module top( in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ , out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ );
  input in_15_ , in_0_ , in_4_ , in_29_ , in_38_ , in_53_ , in_42_ , in_11_ , in_59_ , in_48_ , in_54_ , in_16_ , in_43_ , in_37_ , in_61_ , in_14_ , in_62_ , in_60_ , in_40_ , in_5_ , in_28_ , in_7_ , in_6_ , in_34_ , in_57_ , in_3_ , in_56_ , in_45_ , in_10_ , in_27_ , in_21_ , in_25_ , in_22_ , in_12_ , in_58_ , in_36_ , in_51_ , in_18_ , in_9_ , in_39_ , in_24_ , in_26_ , in_8_ , in_41_ , in_55_ , in_2_ , in_49_ , in_19_ , in_35_ , in_50_ , in_32_ , in_30_ , in_33_ , in_17_ , in_31_ , in_44_ , in_1_ , in_23_ , in_52_ , in_20_ , in_46_ , in_13_ , in_63_ , in_47_ ;
  output out_1_ , out_3_ , out_6_ , out_2_ , out_0_ , out_4_ , out_5_ ;
  wire n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 ;
  assign n65 = in_15_ & in_14_ ;
  assign n66 = in_12_ | in_13_ ;
  assign n67 = in_4_ | in_5_ ;
  assign n68 = in_0_ | in_1_ ;
  assign n69 = in_3_ & in_2_ ;
  assign n70 = ( n67 & n68 ) | ( n67 & n69 ) | ( n68 & n69 ) ;
  assign n71 = ( ~n67 & n68 ) | ( ~n67 & n69 ) | ( n68 & n69 ) ;
  assign n72 = ( n67 & ~n70 ) | ( n67 & n71 ) | ( ~n70 & n71 ) ;
  assign n73 = in_11_ & in_10_ ;
  assign n74 = in_7_ & in_6_ ;
  assign n75 = in_9_ | in_8_ ;
  assign n76 = ( n73 & n74 ) | ( n73 & n75 ) | ( n74 & n75 ) ;
  assign n77 = ( ~n73 & n74 ) | ( ~n73 & n75 ) | ( n74 & n75 ) ;
  assign n78 = ( n73 & ~n76 ) | ( n73 & n77 ) | ( ~n76 & n77 ) ;
  assign n79 = ( n66 & n72 ) | ( n66 & n78 ) | ( n72 & n78 ) ;
  assign n80 = ( ~n66 & n72 ) | ( ~n66 & n78 ) | ( n72 & n78 ) ;
  assign n81 = ( n66 & ~n79 ) | ( n66 & n80 ) | ( ~n79 & n80 ) ;
  assign n82 = n65 & n81 ;
  assign n83 = n65 | n81 ;
  assign n84 = ~n82 & n83 ;
  assign n85 = in_30_ & in_31_ ;
  assign n86 = in_29_ | in_28_ ;
  assign n87 = in_21_ | in_20_ ;
  assign n88 = in_16_ | in_17_ ;
  assign n89 = in_18_ & in_19_ ;
  assign n90 = ( n87 & n88 ) | ( n87 & n89 ) | ( n88 & n89 ) ;
  assign n91 = ( ~n87 & n88 ) | ( ~n87 & n89 ) | ( n88 & n89 ) ;
  assign n92 = ( n87 & ~n90 ) | ( n87 & n91 ) | ( ~n90 & n91 ) ;
  assign n93 = in_27_ & in_26_ ;
  assign n94 = in_22_ & in_23_ ;
  assign n95 = in_25_ | in_24_ ;
  assign n96 = ( n93 & n94 ) | ( n93 & n95 ) | ( n94 & n95 ) ;
  assign n97 = ( ~n93 & n94 ) | ( ~n93 & n95 ) | ( n94 & n95 ) ;
  assign n98 = ( n93 & ~n96 ) | ( n93 & n97 ) | ( ~n96 & n97 ) ;
  assign n99 = ( n86 & n92 ) | ( n86 & n98 ) | ( n92 & n98 ) ;
  assign n100 = ( ~n86 & n92 ) | ( ~n86 & n98 ) | ( n92 & n98 ) ;
  assign n101 = ( n86 & ~n99 ) | ( n86 & n100 ) | ( ~n99 & n100 ) ;
  assign n102 = n85 & n101 ;
  assign n103 = n85 | n101 ;
  assign n104 = ~n102 & n103 ;
  assign n105 = n84 & n104 ;
  assign n106 = n84 | n104 ;
  assign n107 = ~n105 & n106 ;
  assign n108 = in_46_ & in_47_ ;
  assign n109 = in_45_ | in_44_ ;
  assign n110 = in_37_ | in_36_ ;
  assign n111 = in_32_ | in_33_ ;
  assign n112 = in_34_ & in_35_ ;
  assign n113 = ( n110 & n111 ) | ( n110 & n112 ) | ( n111 & n112 ) ;
  assign n114 = ( ~n110 & n111 ) | ( ~n110 & n112 ) | ( n111 & n112 ) ;
  assign n115 = ( n110 & ~n113 ) | ( n110 & n114 ) | ( ~n113 & n114 ) ;
  assign n116 = in_42_ & in_43_ ;
  assign n117 = in_38_ & in_39_ ;
  assign n118 = in_40_ | in_41_ ;
  assign n119 = ( n116 & n117 ) | ( n116 & n118 ) | ( n117 & n118 ) ;
  assign n120 = ( ~n116 & n117 ) | ( ~n116 & n118 ) | ( n117 & n118 ) ;
  assign n121 = ( n116 & ~n119 ) | ( n116 & n120 ) | ( ~n119 & n120 ) ;
  assign n122 = ( n109 & n115 ) | ( n109 & n121 ) | ( n115 & n121 ) ;
  assign n123 = ( ~n109 & n115 ) | ( ~n109 & n121 ) | ( n115 & n121 ) ;
  assign n124 = ( n109 & ~n122 ) | ( n109 & n123 ) | ( ~n122 & n123 ) ;
  assign n125 = n108 & n124 ;
  assign n126 = n108 | n124 ;
  assign n127 = ~n125 & n126 ;
  assign n128 = in_62_ & in_63_ ;
  assign n129 = in_61_ | in_60_ ;
  assign n130 = in_53_ | in_52_ ;
  assign n131 = in_48_ | in_49_ ;
  assign n132 = in_51_ & in_50_ ;
  assign n133 = ( n130 & n131 ) | ( n130 & n132 ) | ( n131 & n132 ) ;
  assign n134 = ( ~n130 & n131 ) | ( ~n130 & n132 ) | ( n131 & n132 ) ;
  assign n135 = ( n130 & ~n133 ) | ( n130 & n134 ) | ( ~n133 & n134 ) ;
  assign n136 = in_59_ & in_58_ ;
  assign n137 = in_54_ & in_55_ ;
  assign n138 = in_57_ | in_56_ ;
  assign n139 = ( n136 & n137 ) | ( n136 & n138 ) | ( n137 & n138 ) ;
  assign n140 = ( ~n136 & n137 ) | ( ~n136 & n138 ) | ( n137 & n138 ) ;
  assign n141 = ( n136 & ~n139 ) | ( n136 & n140 ) | ( ~n139 & n140 ) ;
  assign n142 = ( n129 & n135 ) | ( n129 & n141 ) | ( n135 & n141 ) ;
  assign n143 = ( ~n129 & n135 ) | ( ~n129 & n141 ) | ( n135 & n141 ) ;
  assign n144 = ( n129 & ~n142 ) | ( n129 & n143 ) | ( ~n142 & n143 ) ;
  assign n145 = n128 | n144 ;
  assign n146 = n128 & n144 ;
  assign n147 = n145 & ~n146 ;
  assign n148 = n127 & n147 ;
  assign n149 = n127 | n147 ;
  assign n150 = ~n148 & n149 ;
  assign n151 = n107 & n150 ;
  assign n152 = n107 | n150 ;
  assign n153 = ~n151 & n152 ;
  assign n154 = ( n70 & n76 ) | ( n70 & n79 ) | ( n76 & n79 ) ;
  assign n155 = ( n70 & n76 ) | ( n70 & ~n79 ) | ( n76 & ~n79 ) ;
  assign n156 = ( n79 & ~n154 ) | ( n79 & n155 ) | ( ~n154 & n155 ) ;
  assign n157 = n82 & n156 ;
  assign n158 = n154 & n157 ;
  assign n159 = n154 | n157 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = ( n90 & n96 ) | ( n90 & n99 ) | ( n96 & n99 ) ;
  assign n162 = ( n90 & n96 ) | ( n90 & ~n99 ) | ( n96 & ~n99 ) ;
  assign n163 = ( n99 & ~n161 ) | ( n99 & n162 ) | ( ~n161 & n162 ) ;
  assign n164 = n102 & n163 ;
  assign n165 = n161 & n164 ;
  assign n166 = n161 | n164 ;
  assign n167 = ~n165 & n166 ;
  assign n168 = n160 & n167 ;
  assign n169 = n160 | n167 ;
  assign n170 = ~n168 & n169 ;
  assign n171 = n82 | n156 ;
  assign n172 = ~n157 & n171 ;
  assign n173 = n102 | n163 ;
  assign n174 = ~n164 & n173 ;
  assign n175 = ( n105 & n172 ) | ( n105 & n174 ) | ( n172 & n174 ) ;
  assign n176 = n170 & n175 ;
  assign n177 = n170 | n175 ;
  assign n178 = ~n176 & n177 ;
  assign n179 = ( n113 & n119 ) | ( n113 & n122 ) | ( n119 & n122 ) ;
  assign n180 = ( n113 & n119 ) | ( n113 & ~n122 ) | ( n119 & ~n122 ) ;
  assign n181 = ( n122 & ~n179 ) | ( n122 & n180 ) | ( ~n179 & n180 ) ;
  assign n182 = n125 & n181 ;
  assign n183 = n179 & n182 ;
  assign n184 = n179 | n182 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = ( n133 & n139 ) | ( n133 & n142 ) | ( n139 & n142 ) ;
  assign n187 = ( n133 & n139 ) | ( n133 & ~n142 ) | ( n139 & ~n142 ) ;
  assign n188 = ( n142 & ~n186 ) | ( n142 & n187 ) | ( ~n186 & n187 ) ;
  assign n189 = n146 & n188 ;
  assign n190 = n186 & n189 ;
  assign n191 = n186 | n189 ;
  assign n192 = ~n190 & n191 ;
  assign n193 = n185 & n192 ;
  assign n194 = n185 | n192 ;
  assign n195 = ~n193 & n194 ;
  assign n196 = n125 | n181 ;
  assign n197 = ~n182 & n196 ;
  assign n198 = n146 | n188 ;
  assign n199 = ~n189 & n198 ;
  assign n200 = ( n148 & n197 ) | ( n148 & n199 ) | ( n197 & n199 ) ;
  assign n201 = n195 & n200 ;
  assign n202 = n195 | n200 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = n178 & n203 ;
  assign n205 = n178 | n203 ;
  assign n206 = ~n204 & n205 ;
  assign n207 = n172 & n174 ;
  assign n208 = n172 | n174 ;
  assign n209 = ~n207 & n208 ;
  assign n210 = n105 & n209 ;
  assign n211 = n105 | n209 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n197 & n199 ;
  assign n214 = n197 | n199 ;
  assign n215 = ~n213 & n214 ;
  assign n216 = n148 & n215 ;
  assign n217 = n148 | n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = ( n151 & n212 ) | ( n151 & n218 ) | ( n212 & n218 ) ;
  assign n220 = n206 & n219 ;
  assign n221 = n206 | n219 ;
  assign n222 = ~n220 & n221 ;
  assign n223 = ( n160 & n167 ) | ( n160 & n175 ) | ( n167 & n175 ) ;
  assign n224 = ( n158 & n165 ) | ( n158 & n223 ) | ( n165 & n223 ) ;
  assign n225 = ( n185 & n192 ) | ( n185 & n200 ) | ( n192 & n200 ) ;
  assign n226 = ( n183 & n190 ) | ( n183 & n225 ) | ( n190 & n225 ) ;
  assign n227 = n158 & n165 ;
  assign n228 = n158 | n165 ;
  assign n229 = ~n227 & n228 ;
  assign n230 = n223 & n229 ;
  assign n231 = n223 | n229 ;
  assign n232 = ~n230 & n231 ;
  assign n233 = n183 & n190 ;
  assign n234 = n183 | n190 ;
  assign n235 = ~n233 & n234 ;
  assign n236 = n225 & n235 ;
  assign n237 = n225 | n235 ;
  assign n238 = ~n236 & n237 ;
  assign n239 = ( n178 & n203 ) | ( n178 & n219 ) | ( n203 & n219 ) ;
  assign n240 = ( n232 & n238 ) | ( n232 & n239 ) | ( n238 & n239 ) ;
  assign n241 = ( n224 & n226 ) | ( n224 & n240 ) | ( n226 & n240 ) ;
  assign n242 = n212 & n218 ;
  assign n243 = n212 | n218 ;
  assign n244 = ~n242 & n243 ;
  assign n245 = n151 & n244 ;
  assign n246 = n151 | n244 ;
  assign n247 = ~n245 & n246 ;
  assign n248 = n232 & n238 ;
  assign n249 = n232 | n238 ;
  assign n250 = ~n248 & n249 ;
  assign n251 = n239 & n250 ;
  assign n252 = n239 | n250 ;
  assign n253 = ~n251 & n252 ;
  assign n254 = n224 & n226 ;
  assign n255 = n224 | n226 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = n240 & n256 ;
  assign n258 = n240 | n256 ;
  assign n259 = ~n257 & n258 ;
  assign out_1_ = n153 ;
  assign out_3_ = n222 ;
  assign out_6_ = n241 ;
  assign out_2_ = n247 ;
  assign out_0_ = 1'b0 ;
  assign out_4_ = n253 ;
  assign out_5_ = n259 ;
endmodule
