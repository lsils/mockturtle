module top( N1 , N100 , N103 , N106 , N109 , N110 , N111 , N112 , N113 , N114 , N115 , N118 , N12 , N121 , N124 , N127 , N130 , N133 , N134 , N135 , N138 , N141 , N144 , N147 , N15 , N150 , N151 , N152 , N153 , N154 , N155 , N156 , N157 , N158 , N159 , N160 , N161 , N162 , N163 , N164 , N165 , N166 , N167 , N168 , N169 , N170 , N171 , N172 , N173 , N174 , N175 , N176 , N177 , N178 , N179 , N18 , N180 , N181 , N182 , N183 , N184 , N185 , N186 , N187 , N188 , N189 , N190 , N191 , N192 , N193 , N194 , N195 , N196 , N197 , N198 , N199 , N200 , N201 , N202 , N203 , N204 , N205 , N206 , N207 , N208 , N209 , N210 , N211 , N212 , N213 , N214 , N215 , N216 , N217 , N218 , N219 , N220 , N221 , N222 , N223 , N224 , N225 , N226 , N227 , N228 , N229 , N23 , N230 , N231 , N232 , N233 , N234 , N235 , N236 , N237 , N238 , N239 , N240 , N241_I , N242 , N245 , N248 , N251 , N254 , N257 , N26 , N260 , N263 , N267 , N271 , N274 , N277 , N280 , N283 , N286 , N289 , N29 , N293 , N296 , N299 , N303 , N307 , N310 , N313 , N316 , N319 , N32 , N322 , N325 , N328 , N331 , N334 , N337 , N340 , N343 , N346 , N349 , N35 , N352 , N355 , N358 , N361 , N364 , N367 , N38 , N382 , N41 , N44 , N47 , N5 , N50 , N53 , N54 , N55 , N56 , N57 , N58 , N59 , N60 , N61 , N62 , N63 , N64 , N65 , N66 , N69 , N70 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 , N85 , N86 , N87 , N88 , N89 , N9 , N94 , N97 , N10025 , N10101 , N10102 , N10103 , N10104 , N10109 , N10110 , N10111 , N10112 , N10350 , N10351 , N10352 , N10353 , N10574 , N10575 , N10576 , N10628 , N10632 , N10641 , N10704 , N10706 , N10711 , N10712 , N10713 , N10714 , N10715 , N10716 , N10717 , N10718 , N10729 , N10759 , N10760 , N10761 , N10762 , N10763 , N10827 , N10837 , N10838 , N10839 , N10840 , N10868 , N10869 , N10870 , N10871 , N10905 , N10906 , N10907 , N10908 , N1110 , N1111 , N1112 , N1113 , N1114 , N11333 , N11334 , N11340 , N11342 , N1489 , N1490 , N1781 , N241_O , N387 , N388 , N478 , N482 , N484 , N486 , N489 , N492 , N501 , N505 , N507 , N509 , N511 , N513 , N515 , N517 , N519 , N535 , N537 , N539 , N541 , N543 , N545 , N547 , N549 , N551 , N553 , N556 , N559 , N561 , N563 , N565 , N567 , N569 , N571 , N573 , N582 , N643 , N707 , N813 , N881 , N882 , N883 , N884 , N885 , N889 , N945 );
  input N1 , N100 , N103 , N106 , N109 , N110 , N111 , N112 , N113 , N114 , N115 , N118 , N12 , N121 , N124 , N127 , N130 , N133 , N134 , N135 , N138 , N141 , N144 , N147 , N15 , N150 , N151 , N152 , N153 , N154 , N155 , N156 , N157 , N158 , N159 , N160 , N161 , N162 , N163 , N164 , N165 , N166 , N167 , N168 , N169 , N170 , N171 , N172 , N173 , N174 , N175 , N176 , N177 , N178 , N179 , N18 , N180 , N181 , N182 , N183 , N184 , N185 , N186 , N187 , N188 , N189 , N190 , N191 , N192 , N193 , N194 , N195 , N196 , N197 , N198 , N199 , N200 , N201 , N202 , N203 , N204 , N205 , N206 , N207 , N208 , N209 , N210 , N211 , N212 , N213 , N214 , N215 , N216 , N217 , N218 , N219 , N220 , N221 , N222 , N223 , N224 , N225 , N226 , N227 , N228 , N229 , N23 , N230 , N231 , N232 , N233 , N234 , N235 , N236 , N237 , N238 , N239 , N240 , N241_I , N242 , N245 , N248 , N251 , N254 , N257 , N26 , N260 , N263 , N267 , N271 , N274 , N277 , N280 , N283 , N286 , N289 , N29 , N293 , N296 , N299 , N303 , N307 , N310 , N313 , N316 , N319 , N32 , N322 , N325 , N328 , N331 , N334 , N337 , N340 , N343 , N346 , N349 , N35 , N352 , N355 , N358 , N361 , N364 , N367 , N38 , N382 , N41 , N44 , N47 , N5 , N50 , N53 , N54 , N55 , N56 , N57 , N58 , N59 , N60 , N61 , N62 , N63 , N64 , N65 , N66 , N69 , N70 , N73 , N74 , N75 , N76 , N77 , N78 , N79 , N80 , N81 , N82 , N83 , N84 , N85 , N86 , N87 , N88 , N89 , N9 , N94 , N97 ;
  output N10025 , N10101 , N10102 , N10103 , N10104 , N10109 , N10110 , N10111 , N10112 , N10350 , N10351 , N10352 , N10353 , N10574 , N10575 , N10576 , N10628 , N10632 , N10641 , N10704 , N10706 , N10711 , N10712 , N10713 , N10714 , N10715 , N10716 , N10717 , N10718 , N10729 , N10759 , N10760 , N10761 , N10762 , N10763 , N10827 , N10837 , N10838 , N10839 , N10840 , N10868 , N10869 , N10870 , N10871 , N10905 , N10906 , N10907 , N10908 , N1110 , N1111 , N1112 , N1113 , N1114 , N11333 , N11334 , N11340 , N11342 , N1489 , N1490 , N1781 , N241_O , N387 , N388 , N478 , N482 , N484 , N486 , N489 , N492 , N501 , N505 , N507 , N509 , N511 , N513 , N515 , N517 , N519 , N535 , N537 , N539 , N541 , N543 , N545 , N547 , N549 , N551 , N553 , N556 , N559 , N561 , N563 , N565 , N567 , N569 , N571 , N573 , N582 , N643 , N707 , N813 , N881 , N882 , N883 , N884 , N885 , N889 , N945 ;
  wire n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 ;
  assign n208 = ~N18 & N41 ;
  assign n209 = ~N310 & n208 ;
  assign n210 = N18 | N41 ;
  assign n211 = N310 & ~n210 ;
  assign n212 = n209 | n211 ;
  assign n213 = N367 & ~n212 ;
  assign n214 = ~N367 & n212 ;
  assign n215 = n213 | n214 ;
  assign n216 = N267 & N382 ;
  assign n217 = ~N38 & n216 ;
  assign n218 = N263 & n216 ;
  assign n219 = N38 & ~n218 ;
  assign n220 = N263 & N382 ;
  assign n221 = N38 & n220 ;
  assign n222 = N38 | n220 ;
  assign n223 = ~n221 & n222 ;
  assign n224 = N12 & N9 ;
  assign n225 = N18 & ~N213 ;
  assign n226 = n224 | n225 ;
  assign n227 = N260 | n226 ;
  assign n228 = N18 & ~N214 ;
  assign n229 = n224 | n228 ;
  assign n230 = N257 | n229 ;
  assign n231 = N260 & n226 ;
  assign n232 = n230 | n231 ;
  assign n233 = n227 & n232 ;
  assign n234 = N18 & ~N215 ;
  assign n235 = n224 | n234 ;
  assign n236 = N106 | n235 ;
  assign n237 = N106 & n235 ;
  assign n238 = N18 & ~N216 ;
  assign n239 = n224 | n238 ;
  assign n240 = N254 & n239 ;
  assign n241 = N18 & ~N209 ;
  assign n242 = n224 | n241 ;
  assign n243 = N251 | n242 ;
  assign n244 = N254 | n239 ;
  assign n245 = n243 & n244 ;
  assign n246 = n240 | n245 ;
  assign n247 = n237 | n246 ;
  assign n248 = n236 & n247 ;
  assign n249 = N257 & n229 ;
  assign n250 = n230 & ~n249 ;
  assign n251 = n227 & ~n231 ;
  assign n252 = n250 & n251 ;
  assign n253 = ~n248 & n252 ;
  assign n254 = n233 & ~n253 ;
  assign n255 = ~N153 & N18 ;
  assign n256 = n224 | n255 ;
  assign n257 = N303 & n256 ;
  assign n258 = N303 | n256 ;
  assign n259 = ~N154 & N18 ;
  assign n260 = n224 | n259 ;
  assign n261 = N299 & n260 ;
  assign n262 = N299 | n260 ;
  assign n263 = ~N155 & N18 ;
  assign n264 = n224 | n263 ;
  assign n265 = N296 & n264 ;
  assign n266 = N296 | n264 ;
  assign n267 = ~N156 & N18 ;
  assign n268 = n224 | n267 ;
  assign n269 = N293 | n268 ;
  assign n270 = n266 & n269 ;
  assign n271 = n265 | n270 ;
  assign n272 = n262 & n271 ;
  assign n273 = n261 | n272 ;
  assign n274 = N293 & n268 ;
  assign n275 = n265 | n274 ;
  assign n276 = n270 & ~n275 ;
  assign n277 = ~n261 & n262 ;
  assign n278 = n276 & n277 ;
  assign n279 = n273 & ~n278 ;
  assign n280 = ~N157 & N18 ;
  assign n281 = n224 | n280 ;
  assign n282 = N289 & n281 ;
  assign n283 = N289 | n281 ;
  assign n284 = N135 & ~N18 ;
  assign n285 = N158 & N18 ;
  assign n286 = n284 | n285 ;
  assign n287 = N286 & ~n286 ;
  assign n288 = ~N286 & n286 ;
  assign n289 = N144 & ~N18 ;
  assign n290 = N159 & N18 ;
  assign n291 = n289 | n290 ;
  assign n292 = ~N283 & n291 ;
  assign n293 = N283 & ~n291 ;
  assign n294 = N138 & ~N18 ;
  assign n295 = N160 & N18 ;
  assign n296 = n294 | n295 ;
  assign n297 = ~N280 & n296 ;
  assign n298 = N147 & ~N18 ;
  assign n299 = N151 & N18 ;
  assign n300 = n298 | n299 ;
  assign n301 = ~N277 & n300 ;
  assign n302 = N280 & ~n296 ;
  assign n303 = n301 & ~n302 ;
  assign n304 = n297 | n303 ;
  assign n305 = ~n293 & n304 ;
  assign n306 = n292 | n305 ;
  assign n307 = n288 | n306 ;
  assign n308 = ~n287 & n307 ;
  assign n309 = n283 & ~n308 ;
  assign n310 = N277 & ~n300 ;
  assign n311 = n301 | n310 ;
  assign n312 = n297 | n302 ;
  assign n313 = n311 | n312 ;
  assign n314 = n287 | n288 ;
  assign n315 = n292 | n293 ;
  assign n316 = n314 | n315 ;
  assign n317 = n313 | n316 ;
  assign n318 = n309 & n317 ;
  assign n319 = n282 | n318 ;
  assign n320 = N18 & N219 ;
  assign n321 = ~N18 & N66 ;
  assign n322 = n320 | n321 ;
  assign n323 = ~N364 & n322 ;
  assign n324 = N364 & ~n322 ;
  assign n325 = N18 & N220 ;
  assign n326 = ~N18 & N50 ;
  assign n327 = n325 | n326 ;
  assign n328 = N361 & ~n327 ;
  assign n329 = ~N361 & n327 ;
  assign n330 = N18 & N221 ;
  assign n331 = ~N18 & N32 ;
  assign n332 = n330 | n331 ;
  assign n333 = N358 & ~n332 ;
  assign n334 = ~N358 & n332 ;
  assign n335 = N18 & N222 ;
  assign n336 = ~N18 & N35 ;
  assign n337 = n335 | n336 ;
  assign n338 = ~N355 & n337 ;
  assign n339 = n334 | n338 ;
  assign n340 = ~n333 & n339 ;
  assign n341 = n329 | n340 ;
  assign n342 = ~n328 & n341 ;
  assign n343 = n333 | n334 ;
  assign n344 = N355 & ~n337 ;
  assign n345 = n338 | n344 ;
  assign n346 = n343 | n345 ;
  assign n347 = n328 | n346 ;
  assign n348 = ~n342 & n347 ;
  assign n349 = N18 & N217 ;
  assign n350 = N118 & ~N18 ;
  assign n351 = n349 | n350 ;
  assign n352 = ~N340 & n351 ;
  assign n353 = N18 & N226 ;
  assign n354 = ~N18 & N97 ;
  assign n355 = n353 | n354 ;
  assign n356 = N343 & ~n355 ;
  assign n357 = n352 | n356 ;
  assign n358 = N340 & ~n351 ;
  assign n359 = ~N343 & n355 ;
  assign n360 = n358 | n359 ;
  assign n361 = n357 | n360 ;
  assign n362 = N18 & N224 ;
  assign n363 = N121 & ~N18 ;
  assign n364 = n362 | n363 ;
  assign n365 = N349 & ~n364 ;
  assign n366 = ~N349 & n364 ;
  assign n367 = n365 | n366 ;
  assign n368 = N18 & N225 ;
  assign n369 = ~N18 & N94 ;
  assign n370 = n368 | n369 ;
  assign n371 = N346 & ~n370 ;
  assign n372 = ~N346 & n370 ;
  assign n373 = n371 | n372 ;
  assign n374 = n367 | n373 ;
  assign n375 = n361 | n374 ;
  assign n376 = N18 & N223 ;
  assign n377 = ~N18 & N47 ;
  assign n378 = n376 | n377 ;
  assign n379 = ~N352 & n378 ;
  assign n380 = N352 & ~n378 ;
  assign n381 = n379 | n380 ;
  assign n382 = n375 | n381 ;
  assign n383 = N18 & N231 ;
  assign n384 = N100 & ~N18 ;
  assign n385 = n383 | n384 ;
  assign n386 = N334 & ~n385 ;
  assign n387 = ~N334 & n385 ;
  assign n388 = N18 & N232 ;
  assign n389 = N124 & ~N18 ;
  assign n390 = n388 | n389 ;
  assign n391 = N331 & ~n390 ;
  assign n392 = ~N331 & n390 ;
  assign n393 = N18 & N233 ;
  assign n394 = N127 & ~N18 ;
  assign n395 = n393 | n394 ;
  assign n396 = N328 & ~n395 ;
  assign n397 = ~N328 & n395 ;
  assign n398 = N18 & N234 ;
  assign n399 = N130 & ~N18 ;
  assign n400 = n398 | n399 ;
  assign n401 = ~N325 & n400 ;
  assign n402 = n397 | n401 ;
  assign n403 = ~n396 & n402 ;
  assign n404 = n392 | n403 ;
  assign n405 = ~n391 & n404 ;
  assign n406 = n387 | n405 ;
  assign n407 = ~n386 & n406 ;
  assign n408 = N18 & N235 ;
  assign n409 = N103 & ~N18 ;
  assign n410 = n408 | n409 ;
  assign n411 = ~N322 & n410 ;
  assign n412 = N322 & ~n410 ;
  assign n413 = N18 & N236 ;
  assign n414 = ~N18 & N23 ;
  assign n415 = n413 | n414 ;
  assign n416 = N319 & ~n415 ;
  assign n417 = ~N319 & n415 ;
  assign n418 = N18 & N237 ;
  assign n419 = ~N18 & N26 ;
  assign n420 = n418 | n419 ;
  assign n421 = N316 & ~n420 ;
  assign n422 = N18 & N238 ;
  assign n423 = ~N18 & N29 ;
  assign n424 = n422 | n423 ;
  assign n425 = N313 & ~n424 ;
  assign n426 = n209 & ~n425 ;
  assign n427 = ~N316 & n420 ;
  assign n428 = ~N313 & n424 ;
  assign n429 = n427 | n428 ;
  assign n430 = n426 | n429 ;
  assign n431 = ~n421 & n430 ;
  assign n432 = n417 | n431 ;
  assign n433 = ~n416 & n432 ;
  assign n434 = ~n412 & n433 ;
  assign n435 = n411 | n434 ;
  assign n436 = N367 | n435 ;
  assign n437 = n421 | n427 ;
  assign n438 = n425 | n428 ;
  assign n439 = n212 | n438 ;
  assign n440 = n437 | n439 ;
  assign n441 = n416 | n417 ;
  assign n442 = n440 | n441 ;
  assign n443 = ~n433 & n442 ;
  assign n444 = n412 | n443 ;
  assign n445 = ~n411 & n444 ;
  assign n446 = n436 & ~n445 ;
  assign n447 = n396 | n397 ;
  assign n448 = N325 & ~n400 ;
  assign n449 = n401 | n448 ;
  assign n450 = n447 | n449 ;
  assign n451 = n391 | n392 ;
  assign n452 = n386 | n387 ;
  assign n453 = n451 | n452 ;
  assign n454 = n450 | n453 ;
  assign n455 = n446 & ~n454 ;
  assign n456 = n407 | n455 ;
  assign n457 = ~n382 & n456 ;
  assign n458 = n352 | n359 ;
  assign n459 = ~n356 & n458 ;
  assign n460 = ~n371 & n459 ;
  assign n461 = n372 | n460 ;
  assign n462 = ~n365 & n461 ;
  assign n463 = n366 | n462 ;
  assign n464 = ~n380 & n463 ;
  assign n465 = n379 | n464 ;
  assign n466 = n457 | n465 ;
  assign n467 = n342 | n466 ;
  assign n468 = ~n348 & n467 ;
  assign n469 = ~n324 & n468 ;
  assign n470 = n323 | n469 ;
  assign n471 = n309 & ~n470 ;
  assign n472 = n319 | n471 ;
  assign n473 = n273 & n472 ;
  assign n474 = n279 | n473 ;
  assign n475 = n258 & n474 ;
  assign n476 = n257 | n475 ;
  assign n477 = n236 & ~n237 ;
  assign n478 = N251 & n242 ;
  assign n479 = n243 & ~n478 ;
  assign n480 = ~n240 & n244 ;
  assign n481 = n479 & n480 ;
  assign n482 = n477 & n481 ;
  assign n483 = ~n476 & n482 ;
  assign n484 = n252 & n483 ;
  assign n485 = n254 & ~n484 ;
  assign n486 = n223 | n485 ;
  assign n487 = ~n219 & n486 ;
  assign n488 = n217 | n487 ;
  assign n489 = N245 & N271 ;
  assign n490 = ~N38 & N382 ;
  assign n491 = ~n489 & n490 ;
  assign n492 = ~N18 & N53 ;
  assign n493 = N18 & ~N325 ;
  assign n494 = n492 | n493 ;
  assign n495 = N18 & N203 ;
  assign n496 = n399 | n495 ;
  assign n497 = n494 | n496 ;
  assign n498 = ~N18 & N73 ;
  assign n499 = N18 & ~N322 ;
  assign n500 = n498 | n499 ;
  assign n501 = N18 & N204 ;
  assign n502 = n409 | n501 ;
  assign n503 = n500 & n502 ;
  assign n504 = ~N18 & N74 ;
  assign n505 = N18 & ~N313 ;
  assign n506 = n504 | n505 ;
  assign n507 = N18 & N207 ;
  assign n508 = n423 | n507 ;
  assign n509 = n506 & n508 ;
  assign n510 = N70 | N89 ;
  assign n511 = n208 & n510 ;
  assign n512 = N18 | N70 ;
  assign n513 = N89 & n512 ;
  assign n514 = n511 | n513 ;
  assign n515 = n509 | n514 ;
  assign n516 = ~N18 & N76 ;
  assign n517 = N18 & ~N316 ;
  assign n518 = n516 | n517 ;
  assign n519 = N18 & N206 ;
  assign n520 = n419 | n519 ;
  assign n521 = n518 | n520 ;
  assign n522 = n506 | n508 ;
  assign n523 = n521 & n522 ;
  assign n524 = n515 & n523 ;
  assign n525 = n518 & n520 ;
  assign n526 = ~N18 & N75 ;
  assign n527 = N18 & ~N319 ;
  assign n528 = n526 | n527 ;
  assign n529 = N18 & N205 ;
  assign n530 = n414 | n529 ;
  assign n531 = n528 & n530 ;
  assign n532 = n525 | n531 ;
  assign n533 = n524 | n532 ;
  assign n534 = n500 | n502 ;
  assign n535 = n528 | n530 ;
  assign n536 = n534 & n535 ;
  assign n537 = n533 & n536 ;
  assign n538 = n503 | n537 ;
  assign n539 = n497 & n538 ;
  assign n540 = ~N18 & N54 ;
  assign n541 = N18 & ~N328 ;
  assign n542 = n540 | n541 ;
  assign n543 = N18 & N202 ;
  assign n544 = n394 | n543 ;
  assign n545 = n542 & n544 ;
  assign n546 = n494 & n496 ;
  assign n547 = n545 | n546 ;
  assign n548 = n539 | n547 ;
  assign n549 = ~N18 & N56 ;
  assign n550 = N18 & ~N334 ;
  assign n551 = n549 | n550 ;
  assign n552 = N18 & N200 ;
  assign n553 = n384 | n552 ;
  assign n554 = n551 | n553 ;
  assign n555 = ~N18 & N55 ;
  assign n556 = N18 & ~N331 ;
  assign n557 = n555 | n556 ;
  assign n558 = N18 & N201 ;
  assign n559 = n389 | n558 ;
  assign n560 = n557 & n559 ;
  assign n561 = n554 & ~n560 ;
  assign n562 = n542 | n544 ;
  assign n563 = n557 | n559 ;
  assign n564 = n562 & n563 ;
  assign n565 = n561 & n564 ;
  assign n566 = n548 & n565 ;
  assign n567 = n554 & n560 ;
  assign n568 = n551 & n553 ;
  assign n569 = ~N18 & N77 ;
  assign n570 = N18 & ~N340 ;
  assign n571 = n569 | n570 ;
  assign n572 = N18 & N187 ;
  assign n573 = n350 | n572 ;
  assign n574 = n571 & n573 ;
  assign n575 = n568 | n574 ;
  assign n576 = n567 | n575 ;
  assign n577 = n566 | n576 ;
  assign n578 = ~N18 & N81 ;
  assign n579 = N18 & ~N349 ;
  assign n580 = n578 | n579 ;
  assign n581 = N18 & N194 ;
  assign n582 = n363 | n581 ;
  assign n583 = n580 & n582 ;
  assign n584 = ~N18 & N80 ;
  assign n585 = N18 & ~N352 ;
  assign n586 = n584 | n585 ;
  assign n587 = N18 & N193 ;
  assign n588 = n377 | n587 ;
  assign n589 = n586 & n588 ;
  assign n590 = n583 | n589 ;
  assign n591 = ~N18 & N59 ;
  assign n592 = N18 & ~N346 ;
  assign n593 = n591 | n592 ;
  assign n594 = N18 & N195 ;
  assign n595 = n369 | n594 ;
  assign n596 = n593 | n595 ;
  assign n597 = n580 | n582 ;
  assign n598 = n586 | n588 ;
  assign n599 = n597 & n598 ;
  assign n600 = n596 & n599 ;
  assign n601 = ~n590 & n600 ;
  assign n602 = ~N18 & N78 ;
  assign n603 = N18 & ~N343 ;
  assign n604 = n602 | n603 ;
  assign n605 = N18 & N196 ;
  assign n606 = n354 | n605 ;
  assign n607 = n604 & n606 ;
  assign n608 = n593 & n595 ;
  assign n609 = n607 | n608 ;
  assign n610 = n571 | n573 ;
  assign n611 = n604 | n606 ;
  assign n612 = n610 & n611 ;
  assign n613 = ~n609 & n612 ;
  assign n614 = n601 & n613 ;
  assign n615 = n577 & n614 ;
  assign n616 = n601 & n609 ;
  assign n617 = n590 & n598 ;
  assign n618 = n616 | n617 ;
  assign n619 = n615 | n618 ;
  assign n620 = ~N18 & N62 ;
  assign n621 = N18 & ~N364 ;
  assign n622 = n620 | n621 ;
  assign n623 = N18 & N189 ;
  assign n624 = n321 | n623 ;
  assign n625 = n622 | n624 ;
  assign n626 = ~N18 & N61 ;
  assign n627 = N18 & ~N361 ;
  assign n628 = n626 | n627 ;
  assign n629 = N18 & N190 ;
  assign n630 = n326 | n629 ;
  assign n631 = n628 & n630 ;
  assign n632 = n625 & ~n631 ;
  assign n633 = n622 & n624 ;
  assign n634 = n628 | n630 ;
  assign n635 = ~n633 & n634 ;
  assign n636 = n632 & n635 ;
  assign n637 = ~N18 & N60 ;
  assign n638 = N18 & ~N358 ;
  assign n639 = n637 | n638 ;
  assign n640 = N18 & N191 ;
  assign n641 = n331 | n640 ;
  assign n642 = n639 & n641 ;
  assign n643 = ~N18 & N79 ;
  assign n644 = N18 & ~N355 ;
  assign n645 = n643 | n644 ;
  assign n646 = N18 & N192 ;
  assign n647 = n336 | n646 ;
  assign n648 = n645 & n647 ;
  assign n649 = n642 | n648 ;
  assign n650 = n639 | n641 ;
  assign n651 = n645 | n647 ;
  assign n652 = n650 & n651 ;
  assign n653 = ~n649 & n652 ;
  assign n654 = n636 & n653 ;
  assign n655 = n619 & n654 ;
  assign n656 = n649 & n650 ;
  assign n657 = n636 & n656 ;
  assign n658 = n625 & n631 ;
  assign n659 = n633 | n658 ;
  assign n660 = n657 | n659 ;
  assign n661 = n655 | n660 ;
  assign n662 = ~N18 & N64 ;
  assign n663 = N18 & ~N289 ;
  assign n664 = n662 | n663 ;
  assign n665 = ~N177 & N18 ;
  assign n666 = n224 | n665 ;
  assign n667 = n664 & ~n666 ;
  assign n668 = ~N18 & N85 ;
  assign n669 = N18 & ~N286 ;
  assign n670 = n668 | n669 ;
  assign n671 = N178 & N18 ;
  assign n672 = n284 | n671 ;
  assign n673 = n670 & n672 ;
  assign n674 = n667 | n673 ;
  assign n675 = ~n664 & n666 ;
  assign n676 = n670 | n672 ;
  assign n677 = ~n675 & n676 ;
  assign n678 = ~n674 & n677 ;
  assign n679 = ~N18 & N84 ;
  assign n680 = N18 & ~N283 ;
  assign n681 = n679 | n680 ;
  assign n682 = N179 & N18 ;
  assign n683 = n289 | n682 ;
  assign n684 = n681 & n683 ;
  assign n685 = ~N18 & N83 ;
  assign n686 = N18 & ~N280 ;
  assign n687 = n685 | n686 ;
  assign n688 = N18 & N180 ;
  assign n689 = n294 | n688 ;
  assign n690 = n687 & n689 ;
  assign n691 = n684 | n690 ;
  assign n692 = n681 | n683 ;
  assign n693 = n687 | n689 ;
  assign n694 = n692 & n693 ;
  assign n695 = ~n691 & n694 ;
  assign n696 = n678 & n695 ;
  assign n697 = ~N18 & N65 ;
  assign n698 = N18 & ~N277 ;
  assign n699 = n697 | n698 ;
  assign n700 = N171 & N18 ;
  assign n701 = n298 | n700 ;
  assign n702 = n699 & n701 ;
  assign n703 = n699 | n701 ;
  assign n704 = ~n702 & n703 ;
  assign n705 = n696 & n704 ;
  assign n706 = n661 & n705 ;
  assign n707 = n696 & n702 ;
  assign n708 = n691 & n692 ;
  assign n709 = n678 & n708 ;
  assign n710 = n674 & ~n675 ;
  assign n711 = n709 | n710 ;
  assign n712 = n707 | n711 ;
  assign n713 = n706 | n712 ;
  assign n714 = N109 & ~N18 ;
  assign n715 = N18 & ~N299 ;
  assign n716 = n714 | n715 ;
  assign n717 = ~N174 & N18 ;
  assign n718 = n224 | n717 ;
  assign n719 = n716 & ~n718 ;
  assign n720 = N110 & ~N18 ;
  assign n721 = N18 & ~N303 ;
  assign n722 = n720 | n721 ;
  assign n723 = ~N173 & N18 ;
  assign n724 = n224 | n723 ;
  assign n725 = n722 & ~n724 ;
  assign n726 = n719 | n725 ;
  assign n727 = ~n716 & n718 ;
  assign n728 = ~n722 & n724 ;
  assign n729 = n727 | n728 ;
  assign n730 = n726 | n729 ;
  assign n731 = ~N18 & N86 ;
  assign n732 = N18 & ~N296 ;
  assign n733 = n731 | n732 ;
  assign n734 = ~N175 & N18 ;
  assign n735 = n224 | n734 ;
  assign n736 = n733 & ~n735 ;
  assign n737 = ~N18 & N63 ;
  assign n738 = N18 & ~N293 ;
  assign n739 = n737 | n738 ;
  assign n740 = ~N176 & N18 ;
  assign n741 = n224 | n740 ;
  assign n742 = n739 & ~n741 ;
  assign n743 = n736 | n742 ;
  assign n744 = ~n733 & n735 ;
  assign n745 = ~n739 & n741 ;
  assign n746 = n744 | n745 ;
  assign n747 = n743 | n746 ;
  assign n748 = n730 | n747 ;
  assign n749 = n713 & ~n748 ;
  assign n750 = n743 & ~n744 ;
  assign n751 = ~n730 & n750 ;
  assign n752 = n726 & ~n728 ;
  assign n753 = n751 | n752 ;
  assign n754 = n749 | n753 ;
  assign n755 = ~N18 & N87 ;
  assign n756 = ~N106 & N18 ;
  assign n757 = n755 | n756 ;
  assign n758 = ~N168 & N18 ;
  assign n759 = n224 | n758 ;
  assign n760 = ~n757 & n759 ;
  assign n761 = ~N18 & N88 ;
  assign n762 = N18 & ~N260 ;
  assign n763 = n761 | n762 ;
  assign n764 = ~N166 & N18 ;
  assign n765 = n224 | n764 ;
  assign n766 = ~n763 & n765 ;
  assign n767 = n763 & ~n765 ;
  assign n768 = n766 | n767 ;
  assign n769 = N112 & ~N18 ;
  assign n770 = N18 & ~N257 ;
  assign n771 = n769 | n770 ;
  assign n772 = ~N167 & N18 ;
  assign n773 = n224 | n772 ;
  assign n774 = n771 & ~n773 ;
  assign n775 = ~n771 & n773 ;
  assign n776 = n774 | n775 ;
  assign n777 = n768 | n776 ;
  assign n778 = n760 | n777 ;
  assign n779 = N113 & ~N18 ;
  assign n780 = N18 & ~N251 ;
  assign n781 = n779 | n780 ;
  assign n782 = ~n224 & n781 ;
  assign n783 = N111 & ~N18 ;
  assign n784 = N18 & ~N254 ;
  assign n785 = n783 | n784 ;
  assign n786 = ~N169 & N18 ;
  assign n787 = n224 | n786 ;
  assign n788 = n785 & ~n787 ;
  assign n789 = n782 | n788 ;
  assign n790 = n224 & ~n781 ;
  assign n791 = n757 & ~n759 ;
  assign n792 = ~n785 & n787 ;
  assign n793 = n791 | n792 ;
  assign n794 = n790 | n793 ;
  assign n795 = n789 | n794 ;
  assign n796 = n778 | n795 ;
  assign n797 = n754 & ~n796 ;
  assign n798 = n789 & ~n792 ;
  assign n799 = n791 | n798 ;
  assign n800 = ~n778 & n799 ;
  assign n801 = N245 | N271 ;
  assign n802 = N382 & ~n801 ;
  assign n803 = N38 & ~n802 ;
  assign n804 = n767 | n774 ;
  assign n805 = ~n766 & n804 ;
  assign n806 = n803 | n805 ;
  assign n807 = n800 | n806 ;
  assign n808 = n797 | n807 ;
  assign n809 = ~n491 & n808 ;
  assign n810 = n411 | n412 ;
  assign n811 = N367 & ~n440 ;
  assign n812 = n432 | n811 ;
  assign n813 = ~n416 & n812 ;
  assign n814 = ~n810 & n813 ;
  assign n815 = n810 & ~n813 ;
  assign n816 = n814 | n815 ;
  assign n817 = n431 | n811 ;
  assign n818 = n441 & n817 ;
  assign n819 = n441 | n817 ;
  assign n820 = ~n818 & n819 ;
  assign n821 = n209 | n428 ;
  assign n822 = n213 | n821 ;
  assign n823 = ~n425 & n822 ;
  assign n824 = n437 & n823 ;
  assign n825 = n437 | n823 ;
  assign n826 = ~n824 & n825 ;
  assign n827 = n209 | n213 ;
  assign n828 = n438 | n827 ;
  assign n829 = n438 & n827 ;
  assign n830 = n828 & ~n829 ;
  assign n831 = n450 | n451 ;
  assign n832 = n446 & ~n831 ;
  assign n833 = n405 | n832 ;
  assign n834 = n452 | n833 ;
  assign n835 = n452 & n833 ;
  assign n836 = n834 & ~n835 ;
  assign n837 = n446 & ~n448 ;
  assign n838 = ~n447 & n837 ;
  assign n839 = n403 | n838 ;
  assign n840 = n451 | n839 ;
  assign n841 = n451 & n839 ;
  assign n842 = n840 & ~n841 ;
  assign n843 = n401 | n837 ;
  assign n844 = n447 | n843 ;
  assign n845 = n447 & n843 ;
  assign n846 = n844 & ~n845 ;
  assign n847 = n446 & n449 ;
  assign n848 = n446 | n449 ;
  assign n849 = ~n847 & n848 ;
  assign n850 = n255 & ~n260 ;
  assign n851 = ~n256 & n259 ;
  assign n852 = n850 | n851 ;
  assign n853 = n263 & ~n268 ;
  assign n854 = ~n264 & n267 ;
  assign n855 = n853 | n854 ;
  assign n856 = N141 & ~N18 ;
  assign n857 = N161 & N18 ;
  assign n858 = n856 | n857 ;
  assign n859 = n300 | n858 ;
  assign n860 = n300 & n858 ;
  assign n861 = n859 & ~n860 ;
  assign n862 = n855 | n861 ;
  assign n863 = n855 & n861 ;
  assign n864 = n862 & ~n863 ;
  assign n865 = n852 & ~n864 ;
  assign n866 = ~n852 & n864 ;
  assign n867 = n865 | n866 ;
  assign n868 = n281 & ~n286 ;
  assign n869 = ~n281 & n286 ;
  assign n870 = n868 | n869 ;
  assign n871 = n291 & n296 ;
  assign n872 = n291 | n296 ;
  assign n873 = ~n871 & n872 ;
  assign n874 = n870 & n873 ;
  assign n875 = n870 | n873 ;
  assign n876 = ~n874 & n875 ;
  assign n877 = ~n867 & n876 ;
  assign n878 = ~n224 & n241 ;
  assign n879 = n225 & ~n229 ;
  assign n880 = ~n226 & n228 ;
  assign n881 = n879 | n880 ;
  assign n882 = n878 | n881 ;
  assign n883 = n878 & n881 ;
  assign n884 = n882 & ~n883 ;
  assign n885 = n234 & ~n239 ;
  assign n886 = ~n235 & n238 ;
  assign n887 = n885 | n886 ;
  assign n888 = N18 & ~n224 ;
  assign n889 = N211 | N212 ;
  assign n890 = N211 & N212 ;
  assign n891 = n889 & ~n890 ;
  assign n892 = n888 & n891 ;
  assign n893 = ~n887 & n892 ;
  assign n894 = n887 & ~n892 ;
  assign n895 = n893 | n894 ;
  assign n896 = n884 | n895 ;
  assign n897 = n884 & n895 ;
  assign n898 = n896 & ~n897 ;
  assign n899 = n867 & ~n876 ;
  assign n900 = n898 | n899 ;
  assign n901 = n877 | n900 ;
  assign n902 = N18 & N229 ;
  assign n903 = n208 | n902 ;
  assign n904 = ~n390 & n903 ;
  assign n905 = n390 & ~n903 ;
  assign n906 = n904 | n905 ;
  assign n907 = n385 & ~n415 ;
  assign n908 = ~n385 & n415 ;
  assign n909 = n907 | n908 ;
  assign n910 = ~n906 & n909 ;
  assign n911 = n906 & ~n909 ;
  assign n912 = n910 | n911 ;
  assign n913 = ~n410 & n420 ;
  assign n914 = n410 & ~n420 ;
  assign n915 = n913 | n914 ;
  assign n916 = n395 & ~n400 ;
  assign n917 = ~n395 & n400 ;
  assign n918 = n916 | n917 ;
  assign n919 = N18 & N239 ;
  assign n920 = ~N18 & N44 ;
  assign n921 = n919 | n920 ;
  assign n922 = n424 | n921 ;
  assign n923 = n424 & n921 ;
  assign n924 = n922 & ~n923 ;
  assign n925 = n918 & ~n924 ;
  assign n926 = ~n918 & n924 ;
  assign n927 = n925 | n926 ;
  assign n928 = n915 | n927 ;
  assign n929 = n915 & n927 ;
  assign n930 = n928 & ~n929 ;
  assign n931 = ~n912 & n930 ;
  assign n932 = n912 & ~n930 ;
  assign n933 = n931 | n932 ;
  assign n934 = ~n364 & n378 ;
  assign n935 = n364 & ~n378 ;
  assign n936 = n934 | n935 ;
  assign n937 = n355 & n370 ;
  assign n938 = n355 | n370 ;
  assign n939 = ~n937 & n938 ;
  assign n940 = n936 & ~n939 ;
  assign n941 = ~n936 & n939 ;
  assign n942 = n940 | n941 ;
  assign n943 = N18 & N227 ;
  assign n944 = N115 & ~N18 ;
  assign n945 = n943 | n944 ;
  assign n946 = n351 | n945 ;
  assign n947 = n351 & n945 ;
  assign n948 = n946 & ~n947 ;
  assign n949 = n322 & ~n327 ;
  assign n950 = ~n322 & n327 ;
  assign n951 = n949 | n950 ;
  assign n952 = n332 & n337 ;
  assign n953 = n332 | n337 ;
  assign n954 = ~n952 & n953 ;
  assign n955 = n951 | n954 ;
  assign n956 = n951 & n954 ;
  assign n957 = n955 & ~n956 ;
  assign n958 = ~n948 & n957 ;
  assign n959 = n948 & ~n957 ;
  assign n960 = n958 | n959 ;
  assign n961 = n942 & ~n960 ;
  assign n962 = ~n942 & n960 ;
  assign n963 = n961 | n962 ;
  assign n964 = n933 & n963 ;
  assign n965 = ~n901 & n964 ;
  assign n966 = N114 & ~N18 ;
  assign n967 = N18 & ~N248 ;
  assign n968 = n966 | n967 ;
  assign n969 = n781 & n968 ;
  assign n970 = n781 | n968 ;
  assign n971 = ~n969 & n970 ;
  assign n972 = n763 & ~n771 ;
  assign n973 = ~n763 & n771 ;
  assign n974 = n972 | n973 ;
  assign n975 = ~n971 & n974 ;
  assign n976 = n971 & ~n974 ;
  assign n977 = n975 | n976 ;
  assign n978 = n757 & n785 ;
  assign n979 = n757 | n785 ;
  assign n980 = ~n978 & n979 ;
  assign n981 = N263 & ~N267 ;
  assign n982 = ~N263 & N267 ;
  assign n983 = n981 | n982 ;
  assign n984 = N18 & n983 ;
  assign n985 = N18 | n489 ;
  assign n986 = n801 & ~n985 ;
  assign n987 = n984 | n986 ;
  assign n988 = ~n980 & n987 ;
  assign n989 = n980 & ~n987 ;
  assign n990 = n988 | n989 ;
  assign n991 = ~n977 & n990 ;
  assign n992 = n977 & ~n990 ;
  assign n993 = n991 | n992 ;
  assign n994 = N18 & N310 ;
  assign n995 = n512 & ~n994 ;
  assign n996 = ~N18 & N69 ;
  assign n997 = N18 & ~N307 ;
  assign n998 = n996 | n997 ;
  assign n999 = n995 & n998 ;
  assign n1000 = n995 | n998 ;
  assign n1001 = ~n999 & n1000 ;
  assign n1002 = n506 & n518 ;
  assign n1003 = n506 | n518 ;
  assign n1004 = ~n1002 & n1003 ;
  assign n1005 = n1001 & ~n1004 ;
  assign n1006 = ~n1001 & n1004 ;
  assign n1007 = n1005 | n1006 ;
  assign n1008 = n551 & ~n557 ;
  assign n1009 = ~n551 & n557 ;
  assign n1010 = n1008 | n1009 ;
  assign n1011 = n542 & ~n1010 ;
  assign n1012 = ~n542 & n1010 ;
  assign n1013 = n1011 | n1012 ;
  assign n1014 = n494 & n500 ;
  assign n1015 = n494 | n500 ;
  assign n1016 = ~n1014 & n1015 ;
  assign n1017 = n528 & n1016 ;
  assign n1018 = n528 | n1016 ;
  assign n1019 = ~n1017 & n1018 ;
  assign n1020 = ~n1013 & n1019 ;
  assign n1021 = n1013 & ~n1019 ;
  assign n1022 = n1020 | n1021 ;
  assign n1023 = ~n1007 & n1022 ;
  assign n1024 = n1007 & ~n1022 ;
  assign n1025 = n1023 | n1024 ;
  assign n1026 = n993 & n1025 ;
  assign n1027 = n580 & n586 ;
  assign n1028 = n580 | n586 ;
  assign n1029 = ~n1027 & n1028 ;
  assign n1030 = n622 & ~n628 ;
  assign n1031 = ~n622 & n628 ;
  assign n1032 = n1030 | n1031 ;
  assign n1033 = n1029 | n1032 ;
  assign n1034 = n1029 & n1032 ;
  assign n1035 = n1033 & ~n1034 ;
  assign n1036 = n593 & n604 ;
  assign n1037 = n593 | n604 ;
  assign n1038 = ~n1036 & n1037 ;
  assign n1039 = ~n1035 & n1038 ;
  assign n1040 = n1035 & ~n1038 ;
  assign n1041 = n1039 | n1040 ;
  assign n1042 = n639 & n645 ;
  assign n1043 = n639 | n645 ;
  assign n1044 = ~n1042 & n1043 ;
  assign n1045 = ~N18 & N58 ;
  assign n1046 = N18 & ~N337 ;
  assign n1047 = n1045 | n1046 ;
  assign n1048 = n571 & n1047 ;
  assign n1049 = n571 | n1047 ;
  assign n1050 = ~n1048 & n1049 ;
  assign n1051 = n1044 | n1050 ;
  assign n1052 = n1044 & n1050 ;
  assign n1053 = n1051 & ~n1052 ;
  assign n1054 = n1041 & ~n1053 ;
  assign n1055 = ~n1041 & n1053 ;
  assign n1056 = n1054 | n1055 ;
  assign n1057 = n664 & n670 ;
  assign n1058 = n664 | n670 ;
  assign n1059 = ~n1057 & n1058 ;
  assign n1060 = ~n716 & n722 ;
  assign n1061 = n716 & ~n722 ;
  assign n1062 = n1060 | n1061 ;
  assign n1063 = ~n1059 & n1062 ;
  assign n1064 = n1059 & ~n1062 ;
  assign n1065 = n1063 | n1064 ;
  assign n1066 = ~N18 & N82 ;
  assign n1067 = N18 & ~N274 ;
  assign n1068 = n1066 | n1067 ;
  assign n1069 = n699 & ~n1068 ;
  assign n1070 = ~n699 & n1068 ;
  assign n1071 = n1069 | n1070 ;
  assign n1072 = n681 | n1071 ;
  assign n1073 = n681 & n1071 ;
  assign n1074 = n1072 & ~n1073 ;
  assign n1075 = n733 & ~n739 ;
  assign n1076 = ~n733 & n739 ;
  assign n1077 = n1075 | n1076 ;
  assign n1078 = n687 & n1077 ;
  assign n1079 = n687 | n1077 ;
  assign n1080 = ~n1078 & n1079 ;
  assign n1081 = n1074 & n1080 ;
  assign n1082 = n1074 | n1080 ;
  assign n1083 = ~n1081 & n1082 ;
  assign n1084 = n1065 & n1083 ;
  assign n1085 = n1065 | n1083 ;
  assign n1086 = ~n1084 & n1085 ;
  assign n1087 = n1056 & n1086 ;
  assign n1088 = n1026 & n1087 ;
  assign n1089 = ~N170 & n888 ;
  assign n1090 = n764 & ~n773 ;
  assign n1091 = ~n765 & n772 ;
  assign n1092 = n1090 | n1091 ;
  assign n1093 = ~n1089 & n1092 ;
  assign n1094 = n1089 & ~n1092 ;
  assign n1095 = n1093 | n1094 ;
  assign n1096 = n758 & ~n787 ;
  assign n1097 = ~n759 & n786 ;
  assign n1098 = n1096 | n1097 ;
  assign n1099 = ~N164 & N165 ;
  assign n1100 = N164 & ~N165 ;
  assign n1101 = n1099 | n1100 ;
  assign n1102 = n888 & n1101 ;
  assign n1103 = n1098 | n1102 ;
  assign n1104 = n1098 & n1102 ;
  assign n1105 = n1103 & ~n1104 ;
  assign n1106 = n1095 | n1105 ;
  assign n1107 = n1095 & n1105 ;
  assign n1108 = n1106 & ~n1107 ;
  assign n1109 = n595 & n606 ;
  assign n1110 = n595 | n606 ;
  assign n1111 = ~n1109 & n1110 ;
  assign n1112 = n624 & ~n630 ;
  assign n1113 = ~n624 & n630 ;
  assign n1114 = n1112 | n1113 ;
  assign n1115 = n641 & n647 ;
  assign n1116 = n641 | n647 ;
  assign n1117 = ~n1115 & n1116 ;
  assign n1118 = ~n1114 & n1117 ;
  assign n1119 = n1114 & ~n1117 ;
  assign n1120 = n1118 | n1119 ;
  assign n1121 = n1111 & n1120 ;
  assign n1122 = n1111 | n1120 ;
  assign n1123 = ~n1121 & n1122 ;
  assign n1124 = n582 & n588 ;
  assign n1125 = n582 | n588 ;
  assign n1126 = ~n1124 & n1125 ;
  assign n1127 = N18 & N197 ;
  assign n1128 = n944 | n1127 ;
  assign n1129 = n573 | n1128 ;
  assign n1130 = n573 & n1128 ;
  assign n1131 = n1129 & ~n1130 ;
  assign n1132 = ~n1126 & n1131 ;
  assign n1133 = n1126 & ~n1131 ;
  assign n1134 = n1132 | n1133 ;
  assign n1135 = n1123 | n1134 ;
  assign n1136 = n1123 & n1134 ;
  assign n1137 = n1135 & ~n1136 ;
  assign n1138 = ~n1108 & n1137 ;
  assign n1139 = N18 & N181 ;
  assign n1140 = n856 | n1139 ;
  assign n1141 = n701 & ~n1140 ;
  assign n1142 = ~n701 & n1140 ;
  assign n1143 = n1141 | n1142 ;
  assign n1144 = ~n718 & n723 ;
  assign n1145 = n717 & ~n724 ;
  assign n1146 = n1144 | n1145 ;
  assign n1147 = n734 & ~n741 ;
  assign n1148 = ~n735 & n740 ;
  assign n1149 = n1147 | n1148 ;
  assign n1150 = n1146 | n1149 ;
  assign n1151 = n1146 & n1149 ;
  assign n1152 = n1150 & ~n1151 ;
  assign n1153 = ~n1143 & n1152 ;
  assign n1154 = n1143 & ~n1152 ;
  assign n1155 = n1153 | n1154 ;
  assign n1156 = n666 & n672 ;
  assign n1157 = n666 | n672 ;
  assign n1158 = ~n1156 & n1157 ;
  assign n1159 = n683 & n689 ;
  assign n1160 = n683 | n689 ;
  assign n1161 = ~n1159 & n1160 ;
  assign n1162 = ~n1158 & n1161 ;
  assign n1163 = n1158 & ~n1161 ;
  assign n1164 = n1162 | n1163 ;
  assign n1165 = ~n1155 & n1164 ;
  assign n1166 = n1155 & ~n1164 ;
  assign n1167 = n1165 | n1166 ;
  assign n1168 = N18 & N208 ;
  assign n1169 = n920 | n1168 ;
  assign n1170 = N18 & N198 ;
  assign n1171 = n208 | n1170 ;
  assign n1172 = n1169 | n1171 ;
  assign n1173 = n1169 & n1171 ;
  assign n1174 = n1172 & ~n1173 ;
  assign n1175 = n508 & n520 ;
  assign n1176 = n508 | n520 ;
  assign n1177 = ~n1175 & n1176 ;
  assign n1178 = n502 & ~n530 ;
  assign n1179 = ~n502 & n530 ;
  assign n1180 = n1178 | n1179 ;
  assign n1181 = n1177 | n1180 ;
  assign n1182 = n1177 & n1180 ;
  assign n1183 = n1181 & ~n1182 ;
  assign n1184 = n1174 | n1183 ;
  assign n1185 = n1174 & n1183 ;
  assign n1186 = n1184 & ~n1185 ;
  assign n1187 = n553 & ~n559 ;
  assign n1188 = ~n553 & n559 ;
  assign n1189 = n1187 | n1188 ;
  assign n1190 = n496 & n544 ;
  assign n1191 = n496 | n544 ;
  assign n1192 = ~n1190 & n1191 ;
  assign n1193 = n1189 | n1192 ;
  assign n1194 = n1189 & n1192 ;
  assign n1195 = n1193 & ~n1194 ;
  assign n1196 = n1186 & n1195 ;
  assign n1197 = n1186 | n1195 ;
  assign n1198 = ~n1196 & n1197 ;
  assign n1199 = ~n1167 & n1198 ;
  assign n1200 = n1138 & n1199 ;
  assign n1201 = ~n311 & n470 ;
  assign n1202 = n311 & ~n470 ;
  assign n1203 = n1201 | n1202 ;
  assign n1204 = ~n476 & n479 ;
  assign n1205 = n476 & ~n479 ;
  assign n1206 = n1204 | n1205 ;
  assign n1207 = ~n282 & n283 ;
  assign n1208 = n313 | n315 ;
  assign n1209 = n470 & ~n1208 ;
  assign n1210 = ~n314 & n1209 ;
  assign n1211 = n308 | n1210 ;
  assign n1212 = n1207 & ~n1211 ;
  assign n1213 = ~n1207 & n1211 ;
  assign n1214 = n1212 | n1213 ;
  assign n1215 = n306 | n1209 ;
  assign n1216 = n314 | n1215 ;
  assign n1217 = n314 & n1215 ;
  assign n1218 = n1216 & ~n1217 ;
  assign n1219 = ~n313 & n470 ;
  assign n1220 = n304 | n1219 ;
  assign n1221 = n315 & n1220 ;
  assign n1222 = n315 | n1220 ;
  assign n1223 = ~n1221 & n1222 ;
  assign n1224 = n301 | n1201 ;
  assign n1225 = n312 | n1224 ;
  assign n1226 = n312 & n1224 ;
  assign n1227 = n1225 & ~n1226 ;
  assign n1228 = n248 | n249 ;
  assign n1229 = n230 & n1228 ;
  assign n1230 = n250 & n483 ;
  assign n1231 = n1229 & ~n1230 ;
  assign n1232 = n251 & n1231 ;
  assign n1233 = n251 | n1231 ;
  assign n1234 = ~n1232 & n1233 ;
  assign n1235 = n248 & ~n483 ;
  assign n1236 = n250 | n1235 ;
  assign n1237 = n250 & n1235 ;
  assign n1238 = n1236 & ~n1237 ;
  assign n1239 = ~n476 & n481 ;
  assign n1240 = n246 & ~n1239 ;
  assign n1241 = n477 | n1240 ;
  assign n1242 = n477 & n1240 ;
  assign n1243 = n1241 & ~n1242 ;
  assign n1244 = n243 & ~n1204 ;
  assign n1245 = ~n480 & n1244 ;
  assign n1246 = n480 & ~n1244 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = N150 & N184 ;
  assign n1249 = N228 & N240 ;
  assign n1250 = n1248 & n1249 ;
  assign n1251 = N152 & N210 ;
  assign n1252 = N218 & N230 ;
  assign n1253 = n1251 & n1252 ;
  assign n1254 = n1250 & n1253 ;
  assign n1255 = N182 & N183 ;
  assign n1256 = N185 & N186 ;
  assign n1257 = n1255 & n1256 ;
  assign n1258 = N162 & N172 ;
  assign n1259 = N188 & N199 ;
  assign n1260 = n1258 & n1259 ;
  assign n1261 = n1257 & n1260 ;
  assign n1262 = n1254 & n1261 ;
  assign n1263 = n965 & n1262 ;
  assign n1264 = n1088 & n1200 ;
  assign n1265 = n1263 & n1264 ;
  assign n1266 = ~n257 & n258 ;
  assign n1267 = n474 | n1266 ;
  assign n1268 = n474 & n1266 ;
  assign n1269 = n1267 & ~n1268 ;
  assign n1270 = n276 & ~n472 ;
  assign n1271 = n271 & ~n1270 ;
  assign n1272 = n277 & n1271 ;
  assign n1273 = n277 | n1271 ;
  assign n1274 = ~n1272 & n1273 ;
  assign n1275 = ~n265 & n266 ;
  assign n1276 = n274 | n472 ;
  assign n1277 = n269 & n1276 ;
  assign n1278 = n1275 & ~n1277 ;
  assign n1279 = ~n1275 & n1277 ;
  assign n1280 = n1278 | n1279 ;
  assign n1281 = n269 & ~n274 ;
  assign n1282 = ~n472 & n1281 ;
  assign n1283 = n472 & ~n1281 ;
  assign n1284 = n1282 | n1283 ;
  assign n1285 = n352 | n358 ;
  assign n1286 = n456 & ~n1285 ;
  assign n1287 = ~n456 & n1285 ;
  assign n1288 = n1286 | n1287 ;
  assign n1289 = n221 & n485 ;
  assign n1290 = n222 | n485 ;
  assign n1291 = ~n1289 & n1290 ;
  assign n1292 = n216 & n1291 ;
  assign n1293 = n216 | n1291 ;
  assign n1294 = ~n1292 & n1293 ;
  assign n1295 = n223 & n485 ;
  assign n1296 = n486 & ~n1295 ;
  assign n1297 = ~n375 & n456 ;
  assign n1298 = ~n381 & n463 ;
  assign n1299 = n381 & ~n463 ;
  assign n1300 = n1298 | n1299 ;
  assign n1301 = ~n1297 & n1300 ;
  assign n1302 = n457 | n1301 ;
  assign n1303 = n361 | n373 ;
  assign n1304 = n456 & ~n1303 ;
  assign n1305 = n461 | n1304 ;
  assign n1306 = n367 | n1305 ;
  assign n1307 = n367 & n1305 ;
  assign n1308 = n1306 & ~n1307 ;
  assign n1309 = n356 | n359 ;
  assign n1310 = n1286 & ~n1309 ;
  assign n1311 = n459 | n1310 ;
  assign n1312 = n373 & n1311 ;
  assign n1313 = n373 | n1311 ;
  assign n1314 = ~n1312 & n1313 ;
  assign n1315 = n352 | n1286 ;
  assign n1316 = n1309 | n1315 ;
  assign n1317 = n1309 & n1315 ;
  assign n1318 = n1316 & ~n1317 ;
  assign n1319 = n323 | n324 ;
  assign n1320 = ~n468 & n1319 ;
  assign n1321 = n468 & ~n1319 ;
  assign n1322 = n1320 | n1321 ;
  assign n1323 = n328 | n329 ;
  assign n1324 = ~n346 & n466 ;
  assign n1325 = n340 | n1324 ;
  assign n1326 = n1323 | n1325 ;
  assign n1327 = n1323 & n1325 ;
  assign n1328 = n1326 & ~n1327 ;
  assign n1329 = n338 | n466 ;
  assign n1330 = ~n344 & n1329 ;
  assign n1331 = n343 & ~n1330 ;
  assign n1332 = ~n343 & n1330 ;
  assign n1333 = n1331 | n1332 ;
  assign n1334 = ~n345 & n466 ;
  assign n1335 = n345 & ~n466 ;
  assign n1336 = n1334 | n1335 ;
  assign n1337 = N242 & ~N5 ;
  assign n1338 = N134 & ~N5 ;
  assign n1339 = N133 & n1338 ;
  assign n1340 = n311 & n312 ;
  assign n1341 = n313 & ~n1340 ;
  assign n1342 = n308 & n1341 ;
  assign n1343 = n308 | n1341 ;
  assign n1344 = ~n1342 & n1343 ;
  assign n1345 = n317 & ~n1344 ;
  assign n1346 = ~n306 & n1208 ;
  assign n1347 = ~n297 & n310 ;
  assign n1348 = n302 | n310 ;
  assign n1349 = ~n1347 & n1348 ;
  assign n1350 = n1207 & ~n1349 ;
  assign n1351 = ~n1207 & n1349 ;
  assign n1352 = n1350 | n1351 ;
  assign n1353 = n1346 & ~n1352 ;
  assign n1354 = ~n1346 & n1352 ;
  assign n1355 = n1353 | n1354 ;
  assign n1356 = n1345 | n1355 ;
  assign n1357 = n1345 & n1355 ;
  assign n1358 = n1356 & ~n1357 ;
  assign n1359 = n470 & ~n1358 ;
  assign n1360 = n297 | n301 ;
  assign n1361 = ~n303 & n1360 ;
  assign n1362 = n1207 & n1361 ;
  assign n1363 = n1207 | n1361 ;
  assign n1364 = ~n1362 & n1363 ;
  assign n1365 = n306 | n1364 ;
  assign n1366 = n306 & n1364 ;
  assign n1367 = n1365 & ~n1366 ;
  assign n1368 = n1344 & n1367 ;
  assign n1369 = n1344 | n1367 ;
  assign n1370 = ~n1368 & n1369 ;
  assign n1371 = ~n470 & n1370 ;
  assign n1372 = n1359 | n1371 ;
  assign n1373 = n314 & n315 ;
  assign n1374 = n316 & ~n1373 ;
  assign n1375 = n1372 & ~n1374 ;
  assign n1376 = ~n1372 & n1374 ;
  assign n1377 = n1375 | n1376 ;
  assign n1378 = n261 | n271 ;
  assign n1379 = ~n272 & n1378 ;
  assign n1380 = n266 & ~n275 ;
  assign n1381 = n274 & ~n1275 ;
  assign n1382 = n1380 | n1381 ;
  assign n1383 = ~n277 & n1266 ;
  assign n1384 = n277 & ~n1266 ;
  assign n1385 = n1383 | n1384 ;
  assign n1386 = n1382 | n1385 ;
  assign n1387 = n1382 & n1385 ;
  assign n1388 = n1386 & ~n1387 ;
  assign n1389 = ~n1379 & n1388 ;
  assign n1390 = n1379 & ~n1388 ;
  assign n1391 = n1389 | n1390 ;
  assign n1392 = n472 & ~n1391 ;
  assign n1393 = n266 & n274 ;
  assign n1394 = n275 & ~n1393 ;
  assign n1395 = ~n277 & n1394 ;
  assign n1396 = n277 & ~n1394 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = n1275 | n1281 ;
  assign n1399 = ~n276 & n1398 ;
  assign n1400 = n1266 & n1399 ;
  assign n1401 = n1266 | n1399 ;
  assign n1402 = ~n1400 & n1401 ;
  assign n1403 = n279 | n1402 ;
  assign n1404 = n279 & n1402 ;
  assign n1405 = n1403 & ~n1404 ;
  assign n1406 = n1397 & n1405 ;
  assign n1407 = n1397 | n1405 ;
  assign n1408 = ~n1406 & n1407 ;
  assign n1409 = ~n472 & n1408 ;
  assign n1410 = n1392 | n1409 ;
  assign n1411 = n1377 & ~n1410 ;
  assign n1412 = ~n1377 & n1410 ;
  assign n1413 = n1411 | n1412 ;
  assign n1414 = n222 & n485 ;
  assign n1415 = n221 | n1414 ;
  assign n1416 = ~n250 & n477 ;
  assign n1417 = n250 & ~n477 ;
  assign n1418 = n1416 | n1417 ;
  assign n1419 = ~n216 & n1418 ;
  assign n1420 = n216 & ~n1418 ;
  assign n1421 = n1419 | n1420 ;
  assign n1422 = n479 | n480 ;
  assign n1423 = ~n481 & n1422 ;
  assign n1424 = n1229 & ~n1423 ;
  assign n1425 = ~n1229 & n1423 ;
  assign n1426 = n1424 | n1425 ;
  assign n1427 = n250 & n482 ;
  assign n1428 = n1426 & ~n1427 ;
  assign n1429 = n248 & ~n482 ;
  assign n1430 = n240 | n478 ;
  assign n1431 = n244 & n478 ;
  assign n1432 = n1430 & ~n1431 ;
  assign n1433 = n251 & n1432 ;
  assign n1434 = n251 | n1432 ;
  assign n1435 = ~n1433 & n1434 ;
  assign n1436 = ~n1429 & n1435 ;
  assign n1437 = n1429 & ~n1435 ;
  assign n1438 = n1436 | n1437 ;
  assign n1439 = n1428 & ~n1438 ;
  assign n1440 = ~n1428 & n1438 ;
  assign n1441 = n1439 | n1440 ;
  assign n1442 = n476 | n1441 ;
  assign n1443 = n240 | n243 ;
  assign n1444 = ~n245 & n1443 ;
  assign n1445 = ~n251 & n1444 ;
  assign n1446 = n251 & ~n1444 ;
  assign n1447 = n1445 | n1446 ;
  assign n1448 = n248 | n1447 ;
  assign n1449 = n248 & n1447 ;
  assign n1450 = n1448 & ~n1449 ;
  assign n1451 = n1426 & n1450 ;
  assign n1452 = n1426 | n1450 ;
  assign n1453 = ~n1451 & n1452 ;
  assign n1454 = n476 & n1453 ;
  assign n1455 = n1442 & ~n1454 ;
  assign n1456 = ~n1421 & n1455 ;
  assign n1457 = n1421 & ~n1455 ;
  assign n1458 = n1456 | n1457 ;
  assign n1459 = n1415 | n1458 ;
  assign n1460 = n1415 & n1458 ;
  assign n1461 = n1459 & ~n1460 ;
  assign n1462 = n334 & n338 ;
  assign n1463 = n339 & ~n1462 ;
  assign n1464 = ~n343 & n344 ;
  assign n1465 = n1463 | n1464 ;
  assign n1466 = ~n1319 & n1323 ;
  assign n1467 = n1319 & ~n1323 ;
  assign n1468 = n1466 | n1467 ;
  assign n1469 = n1465 & ~n1468 ;
  assign n1470 = ~n1465 & n1468 ;
  assign n1471 = n1469 | n1470 ;
  assign n1472 = n348 & n1471 ;
  assign n1473 = n348 | n1471 ;
  assign n1474 = ~n1472 & n1473 ;
  assign n1475 = n466 & ~n1474 ;
  assign n1476 = n328 | n340 ;
  assign n1477 = ~n329 & n1476 ;
  assign n1478 = n343 & ~n1477 ;
  assign n1479 = ~n343 & n1477 ;
  assign n1480 = n1478 | n1479 ;
  assign n1481 = n340 & ~n344 ;
  assign n1482 = ~n334 & n344 ;
  assign n1483 = n1481 | n1482 ;
  assign n1484 = n1319 & ~n1483 ;
  assign n1485 = ~n1319 & n1483 ;
  assign n1486 = n1484 | n1485 ;
  assign n1487 = n1480 | n1486 ;
  assign n1488 = n1480 & n1486 ;
  assign n1489 = n1487 & ~n1488 ;
  assign n1490 = n466 | n1489 ;
  assign n1491 = ~n1475 & n1490 ;
  assign n1492 = n372 | n459 ;
  assign n1493 = ~n460 & n1492 ;
  assign n1494 = n358 | n1309 ;
  assign n1495 = n358 & n1309 ;
  assign n1496 = n1494 & ~n1495 ;
  assign n1497 = n1493 & n1496 ;
  assign n1498 = n1493 | n1496 ;
  assign n1499 = ~n1497 & n1498 ;
  assign n1500 = n1300 | n1499 ;
  assign n1501 = n1300 & n1499 ;
  assign n1502 = n1500 & ~n1501 ;
  assign n1503 = n456 | n1502 ;
  assign n1504 = n375 & n1300 ;
  assign n1505 = n382 & ~n1504 ;
  assign n1506 = ~n461 & n1303 ;
  assign n1507 = n352 & ~n359 ;
  assign n1508 = ~n357 & n360 ;
  assign n1509 = n1507 | n1508 ;
  assign n1510 = n1506 | n1509 ;
  assign n1511 = n1506 & n1509 ;
  assign n1512 = n1510 & ~n1511 ;
  assign n1513 = n1505 & ~n1512 ;
  assign n1514 = ~n1505 & n1512 ;
  assign n1515 = n1513 | n1514 ;
  assign n1516 = n456 & n1515 ;
  assign n1517 = n1503 & ~n1516 ;
  assign n1518 = n367 & n373 ;
  assign n1519 = n374 & ~n1518 ;
  assign n1520 = n1517 & ~n1519 ;
  assign n1521 = ~n1517 & n1519 ;
  assign n1522 = n1520 | n1521 ;
  assign n1523 = ~n1491 & n1522 ;
  assign n1524 = n1491 & ~n1522 ;
  assign n1525 = n1523 | n1524 ;
  assign n1526 = n403 | n448 ;
  assign n1527 = n397 & n448 ;
  assign n1528 = n1526 & ~n1527 ;
  assign n1529 = n405 | n1528 ;
  assign n1530 = n405 & n1528 ;
  assign n1531 = n1529 & ~n1530 ;
  assign n1532 = n451 & n452 ;
  assign n1533 = n453 & ~n1532 ;
  assign n1534 = n447 & ~n1533 ;
  assign n1535 = ~n447 & n1533 ;
  assign n1536 = n1534 | n1535 ;
  assign n1537 = n1531 & n1536 ;
  assign n1538 = n1531 | n1536 ;
  assign n1539 = ~n1537 & n1538 ;
  assign n1540 = n445 & ~n1539 ;
  assign n1541 = n396 & ~n401 ;
  assign n1542 = n397 & n401 ;
  assign n1543 = n1541 | n1542 ;
  assign n1544 = n450 & ~n1543 ;
  assign n1545 = n405 & n1544 ;
  assign n1546 = n831 & ~n1544 ;
  assign n1547 = ~n405 & n1546 ;
  assign n1548 = n1545 | n1547 ;
  assign n1549 = ~n1533 & n1548 ;
  assign n1550 = n1533 & ~n1548 ;
  assign n1551 = n1549 | n1550 ;
  assign n1552 = n445 | n1551 ;
  assign n1553 = N367 & n1552 ;
  assign n1554 = ~n1540 & n1553 ;
  assign n1555 = ~n436 & n1539 ;
  assign n1556 = ~N367 & n435 ;
  assign n1557 = n1551 & n1556 ;
  assign n1558 = n1555 | n1557 ;
  assign n1559 = n1554 | n1558 ;
  assign n1560 = ~n416 & n431 ;
  assign n1561 = n432 & ~n1560 ;
  assign n1562 = ~n426 & n821 ;
  assign n1563 = n212 & n438 ;
  assign n1564 = n439 & ~n1563 ;
  assign n1565 = n810 & n1564 ;
  assign n1566 = n810 | n1564 ;
  assign n1567 = ~n1565 & n1566 ;
  assign n1568 = ~n1562 & n1567 ;
  assign n1569 = n1562 & ~n1567 ;
  assign n1570 = n1568 | n1569 ;
  assign n1571 = n1561 & ~n1570 ;
  assign n1572 = ~n1561 & n1570 ;
  assign n1573 = N367 | n1572 ;
  assign n1574 = n1571 | n1573 ;
  assign n1575 = ~n431 & n440 ;
  assign n1576 = n211 | n425 ;
  assign n1577 = n426 | n428 ;
  assign n1578 = n211 & ~n1577 ;
  assign n1579 = n1576 & ~n1578 ;
  assign n1580 = ~n1575 & n1579 ;
  assign n1581 = n1575 & ~n1579 ;
  assign n1582 = n1580 | n1581 ;
  assign n1583 = n443 & ~n1567 ;
  assign n1584 = ~n443 & n1567 ;
  assign n1585 = n1583 | n1584 ;
  assign n1586 = n1582 & n1585 ;
  assign n1587 = n1582 | n1585 ;
  assign n1588 = N367 & n1587 ;
  assign n1589 = ~n1586 & n1588 ;
  assign n1590 = n1574 & ~n1589 ;
  assign n1591 = n437 & n441 ;
  assign n1592 = n437 | n441 ;
  assign n1593 = ~n1591 & n1592 ;
  assign n1594 = n1590 | n1593 ;
  assign n1595 = n1590 & n1593 ;
  assign n1596 = n1594 & ~n1595 ;
  assign n1597 = n1559 | n1596 ;
  assign n1598 = n1559 & n1596 ;
  assign n1599 = n1597 & ~n1598 ;
  assign n1600 = N1 & N163 ;
  assign n1601 = N5 | N57 ;
  assign N10025 = ~n215 ;
  assign N10101 = ~n488 ;
  assign N10102 = n809 ;
  assign N10103 = n809 ;
  assign N10104 = ~n488 ;
  assign N10109 = ~n816 ;
  assign N10110 = ~n820 ;
  assign N10111 = ~n826 ;
  assign N10112 = ~n830 ;
  assign N10350 = ~n836 ;
  assign N10351 = ~n842 ;
  assign N10352 = ~n846 ;
  assign N10353 = ~n849 ;
  assign N10574 = ~n965 ;
  assign N10575 = ~n1088 ;
  assign N10576 = ~n1200 ;
  assign N10628 = n809 ;
  assign N10632 = ~n1203 ;
  assign N10641 = ~n1206 ;
  assign N10704 = n661 ;
  assign N10706 = ~n488 ;
  assign N10711 = n1214 ;
  assign N10712 = ~n1218 ;
  assign N10713 = ~n1223 ;
  assign N10714 = ~n1227 ;
  assign N10715 = ~n1234 ;
  assign N10716 = ~n1238 ;
  assign N10717 = ~n1243 ;
  assign N10718 = ~n1247 ;
  assign N10729 = ~n1265 ;
  assign N10759 = ~n488 ;
  assign N10760 = ~n1269 ;
  assign N10761 = ~n1274 ;
  assign N10762 = ~n1280 ;
  assign N10763 = ~n1284 ;
  assign N10827 = ~n1288 ;
  assign N10837 = n1294 ;
  assign N10838 = n1294 ;
  assign N10839 = n1296 ;
  assign N10840 = n1296 ;
  assign N10868 = ~n1302 ;
  assign N10869 = ~n1308 ;
  assign N10870 = ~n1314 ;
  assign N10871 = ~n1318 ;
  assign N10905 = ~n1322 ;
  assign N10906 = ~n1328 ;
  assign N10907 = ~n1333 ;
  assign N10908 = ~n1336 ;
  assign N1110 = ~n1337 ;
  assign N1111 = ~N15 ;
  assign N1112 = ~n1337 ;
  assign N1113 = ~n1339 ;
  assign N1114 = ~N15 ;
  assign N11333 = ~n1413 ;
  assign N11334 = n1461 ;
  assign N11340 = n1525 ;
  assign N11342 = n1599 ;
  assign N1489 = ~n1339 ;
  assign N1490 = N1 ;
  assign N1781 = n1600 ;
  assign N241_O = N241_I ;
  assign N387 = N1 ;
  assign N388 = N1 ;
  assign N478 = N248 ;
  assign N482 = N254 ;
  assign N484 = N257 ;
  assign N486 = N260 ;
  assign N489 = N263 ;
  assign N492 = N267 ;
  assign N501 = N274 ;
  assign N505 = N280 ;
  assign N507 = N283 ;
  assign N509 = N286 ;
  assign N511 = N289 ;
  assign N513 = N293 ;
  assign N515 = N296 ;
  assign N517 = N299 ;
  assign N519 = N303 ;
  assign N535 = N307 ;
  assign N537 = N310 ;
  assign N539 = N313 ;
  assign N541 = N316 ;
  assign N543 = N319 ;
  assign N545 = N322 ;
  assign N547 = N325 ;
  assign N549 = N328 ;
  assign N551 = N331 ;
  assign N553 = N334 ;
  assign N556 = N337 ;
  assign N559 = N343 ;
  assign N561 = N346 ;
  assign N563 = N349 ;
  assign N565 = N352 ;
  assign N567 = N355 ;
  assign N569 = N358 ;
  assign N571 = N361 ;
  assign N573 = N364 ;
  assign N582 = ~N15 ;
  assign N643 = N251 ;
  assign N707 = N277 ;
  assign N813 = N340 ;
  assign N881 = n1601 ;
  assign N882 = ~n1250 ;
  assign N883 = ~n1253 ;
  assign N884 = ~n1257 ;
  assign N885 = ~n1260 ;
  assign N889 = N1 ;
  assign N945 = N106 ;
endmodule
