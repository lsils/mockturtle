module top( b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ , s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ );
  input b_4_ , a_1_ , a_2_ , b_1_ , b_7_ , a_6_ , a_4_ , b_2_ , a_7_ , a_5_ , b_5_ , b_3_ , b_6_ , b_0_ , a_3_ , a_0_ ;
  output s_1_ , s_8_ , s_3_ , s_5_ , s_9_ , s_2_ , s_11_ , s_15_ , s_4_ , s_10_ , s_14_ , s_7_ , s_13_ , s_12_ , s_6_ , s_0_ ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 ;
  assign n17 = a_1_ & b_0_ ;
  assign n18 = b_1_ & a_0_ ;
  assign n19 = n17 & n18 ;
  assign n20 = n17 | n18 ;
  assign n21 = ~n19 & n20 ;
  assign n22 = a_1_ & b_6_ ;
  assign n23 = b_4_ & a_2_ ;
  assign n24 = b_3_ & a_3_ ;
  assign n25 = n23 & n24 ;
  assign n26 = a_1_ & b_5_ ;
  assign n27 = n23 | n24 ;
  assign n28 = ~n25 & n27 ;
  assign n29 = n26 & n28 ;
  assign n30 = n25 | n29 ;
  assign n31 = n22 & n30 ;
  assign n32 = b_7_ & a_0_ ;
  assign n33 = n22 | n30 ;
  assign n34 = ~n31 & n33 ;
  assign n35 = n32 & n34 ;
  assign n36 = n31 | n35 ;
  assign n37 = a_1_ & b_7_ ;
  assign n38 = a_2_ & b_6_ ;
  assign n39 = b_4_ & a_3_ ;
  assign n40 = a_4_ & b_3_ ;
  assign n41 = n39 & n40 ;
  assign n42 = n39 | n40 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = a_2_ & b_5_ ;
  assign n45 = n43 & n44 ;
  assign n46 = n41 | n45 ;
  assign n47 = n38 & n46 ;
  assign n48 = n38 | n46 ;
  assign n49 = ~n47 & n48 ;
  assign n50 = n37 & n49 ;
  assign n51 = n37 | n49 ;
  assign n52 = ~n50 & n51 ;
  assign n53 = b_5_ & a_3_ ;
  assign n54 = b_4_ & a_4_ ;
  assign n55 = a_5_ & b_3_ ;
  assign n56 = n54 & n55 ;
  assign n57 = n54 | n55 ;
  assign n58 = ~n56 & n57 ;
  assign n59 = n53 & n58 ;
  assign n60 = n53 | n58 ;
  assign n61 = ~n59 & n60 ;
  assign n62 = b_1_ & a_6_ ;
  assign n63 = a_7_ & b_0_ ;
  assign n64 = n62 & n63 ;
  assign n65 = b_2_ & a_5_ ;
  assign n66 = n62 | n63 ;
  assign n67 = ~n64 & n66 ;
  assign n68 = n65 & n67 ;
  assign n69 = n64 | n68 ;
  assign n70 = b_1_ & a_7_ ;
  assign n71 = a_6_ & b_2_ ;
  assign n72 = n70 | n71 ;
  assign n73 = b_2_ & a_7_ ;
  assign n74 = n62 & n73 ;
  assign n75 = n72 & ~n74 ;
  assign n76 = n69 & n75 ;
  assign n77 = n69 | n75 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = n61 & n78 ;
  assign n80 = n61 | n78 ;
  assign n81 = ~n79 & n80 ;
  assign n82 = n65 | n67 ;
  assign n83 = ~n68 & n82 ;
  assign n84 = a_5_ & b_0_ ;
  assign n85 = n62 & n84 ;
  assign n86 = a_4_ & b_2_ ;
  assign n87 = b_1_ & a_5_ ;
  assign n88 = a_6_ & b_0_ ;
  assign n89 = n87 | n88 ;
  assign n90 = ~n85 & n89 ;
  assign n91 = n86 & n90 ;
  assign n92 = n85 | n91 ;
  assign n93 = n83 & n92 ;
  assign n94 = n43 | n44 ;
  assign n95 = ~n45 & n94 ;
  assign n96 = n83 | n92 ;
  assign n97 = ~n93 & n96 ;
  assign n98 = n95 & n97 ;
  assign n99 = n93 | n98 ;
  assign n100 = n81 & n99 ;
  assign n101 = n81 | n99 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = n52 & n102 ;
  assign n104 = n52 | n102 ;
  assign n105 = ~n103 & n104 ;
  assign n106 = n95 | n97 ;
  assign n107 = ~n98 & n106 ;
  assign n108 = n86 | n90 ;
  assign n109 = ~n91 & n108 ;
  assign n110 = b_1_ & a_4_ ;
  assign n111 = n84 & n110 ;
  assign n112 = b_2_ & a_3_ ;
  assign n113 = n84 | n110 ;
  assign n114 = ~n111 & n113 ;
  assign n115 = n112 & n114 ;
  assign n116 = n111 | n115 ;
  assign n117 = n109 & n116 ;
  assign n118 = n26 | n28 ;
  assign n119 = ~n29 & n118 ;
  assign n120 = n109 | n116 ;
  assign n121 = ~n117 & n120 ;
  assign n122 = n119 & n121 ;
  assign n123 = n117 | n122 ;
  assign n124 = n107 & n123 ;
  assign n125 = n32 | n34 ;
  assign n126 = ~n35 & n125 ;
  assign n127 = n107 | n123 ;
  assign n128 = ~n124 & n127 ;
  assign n129 = n126 & n128 ;
  assign n130 = n124 | n129 ;
  assign n131 = n105 & n130 ;
  assign n132 = n105 | n130 ;
  assign n133 = ~n131 & n132 ;
  assign n134 = n36 & n133 ;
  assign n135 = n36 | n133 ;
  assign n136 = ~n134 & n135 ;
  assign n137 = n126 | n128 ;
  assign n138 = ~n129 & n137 ;
  assign n139 = n119 | n121 ;
  assign n140 = ~n122 & n139 ;
  assign n141 = n112 | n114 ;
  assign n142 = ~n115 & n141 ;
  assign n143 = a_4_ & b_0_ ;
  assign n144 = b_1_ & a_3_ ;
  assign n145 = n143 & n144 ;
  assign n146 = a_2_ & b_2_ ;
  assign n147 = n143 | n144 ;
  assign n148 = ~n145 & n147 ;
  assign n149 = n146 & n148 ;
  assign n150 = n145 | n149 ;
  assign n151 = n142 & n150 ;
  assign n152 = b_5_ & a_0_ ;
  assign n153 = b_4_ & a_1_ ;
  assign n154 = a_2_ & b_3_ ;
  assign n155 = n153 | n154 ;
  assign n156 = n153 & n154 ;
  assign n157 = n155 & ~n156 ;
  assign n158 = n152 & n157 ;
  assign n159 = n152 | n157 ;
  assign n160 = ~n158 & n159 ;
  assign n161 = n142 | n150 ;
  assign n162 = ~n151 & n161 ;
  assign n163 = n160 & n162 ;
  assign n164 = n151 | n163 ;
  assign n165 = n140 & n164 ;
  assign n166 = b_6_ & a_0_ ;
  assign n167 = n156 | n158 ;
  assign n168 = n166 & n167 ;
  assign n169 = n166 | n167 ;
  assign n170 = ~n168 & n169 ;
  assign n171 = n140 | n164 ;
  assign n172 = ~n165 & n171 ;
  assign n173 = n170 & n172 ;
  assign n174 = n165 | n173 ;
  assign n175 = n138 & n174 ;
  assign n176 = n138 | n174 ;
  assign n177 = ~n175 & n176 ;
  assign n178 = n168 & n177 ;
  assign n179 = n175 | n178 ;
  assign n180 = n136 | n179 ;
  assign n181 = n136 & n179 ;
  assign n182 = n180 & ~n181 ;
  assign n183 = n168 | n177 ;
  assign n184 = ~n178 & n183 ;
  assign n185 = n170 | n172 ;
  assign n186 = ~n173 & n185 ;
  assign n187 = n160 | n162 ;
  assign n188 = ~n163 & n187 ;
  assign n189 = n146 | n148 ;
  assign n190 = ~n149 & n189 ;
  assign n191 = a_2_ & b_1_ ;
  assign n192 = b_0_ & a_3_ ;
  assign n193 = n191 & n192 ;
  assign n194 = a_1_ & b_2_ ;
  assign n195 = n191 | n192 ;
  assign n196 = ~n193 & n195 ;
  assign n197 = n194 & n196 ;
  assign n198 = n193 | n197 ;
  assign n199 = n190 & n198 ;
  assign n200 = a_1_ & b_3_ ;
  assign n201 = b_4_ & a_0_ ;
  assign n202 = n200 | n201 ;
  assign n203 = b_3_ & a_0_ ;
  assign n204 = n153 & n203 ;
  assign n205 = n202 & ~n204 ;
  assign n206 = n190 | n198 ;
  assign n207 = ~n199 & n206 ;
  assign n208 = n205 & n207 ;
  assign n209 = n199 | n208 ;
  assign n210 = n188 & n209 ;
  assign n211 = n188 | n209 ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n204 & n212 ;
  assign n214 = n210 | n213 ;
  assign n215 = n186 & n214 ;
  assign n216 = n184 & n215 ;
  assign n217 = n184 | n215 ;
  assign n218 = ~n216 & n217 ;
  assign n219 = n186 | n214 ;
  assign n220 = ~n215 & n219 ;
  assign n221 = n204 | n212 ;
  assign n222 = ~n213 & n221 ;
  assign n223 = n205 | n207 ;
  assign n224 = ~n208 & n223 ;
  assign n225 = a_1_ & b_1_ ;
  assign n226 = a_2_ & b_0_ ;
  assign n227 = n225 & n226 ;
  assign n228 = b_2_ & a_0_ ;
  assign n229 = n225 | n226 ;
  assign n230 = ~n227 & n229 ;
  assign n231 = n228 & n230 ;
  assign n232 = n227 | n231 ;
  assign n233 = n194 | n196 ;
  assign n234 = ~n197 & n233 ;
  assign n235 = n232 & n234 ;
  assign n236 = n232 | n234 ;
  assign n237 = ~n235 & n236 ;
  assign n238 = n203 & n237 ;
  assign n239 = n235 | n238 ;
  assign n240 = n224 & n239 ;
  assign n241 = n222 & n240 ;
  assign n242 = n220 & n241 ;
  assign n243 = n220 | n241 ;
  assign n244 = ~n242 & n243 ;
  assign n245 = n222 | n240 ;
  assign n246 = ~n241 & n245 ;
  assign n247 = n224 | n239 ;
  assign n248 = ~n240 & n247 ;
  assign n249 = n228 | n230 ;
  assign n250 = ~n231 & n249 ;
  assign n251 = n19 & n250 ;
  assign n252 = n203 | n237 ;
  assign n253 = ~n238 & n252 ;
  assign n254 = n251 & n253 ;
  assign n255 = n248 & n254 ;
  assign n256 = n246 & n255 ;
  assign n257 = n244 & n256 ;
  assign n258 = n242 | n257 ;
  assign n259 = n218 & n258 ;
  assign n260 = n216 | n259 ;
  assign n261 = n182 & n260 ;
  assign n262 = n182 | n260 ;
  assign n263 = ~n261 & n262 ;
  assign n264 = n251 | n253 ;
  assign n265 = ~n254 & n264 ;
  assign n266 = n246 | n255 ;
  assign n267 = ~n256 & n266 ;
  assign n268 = n181 | n261 ;
  assign n269 = n131 | n134 ;
  assign n270 = n47 | n50 ;
  assign n271 = a_2_ & b_7_ ;
  assign n272 = b_6_ & a_3_ ;
  assign n273 = n56 | n59 ;
  assign n274 = n272 & n273 ;
  assign n275 = n272 | n273 ;
  assign n276 = ~n274 & n275 ;
  assign n277 = n271 & n276 ;
  assign n278 = n271 | n276 ;
  assign n279 = ~n277 & n278 ;
  assign n280 = a_4_ & b_5_ ;
  assign n281 = b_4_ & a_5_ ;
  assign n282 = a_6_ & b_3_ ;
  assign n283 = n281 | n282 ;
  assign n284 = b_4_ & a_6_ ;
  assign n285 = n55 & n284 ;
  assign n286 = n283 & ~n285 ;
  assign n287 = n280 & n286 ;
  assign n288 = n280 | n286 ;
  assign n289 = ~n287 & n288 ;
  assign n290 = ~n62 & n73 ;
  assign n291 = n289 & n290 ;
  assign n292 = n289 | n290 ;
  assign n293 = ~n291 & n292 ;
  assign n294 = n76 | n79 ;
  assign n295 = n293 & n294 ;
  assign n296 = n293 | n294 ;
  assign n297 = ~n295 & n296 ;
  assign n298 = n279 & n297 ;
  assign n299 = n279 | n297 ;
  assign n300 = ~n298 & n299 ;
  assign n301 = n100 | n103 ;
  assign n302 = n300 & n301 ;
  assign n303 = n300 | n301 ;
  assign n304 = ~n302 & n303 ;
  assign n305 = n270 & n304 ;
  assign n306 = n270 | n304 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = n269 & n307 ;
  assign n309 = n269 | n307 ;
  assign n310 = ~n308 & n309 ;
  assign n311 = n268 | n310 ;
  assign n312 = n268 & n310 ;
  assign n313 = n311 & ~n312 ;
  assign n314 = n19 | n250 ;
  assign n315 = ~n251 & n314 ;
  assign n316 = n285 | n287 ;
  assign n317 = a_4_ & b_6_ ;
  assign n318 = n316 & n317 ;
  assign n319 = b_7_ & a_3_ ;
  assign n320 = n316 | n317 ;
  assign n321 = ~n318 & n320 ;
  assign n322 = n319 & n321 ;
  assign n323 = n318 | n322 ;
  assign n324 = a_7_ & b_5_ ;
  assign n325 = n284 & n324 ;
  assign n326 = b_4_ & a_7_ ;
  assign n327 = a_6_ & b_5_ ;
  assign n328 = n326 | n327 ;
  assign n329 = ~n325 & n328 ;
  assign n330 = b_7_ & a_4_ ;
  assign n331 = n282 & n326 ;
  assign n332 = a_5_ & b_5_ ;
  assign n333 = a_7_ & b_3_ ;
  assign n334 = n284 | n333 ;
  assign n335 = ~n331 & n334 ;
  assign n336 = n332 & n335 ;
  assign n337 = n331 | n336 ;
  assign n338 = a_5_ & b_6_ ;
  assign n339 = n337 & n338 ;
  assign n340 = n337 | n338 ;
  assign n341 = ~n339 & n340 ;
  assign n342 = n330 & n341 ;
  assign n343 = n330 | n341 ;
  assign n344 = ~n342 & n343 ;
  assign n345 = n329 & n344 ;
  assign n346 = n329 | n344 ;
  assign n347 = ~n345 & n346 ;
  assign n348 = n74 | n291 ;
  assign n349 = n332 | n335 ;
  assign n350 = ~n336 & n349 ;
  assign n351 = n348 & n350 ;
  assign n352 = n348 | n350 ;
  assign n353 = ~n351 & n352 ;
  assign n354 = n319 | n321 ;
  assign n355 = ~n322 & n354 ;
  assign n356 = n353 & n355 ;
  assign n357 = n351 | n356 ;
  assign n358 = n347 & n357 ;
  assign n359 = n347 | n357 ;
  assign n360 = ~n358 & n359 ;
  assign n361 = n323 & n360 ;
  assign n362 = n323 | n360 ;
  assign n363 = ~n361 & n362 ;
  assign n364 = n295 | n298 ;
  assign n365 = n353 | n355 ;
  assign n366 = ~n356 & n365 ;
  assign n367 = n364 & n366 ;
  assign n368 = n274 | n277 ;
  assign n369 = n364 | n366 ;
  assign n370 = ~n367 & n369 ;
  assign n371 = n368 & n370 ;
  assign n372 = n367 | n371 ;
  assign n373 = n363 & n372 ;
  assign n374 = n363 | n372 ;
  assign n375 = ~n373 & n374 ;
  assign n376 = n302 | n305 ;
  assign n377 = n368 | n370 ;
  assign n378 = ~n371 & n377 ;
  assign n379 = n376 & n378 ;
  assign n380 = n268 | n308 ;
  assign n381 = n309 & n380 ;
  assign n382 = n376 | n378 ;
  assign n383 = ~n379 & n382 ;
  assign n384 = n381 & n383 ;
  assign n385 = n379 | n384 ;
  assign n386 = n375 | n385 ;
  assign n387 = n375 & n385 ;
  assign n388 = n386 & ~n387 ;
  assign n389 = a_6_ & b_6_ ;
  assign n390 = b_7_ & a_7_ ;
  assign n391 = n389 & n390 ;
  assign n392 = ~n389 & n390 ;
  assign n393 = a_7_ & b_6_ ;
  assign n394 = b_7_ & a_6_ ;
  assign n395 = n393 | n394 ;
  assign n396 = ~n391 & n395 ;
  assign n397 = b_7_ & a_5_ ;
  assign n398 = b_6_ & n325 ;
  assign n399 = n325 | n389 ;
  assign n400 = ~n398 & n399 ;
  assign n401 = n397 & n400 ;
  assign n402 = n397 | n400 ;
  assign n403 = ~n401 & n402 ;
  assign n404 = n324 & n403 ;
  assign n405 = n396 & n404 ;
  assign n406 = n398 | n401 ;
  assign n407 = n396 | n404 ;
  assign n408 = ~n405 & n407 ;
  assign n409 = n406 & n408 ;
  assign n410 = n405 | n409 ;
  assign n411 = n392 & n410 ;
  assign n412 = n391 | n411 ;
  assign n413 = n392 | n410 ;
  assign n414 = ~n411 & n413 ;
  assign n415 = n406 | n408 ;
  assign n416 = ~n409 & n415 ;
  assign n417 = n324 | n403 ;
  assign n418 = ~n404 & n417 ;
  assign n419 = n345 & n418 ;
  assign n420 = n339 | n342 ;
  assign n421 = n345 | n418 ;
  assign n422 = ~n419 & n421 ;
  assign n423 = n420 & n422 ;
  assign n424 = n419 | n423 ;
  assign n425 = n416 & n424 ;
  assign n426 = n416 | n424 ;
  assign n427 = ~n425 & n426 ;
  assign n428 = n420 | n422 ;
  assign n429 = ~n423 & n428 ;
  assign n430 = n358 | n361 ;
  assign n431 = n429 & n430 ;
  assign n432 = n429 | n430 ;
  assign n433 = ~n431 & n432 ;
  assign n434 = n373 | n387 ;
  assign n435 = n433 & n434 ;
  assign n436 = n431 | n435 ;
  assign n437 = n427 & n436 ;
  assign n438 = n425 | n437 ;
  assign n439 = n414 & n438 ;
  assign n440 = n412 | n439 ;
  assign n441 = n248 | n254 ;
  assign n442 = ~n255 & n441 ;
  assign n443 = n381 | n383 ;
  assign n444 = ~n384 & n443 ;
  assign n445 = n414 | n438 ;
  assign n446 = ~n439 & n445 ;
  assign n447 = n218 | n258 ;
  assign n448 = ~n259 & n447 ;
  assign n449 = n427 | n436 ;
  assign n450 = ~n437 & n449 ;
  assign n451 = n433 | n434 ;
  assign n452 = ~n435 & n451 ;
  assign n453 = n244 | n256 ;
  assign n454 = ~n257 & n453 ;
  assign n455 = b_0_ & a_0_ ;
  assign s_1_ = n21 ;
  assign s_8_ = n263 ;
  assign s_3_ = n265 ;
  assign s_5_ = n267 ;
  assign s_9_ = n313 ;
  assign s_2_ = n315 ;
  assign s_11_ = n388 ;
  assign s_15_ = n440 ;
  assign s_4_ = n442 ;
  assign s_10_ = n444 ;
  assign s_14_ = n446 ;
  assign s_7_ = n448 ;
  assign s_13_ = n450 ;
  assign s_12_ = n452 ;
  assign s_6_ = n454 ;
  assign s_0_ = n455 ;
endmodule
