module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 ;
  assign n15 = x8 | x10 ;
  assign n16 = x10 & ~x11 ;
  assign n17 = x8 & x9 ;
  assign n18 = n16 & ~n17 ;
  assign n19 = ~x8 & x13 ;
  assign n20 = ( x9 & n16 ) | ( x9 & n19 ) | ( n16 & n19 ) ;
  assign n21 = ~n16 & n20 ;
  assign n22 = x8 & x10 ;
  assign n23 = ~x13 & n22 ;
  assign n24 = ( x9 & x11 ) | ( x9 & n23 ) | ( x11 & n23 ) ;
  assign n25 = ~x9 & n24 ;
  assign n26 = n21 | n25 ;
  assign n27 = ( n16 & ~n18 ) | ( n16 & n26 ) | ( ~n18 & n26 ) ;
  assign n28 = ~x4 & n27 ;
  assign n29 = x9 & ~x11 ;
  assign n30 = x13 | n15 ;
  assign n31 = ( x9 & ~n29 ) | ( x9 & n30 ) | ( ~n29 & n30 ) ;
  assign n32 = ~n28 & n31 ;
  assign n33 = ( x0 & ~n28 ) | ( x0 & n32 ) | ( ~n28 & n32 ) ;
  assign n34 = x0 | x4 ;
  assign n35 = ~x0 & n16 ;
  assign n36 = x4 & n35 ;
  assign n37 = ( ~x4 & n34 ) | ( ~x4 & n36 ) | ( n34 & n36 ) ;
  assign n38 = ( x9 & n19 ) | ( x9 & ~n37 ) | ( n19 & ~n37 ) ;
  assign n39 = n37 & n38 ;
  assign n40 = x8 & ~x9 ;
  assign n41 = ( ~x10 & x13 ) | ( ~x10 & n40 ) | ( x13 & n40 ) ;
  assign n42 = x10 & n41 ;
  assign n43 = ( x11 & x13 ) | ( x11 & ~n42 ) | ( x13 & ~n42 ) ;
  assign n44 = ( n41 & n42 ) | ( n41 & ~n43 ) | ( n42 & ~n43 ) ;
  assign n45 = ( ~x0 & x4 ) | ( ~x0 & n44 ) | ( x4 & n44 ) ;
  assign n46 = ( ~x8 & x9 ) | ( ~x8 & x11 ) | ( x9 & x11 ) ;
  assign n47 = ( ~x8 & x9 ) | ( ~x8 & x10 ) | ( x9 & x10 ) ;
  assign n48 = n46 & ~n47 ;
  assign n49 = ~x8 & n16 ;
  assign n50 = ~x9 & n49 ;
  assign n51 = x13 | n50 ;
  assign n52 = ( n48 & n50 ) | ( n48 & n51 ) | ( n50 & n51 ) ;
  assign n53 = ( x0 & n44 ) | ( x0 & n52 ) | ( n44 & n52 ) ;
  assign n54 = ~n45 & n53 ;
  assign n55 = ( x4 & n44 ) | ( x4 & n54 ) | ( n44 & n54 ) ;
  assign n56 = n39 | n55 ;
  assign n57 = n33 & ~n56 ;
  assign n58 = ( x4 & n15 ) | ( x4 & ~n57 ) | ( n15 & ~n57 ) ;
  assign n59 = ( x8 & x9 ) | ( x8 & ~x10 ) | ( x9 & ~x10 ) ;
  assign n60 = ( x9 & x10 ) | ( x9 & ~x11 ) | ( x10 & ~x11 ) ;
  assign n61 = n59 | n60 ;
  assign n62 = n57 | n61 ;
  assign n63 = ( n15 & ~n58 ) | ( n15 & n62 ) | ( ~n58 & n62 ) ;
  assign n64 = x10 | x11 ;
  assign n65 = ( ~x8 & x11 ) | ( ~x8 & n64 ) | ( x11 & n64 ) ;
  assign n66 = x0 & ~n57 ;
  assign n67 = n22 & n66 ;
  assign n68 = x0 & x4 ;
  assign n69 = n67 | n68 ;
  assign n70 = ( n65 & n67 ) | ( n65 & n69 ) | ( n67 & n69 ) ;
  assign n71 = ~x8 & x11 ;
  assign n72 = x4 & ~n71 ;
  assign n73 = ~x0 & n49 ;
  assign n74 = x4 | n73 ;
  assign n75 = ~n72 & n74 ;
  assign n76 = x8 | x9 ;
  assign n77 = ~x10 & n76 ;
  assign n78 = x8 & ~n64 ;
  assign n79 = ( ~x8 & n15 ) | ( ~x8 & n78 ) | ( n15 & n78 ) ;
  assign n80 = n57 & n79 ;
  assign n81 = x8 & n16 ;
  assign n82 = n80 | n81 ;
  assign n83 = ( ~x4 & n80 ) | ( ~x4 & n82 ) | ( n80 & n82 ) ;
  assign n84 = ( x0 & x4 ) | ( x0 & ~x11 ) | ( x4 & ~x11 ) ;
  assign n85 = x0 & ~n84 ;
  assign n86 = x8 & ~x10 ;
  assign n87 = ( x4 & n85 ) | ( x4 & n86 ) | ( n85 & n86 ) ;
  assign n88 = ( ~n84 & n85 ) | ( ~n84 & n87 ) | ( n85 & n87 ) ;
  assign n89 = ~x9 & n88 ;
  assign n90 = ( ~x9 & n83 ) | ( ~x9 & n89 ) | ( n83 & n89 ) ;
  assign n91 = x0 & x11 ;
  assign n92 = n90 | n91 ;
  assign n93 = ( ~n77 & n90 ) | ( ~n77 & n92 ) | ( n90 & n92 ) ;
  assign n94 = ( ~n70 & n75 ) | ( ~n70 & n93 ) | ( n75 & n93 ) ;
  assign n95 = x9 | n93 ;
  assign n96 = ( n70 & n94 ) | ( n70 & n95 ) | ( n94 & n95 ) ;
  assign n97 = ~x10 & n17 ;
  assign n98 = ~x11 & n97 ;
  assign n99 = x13 & ~n98 ;
  assign n100 = ~x9 & x10 ;
  assign n101 = n71 & n100 ;
  assign n102 = ~x13 & n101 ;
  assign n103 = ( x13 & ~n99 ) | ( x13 & n102 ) | ( ~n99 & n102 ) ;
  assign n104 = ( n63 & n96 ) | ( n63 & n103 ) | ( n96 & n103 ) ;
  assign n105 = x13 & ~n103 ;
  assign n106 = ( n63 & ~n104 ) | ( n63 & n105 ) | ( ~n104 & n105 ) ;
  assign n107 = ( x9 & x11 ) | ( x9 & ~n57 ) | ( x11 & ~n57 ) ;
  assign n108 = ~x11 & n107 ;
  assign n109 = x0 & n107 ;
  assign n110 = ( x0 & n108 ) | ( x0 & ~n109 ) | ( n108 & ~n109 ) ;
  assign n111 = ~n17 & n91 ;
  assign n112 = x9 | x11 ;
  assign n113 = x13 & n71 ;
  assign n114 = x9 & n113 ;
  assign n115 = ~x10 & n114 ;
  assign n116 = x13 & n16 ;
  assign n117 = ( n57 & n76 ) | ( n57 & ~n116 ) | ( n76 & ~n116 ) ;
  assign n118 = ( x8 & ~x9 ) | ( x8 & n66 ) | ( ~x9 & n66 ) ;
  assign n119 = ( x8 & x9 ) | ( x8 & n68 ) | ( x9 & n68 ) ;
  assign n120 = n118 & n119 ;
  assign n121 = n116 & n120 ;
  assign n122 = ( n57 & ~n117 ) | ( n57 & n121 ) | ( ~n117 & n121 ) ;
  assign n123 = ( x0 & n57 ) | ( x0 & ~n122 ) | ( n57 & ~n122 ) ;
  assign n124 = n114 | n122 ;
  assign n125 = ( x0 & ~n123 ) | ( x0 & n124 ) | ( ~n123 & n124 ) ;
  assign n126 = ~x9 & x13 ;
  assign n127 = n81 & n126 ;
  assign n128 = ~n125 & n127 ;
  assign n129 = n68 | n128 ;
  assign n130 = ( n115 & n128 ) | ( n115 & n129 ) | ( n128 & n129 ) ;
  assign n131 = x8 & n130 ;
  assign n132 = ~n112 & n131 ;
  assign n133 = ( x8 & ~x9 ) | ( x8 & x10 ) | ( ~x9 & x10 ) ;
  assign n134 = ( x10 & x11 ) | ( x10 & ~n133 ) | ( x11 & ~n133 ) ;
  assign n135 = ( ~x8 & x11 ) | ( ~x8 & n133 ) | ( x11 & n133 ) ;
  assign n136 = n134 & ~n135 ;
  assign n137 = ( ~n111 & n132 ) | ( ~n111 & n136 ) | ( n132 & n136 ) ;
  assign n138 = x10 | n136 ;
  assign n139 = ( n111 & n137 ) | ( n111 & n138 ) | ( n137 & n138 ) ;
  assign n140 = x8 | n125 ;
  assign n141 = x0 & ~n140 ;
  assign n142 = x4 | n141 ;
  assign n143 = ( n86 & n141 ) | ( n86 & n142 ) | ( n141 & n142 ) ;
  assign n144 = ( n16 & ~n17 ) | ( n16 & n125 ) | ( ~n17 & n125 ) ;
  assign n145 = x9 & ~n15 ;
  assign n146 = x11 & n130 ;
  assign n147 = n145 & n146 ;
  assign n148 = ~n125 & n147 ;
  assign n149 = ( n16 & ~n144 ) | ( n16 & n148 ) | ( ~n144 & n148 ) ;
  assign n150 = x10 & n17 ;
  assign n151 = ( ~x0 & n149 ) | ( ~x0 & n150 ) | ( n149 & n150 ) ;
  assign n152 = x11 & ~n151 ;
  assign n153 = ( x11 & n149 ) | ( x11 & ~n152 ) | ( n149 & ~n152 ) ;
  assign n154 = n112 & ~n153 ;
  assign n155 = ( n143 & n153 ) | ( n143 & ~n154 ) | ( n153 & ~n154 ) ;
  assign n156 = ( n57 & n139 ) | ( n57 & n155 ) | ( n139 & n155 ) ;
  assign n157 = x10 & ~n112 ;
  assign n158 = ( x8 & n130 ) | ( x8 & n157 ) | ( n130 & n157 ) ;
  assign n159 = ~n130 & n158 ;
  assign n160 = ( x0 & n77 ) | ( x0 & ~n159 ) | ( n77 & ~n159 ) ;
  assign n161 = x11 & n160 ;
  assign n162 = ( x11 & n159 ) | ( x11 & ~n161 ) | ( n159 & ~n161 ) ;
  assign n163 = ( ~n57 & n155 ) | ( ~n57 & n162 ) | ( n155 & n162 ) ;
  assign n164 = n156 | n163 ;
  assign n165 = n15 & ~n164 ;
  assign n166 = ( n110 & n164 ) | ( n110 & ~n165 ) | ( n164 & ~n165 ) ;
  assign n167 = ~n130 & n145 ;
  assign n168 = ( x11 & n125 ) | ( x11 & ~n167 ) | ( n125 & ~n167 ) ;
  assign n169 = ~x8 & x10 ;
  assign n170 = ( x0 & ~n112 ) | ( x0 & n169 ) | ( ~n112 & n169 ) ;
  assign n171 = ~x0 & n170 ;
  assign n172 = n125 & n171 ;
  assign n173 = ( n167 & n168 ) | ( n167 & n172 ) | ( n168 & n172 ) ;
  assign n174 = ( x0 & x4 ) | ( x0 & ~n40 ) | ( x4 & ~n40 ) ;
  assign n175 = ( x0 & x4 ) | ( x0 & ~x10 ) | ( x4 & ~x10 ) ;
  assign n176 = ~n174 & n175 ;
  assign n177 = ( x13 & n173 ) | ( x13 & n176 ) | ( n173 & n176 ) ;
  assign n178 = ~n166 & n177 ;
  assign n179 = ( x13 & n166 ) | ( x13 & n178 ) | ( n166 & n178 ) ;
  assign n180 = ~x12 & n179 ;
  assign n181 = ( ~x12 & x13 ) | ( ~x12 & n179 ) | ( x13 & n179 ) ;
  assign n182 = ( n106 & n180 ) | ( n106 & ~n181 ) | ( n180 & ~n181 ) ;
  assign n183 = ( x1 & x11 ) | ( x1 & n77 ) | ( x11 & n77 ) ;
  assign n184 = ~x0 & x4 ;
  assign n185 = ( x8 & n116 ) | ( x8 & n184 ) | ( n116 & n184 ) ;
  assign n186 = ~x8 & n185 ;
  assign n187 = ( ~x9 & n16 ) | ( ~x9 & n52 ) | ( n16 & n52 ) ;
  assign n188 = x13 & ~n187 ;
  assign n189 = ( x13 & n52 ) | ( x13 & ~n188 ) | ( n52 & ~n188 ) ;
  assign n190 = ~x5 & n27 ;
  assign n191 = n31 & ~n190 ;
  assign n192 = ( x1 & ~n190 ) | ( x1 & n191 ) | ( ~n190 & n191 ) ;
  assign n193 = ( x1 & ~x5 ) | ( x1 & n192 ) | ( ~x5 & n192 ) ;
  assign n194 = ~n44 & n192 ;
  assign n195 = ( ~x1 & n193 ) | ( ~x1 & n194 ) | ( n193 & n194 ) ;
  assign n196 = ( x1 & ~x5 ) | ( x1 & n184 ) | ( ~x5 & n184 ) ;
  assign n197 = ( x1 & n184 ) | ( x1 & ~n196 ) | ( n184 & ~n196 ) ;
  assign n198 = n16 | n196 ;
  assign n199 = ( x5 & n196 ) | ( x5 & n198 ) | ( n196 & n198 ) ;
  assign n200 = ~n197 & n199 ;
  assign n201 = x9 & ~n200 ;
  assign n202 = x10 & n91 ;
  assign n203 = x9 | n202 ;
  assign n204 = ~n201 & n203 ;
  assign n205 = ( x8 & n195 ) | ( x8 & ~n204 ) | ( n195 & ~n204 ) ;
  assign n206 = x13 & n205 ;
  assign n207 = ( ~x13 & n195 ) | ( ~x13 & n206 ) | ( n195 & n206 ) ;
  assign n208 = ( n186 & ~n189 ) | ( n186 & n207 ) | ( ~n189 & n207 ) ;
  assign n209 = x1 & x5 ;
  assign n210 = n207 & ~n209 ;
  assign n211 = ( ~n186 & n208 ) | ( ~n186 & n210 ) | ( n208 & n210 ) ;
  assign n212 = x9 & ~n211 ;
  assign n213 = n22 & n212 ;
  assign n214 = x1 & n213 ;
  assign n215 = ( ~n77 & n183 ) | ( ~n77 & n214 ) | ( n183 & n214 ) ;
  assign n216 = ~n79 & n211 ;
  assign n217 = ~x5 & n81 ;
  assign n218 = ( x1 & x5 ) | ( x1 & ~x11 ) | ( x5 & ~x11 ) ;
  assign n219 = x1 & ~n218 ;
  assign n220 = ( x5 & n86 ) | ( x5 & n219 ) | ( n86 & n219 ) ;
  assign n221 = ( ~n218 & n219 ) | ( ~n218 & n220 ) | ( n219 & n220 ) ;
  assign n222 = n217 | n221 ;
  assign n223 = ( n211 & ~n216 ) | ( n211 & n222 ) | ( ~n216 & n222 ) ;
  assign n224 = ( x5 & n15 ) | ( x5 & ~n211 ) | ( n15 & ~n211 ) ;
  assign n225 = n61 | n211 ;
  assign n226 = ( n15 & ~n224 ) | ( n15 & n225 ) | ( ~n224 & n225 ) ;
  assign n227 = ( x9 & ~n223 ) | ( x9 & n226 ) | ( ~n223 & n226 ) ;
  assign n228 = ~x1 & x5 ;
  assign n229 = x5 & ~n228 ;
  assign n230 = n65 & n229 ;
  assign n231 = ( n49 & ~n228 ) | ( n49 & n229 ) | ( ~n228 & n229 ) ;
  assign n232 = ( ~x1 & n230 ) | ( ~x1 & n231 ) | ( n230 & n231 ) ;
  assign n233 = x5 | n232 ;
  assign n234 = ( n71 & n232 ) | ( n71 & n233 ) | ( n232 & n233 ) ;
  assign n235 = ( x9 & ~n226 ) | ( x9 & n234 ) | ( ~n226 & n234 ) ;
  assign n236 = n227 & ~n235 ;
  assign n237 = ( ~n103 & n215 ) | ( ~n103 & n236 ) | ( n215 & n236 ) ;
  assign n238 = ( n105 & ~n215 ) | ( n105 & n237 ) | ( ~n215 & n237 ) ;
  assign n239 = ( ~x8 & x9 ) | ( ~x8 & n211 ) | ( x9 & n211 ) ;
  assign n240 = ( x5 & x8 ) | ( x5 & x9 ) | ( x8 & x9 ) ;
  assign n241 = ~n239 & n240 ;
  assign n242 = x1 & n241 ;
  assign n243 = n211 | n242 ;
  assign n244 = ( ~n76 & n242 ) | ( ~n76 & n243 ) | ( n242 & n243 ) ;
  assign n245 = x1 & n114 ;
  assign n246 = ( n114 & ~n211 ) | ( n114 & n245 ) | ( ~n211 & n245 ) ;
  assign n247 = n116 | n246 ;
  assign n248 = ( n244 & n246 ) | ( n244 & n247 ) | ( n246 & n247 ) ;
  assign n249 = x0 & n125 ;
  assign n250 = n248 | n249 ;
  assign n251 = n248 & ~n249 ;
  assign n252 = ( ~n248 & n250 ) | ( ~n248 & n251 ) | ( n250 & n251 ) ;
  assign n253 = ( n112 & ~n169 ) | ( n112 & n252 ) | ( ~n169 & n252 ) ;
  assign n254 = n252 & ~n253 ;
  assign n255 = ~n66 & n211 ;
  assign n256 = x11 & ~n59 ;
  assign n257 = ( ~n66 & n211 ) | ( ~n66 & n256 ) | ( n211 & n256 ) ;
  assign n258 = ( n254 & ~n255 ) | ( n254 & n257 ) | ( ~n255 & n257 ) ;
  assign n259 = ( x1 & ~x13 ) | ( x1 & n258 ) | ( ~x13 & n258 ) ;
  assign n260 = ~x5 & n86 ;
  assign n261 = ~n57 & n130 ;
  assign n262 = n127 & ~n248 ;
  assign n263 = n209 | n262 ;
  assign n264 = ( n115 & n262 ) | ( n115 & n263 ) | ( n262 & n263 ) ;
  assign n265 = ( n211 & ~n261 ) | ( n211 & n264 ) | ( ~n261 & n264 ) ;
  assign n266 = ( n211 & n261 ) | ( n211 & ~n264 ) | ( n261 & ~n264 ) ;
  assign n267 = ( ~n211 & n265 ) | ( ~n211 & n266 ) | ( n265 & n266 ) ;
  assign n268 = n22 & ~n267 ;
  assign n269 = x8 | n252 ;
  assign n270 = x1 & ~n269 ;
  assign n271 = n268 | n270 ;
  assign n272 = ( n86 & ~n260 ) | ( n86 & n271 ) | ( ~n260 & n271 ) ;
  assign n273 = n112 & n272 ;
  assign n274 = x0 | x1 ;
  assign n275 = ( ~x11 & n150 ) | ( ~x11 & n274 ) | ( n150 & n274 ) ;
  assign n276 = ~x9 & n86 ;
  assign n277 = ~x5 & n68 ;
  assign n278 = ( x1 & n276 ) | ( x1 & n277 ) | ( n276 & n277 ) ;
  assign n279 = ~x1 & n278 ;
  assign n280 = x11 & n279 ;
  assign n281 = ( n150 & ~n275 ) | ( n150 & n280 ) | ( ~n275 & n280 ) ;
  assign n282 = ~n91 & n150 ;
  assign n283 = x11 | n17 ;
  assign n284 = x10 | n283 ;
  assign n285 = ~n68 & n276 ;
  assign n286 = ~x5 & n285 ;
  assign n287 = n284 & ~n286 ;
  assign n288 = ( ~n150 & n282 ) | ( ~n150 & n287 ) | ( n282 & n287 ) ;
  assign n289 = n66 & n211 ;
  assign n290 = x10 & ~n256 ;
  assign n291 = ( n76 & ~n256 ) | ( n76 & n290 ) | ( ~n256 & n290 ) ;
  assign n292 = ( n66 & n211 ) | ( n66 & ~n291 ) | ( n211 & ~n291 ) ;
  assign n293 = ( n288 & n289 ) | ( n288 & ~n292 ) | ( n289 & ~n292 ) ;
  assign n294 = x1 | n293 ;
  assign n295 = ~x10 & n71 ;
  assign n296 = x9 & n295 ;
  assign n297 = n125 & n130 ;
  assign n298 = ( n248 & ~n264 ) | ( n248 & n297 ) | ( ~n264 & n297 ) ;
  assign n299 = ( n248 & n264 ) | ( n248 & ~n297 ) | ( n264 & ~n297 ) ;
  assign n300 = ( ~n248 & n298 ) | ( ~n248 & n299 ) | ( n298 & n299 ) ;
  assign n301 = n296 & n300 ;
  assign n302 = ( ~n125 & n150 ) | ( ~n125 & n248 ) | ( n150 & n248 ) ;
  assign n303 = n125 & n302 ;
  assign n304 = ( ~n248 & n302 ) | ( ~n248 & n303 ) | ( n302 & n303 ) ;
  assign n305 = n145 | n304 ;
  assign n306 = ( ~n211 & n304 ) | ( ~n211 & n305 ) | ( n304 & n305 ) ;
  assign n307 = x11 & n306 ;
  assign n308 = ( x1 & ~n68 ) | ( x1 & n276 ) | ( ~n68 & n276 ) ;
  assign n309 = ( ~x1 & x5 ) | ( ~x1 & n68 ) | ( x5 & n68 ) ;
  assign n310 = n308 & n309 ;
  assign n311 = ~n57 & n211 ;
  assign n312 = n211 & ~n311 ;
  assign n313 = n136 & n312 ;
  assign n314 = ( x8 & x9 ) | ( x8 & ~x11 ) | ( x9 & ~x11 ) ;
  assign n315 = ~x8 & n314 ;
  assign n316 = ( ~x10 & x11 ) | ( ~x10 & n315 ) | ( x11 & n315 ) ;
  assign n317 = ( n314 & n315 ) | ( n314 & n316 ) | ( n315 & n316 ) ;
  assign n318 = ( ~n311 & n312 ) | ( ~n311 & n317 ) | ( n312 & n317 ) ;
  assign n319 = ( ~n57 & n313 ) | ( ~n57 & n318 ) | ( n313 & n318 ) ;
  assign n320 = n310 | n319 ;
  assign n321 = ( n306 & ~n307 ) | ( n306 & n320 ) | ( ~n307 & n320 ) ;
  assign n322 = n301 | n321 ;
  assign n323 = ( ~n293 & n294 ) | ( ~n293 & n322 ) | ( n294 & n322 ) ;
  assign n324 = n281 | n323 ;
  assign n325 = ( n272 & ~n273 ) | ( n272 & n324 ) | ( ~n273 & n324 ) ;
  assign n326 = x13 & n325 ;
  assign n327 = ( n258 & ~n259 ) | ( n258 & n326 ) | ( ~n259 & n326 ) ;
  assign n328 = n180 | n327 ;
  assign n329 = ( ~x13 & n180 ) | ( ~x13 & n327 ) | ( n180 & n327 ) ;
  assign n330 = ( n238 & ~n328 ) | ( n238 & n329 ) | ( ~n328 & n329 ) ;
  assign n331 = x9 & n77 ;
  assign n332 = ( x6 & n77 ) | ( x6 & n331 ) | ( n77 & n331 ) ;
  assign n333 = x11 & ~n332 ;
  assign n334 = x2 & n333 ;
  assign n335 = x9 & ~n71 ;
  assign n336 = x11 & n86 ;
  assign n337 = ~x2 & n336 ;
  assign n338 = x9 | n337 ;
  assign n339 = ~n335 & n338 ;
  assign n340 = ~x6 & n339 ;
  assign n341 = ( ~x1 & x5 ) | ( ~x1 & n184 ) | ( x5 & n184 ) ;
  assign n342 = x6 & ~n341 ;
  assign n343 = x6 & ~n342 ;
  assign n344 = n16 & n343 ;
  assign n345 = ( x9 & ~n342 ) | ( x9 & n343 ) | ( ~n342 & n343 ) ;
  assign n346 = ( ~n341 & n344 ) | ( ~n341 & n345 ) | ( n344 & n345 ) ;
  assign n347 = ( ~x2 & x8 ) | ( ~x2 & n346 ) | ( x8 & n346 ) ;
  assign n348 = x1 & x11 ;
  assign n349 = ( x9 & x10 ) | ( x9 & n348 ) | ( x10 & n348 ) ;
  assign n350 = ~x9 & n349 ;
  assign n351 = x6 | n341 ;
  assign n352 = n16 & ~n341 ;
  assign n353 = x6 & n352 ;
  assign n354 = ( ~x6 & n351 ) | ( ~x6 & n353 ) | ( n351 & n353 ) ;
  assign n355 = ( ~x2 & n350 ) | ( ~x2 & n354 ) | ( n350 & n354 ) ;
  assign n356 = x9 & ~n355 ;
  assign n357 = ( x9 & n350 ) | ( x9 & ~n356 ) | ( n350 & ~n356 ) ;
  assign n358 = ~x8 & n357 ;
  assign n359 = ( n346 & ~n347 ) | ( n346 & n358 ) | ( ~n347 & n358 ) ;
  assign n360 = ~x13 & n359 ;
  assign n361 = x2 & ~n44 ;
  assign n362 = ( x2 & x6 ) | ( x2 & n44 ) | ( x6 & n44 ) ;
  assign n363 = x2 | n31 ;
  assign n364 = ( n361 & ~n362 ) | ( n361 & n363 ) | ( ~n362 & n363 ) ;
  assign n365 = x6 | n27 ;
  assign n366 = x2 & n189 ;
  assign n367 = x6 & ~n366 ;
  assign n368 = n365 & ~n367 ;
  assign n369 = n364 & ~n368 ;
  assign n370 = ( ~n359 & n360 ) | ( ~n359 & n369 ) | ( n360 & n369 ) ;
  assign n371 = ( x6 & n15 ) | ( x6 & ~n370 ) | ( n15 & ~n370 ) ;
  assign n372 = ( x2 & n22 ) | ( x2 & ~n61 ) | ( n22 & ~n61 ) ;
  assign n373 = x9 & ~n372 ;
  assign n374 = ( ~x9 & n61 ) | ( ~x9 & n373 ) | ( n61 & n373 ) ;
  assign n375 = n370 | n374 ;
  assign n376 = ( n15 & ~n371 ) | ( n15 & n375 ) | ( ~n371 & n375 ) ;
  assign n377 = ~x2 & x6 ;
  assign n378 = x6 & ~n377 ;
  assign n379 = n65 & n378 ;
  assign n380 = ( n49 & ~n377 ) | ( n49 & n378 ) | ( ~n377 & n378 ) ;
  assign n381 = ( ~x2 & n379 ) | ( ~x2 & n380 ) | ( n379 & n380 ) ;
  assign n382 = x9 & n381 ;
  assign n383 = n79 & n370 ;
  assign n384 = n81 | n383 ;
  assign n385 = ( ~x6 & n383 ) | ( ~x6 & n384 ) | ( n383 & n384 ) ;
  assign n386 = x9 | n385 ;
  assign n387 = ( ~x9 & n382 ) | ( ~x9 & n386 ) | ( n382 & n386 ) ;
  assign n388 = n376 & ~n387 ;
  assign n389 = ( ~n339 & n340 ) | ( ~n339 & n388 ) | ( n340 & n388 ) ;
  assign n390 = ( ~n103 & n334 ) | ( ~n103 & n389 ) | ( n334 & n389 ) ;
  assign n391 = ( n105 & ~n334 ) | ( n105 & n390 ) | ( ~n334 & n390 ) ;
  assign n392 = n180 & n327 ;
  assign n393 = ( x1 & n66 ) | ( x1 & ~n211 ) | ( n66 & ~n211 ) ;
  assign n394 = x2 | n393 ;
  assign n395 = ~n393 & n394 ;
  assign n396 = ~n291 & n395 ;
  assign n397 = ( n256 & n394 ) | ( n256 & n395 ) | ( n394 & n395 ) ;
  assign n398 = ( ~x2 & n396 ) | ( ~x2 & n397 ) | ( n396 & n397 ) ;
  assign n399 = ( x13 & n370 ) | ( x13 & ~n398 ) | ( n370 & ~n398 ) ;
  assign n400 = ( x1 & x5 ) | ( x1 & n68 ) | ( x5 & n68 ) ;
  assign n401 = ~x2 & x11 ;
  assign n402 = ( x2 & n400 ) | ( x2 & ~n401 ) | ( n400 & ~n401 ) ;
  assign n403 = ( x6 & n400 ) | ( x6 & ~n402 ) | ( n400 & ~n402 ) ;
  assign n404 = ( x6 & n400 ) | ( x6 & ~n403 ) | ( n400 & ~n403 ) ;
  assign n405 = ( x2 & n403 ) | ( x2 & ~n404 ) | ( n403 & ~n404 ) ;
  assign n406 = ( x1 & n248 ) | ( x1 & n249 ) | ( n248 & n249 ) ;
  assign n407 = ( ~x8 & x9 ) | ( ~x8 & n370 ) | ( x9 & n370 ) ;
  assign n408 = ( x6 & x8 ) | ( x6 & x9 ) | ( x8 & x9 ) ;
  assign n409 = ~n407 & n408 ;
  assign n410 = x2 & n409 ;
  assign n411 = n370 | n410 ;
  assign n412 = ( ~n76 & n410 ) | ( ~n76 & n411 ) | ( n410 & n411 ) ;
  assign n413 = x2 & n114 ;
  assign n414 = ( n114 & ~n370 ) | ( n114 & n413 ) | ( ~n370 & n413 ) ;
  assign n415 = n116 | n414 ;
  assign n416 = ( n412 & n414 ) | ( n412 & n415 ) | ( n414 & n415 ) ;
  assign n417 = ~n406 & n416 ;
  assign n418 = n406 & n416 ;
  assign n419 = ( n406 & n417 ) | ( n406 & ~n418 ) | ( n417 & ~n418 ) ;
  assign n420 = ( n112 & ~n169 ) | ( n112 & n419 ) | ( ~n169 & n419 ) ;
  assign n421 = n419 & ~n420 ;
  assign n422 = ( n370 & n393 ) | ( n370 & ~n421 ) | ( n393 & ~n421 ) ;
  assign n423 = n256 & n422 ;
  assign n424 = ( n256 & n421 ) | ( n256 & ~n423 ) | ( n421 & ~n423 ) ;
  assign n425 = x2 & n424 ;
  assign n426 = ( n248 & n264 ) | ( n248 & n297 ) | ( n264 & n297 ) ;
  assign n427 = x6 & n115 ;
  assign n428 = x2 & n427 ;
  assign n429 = n127 | n428 ;
  assign n430 = ( ~n416 & n428 ) | ( ~n416 & n429 ) | ( n428 & n429 ) ;
  assign n431 = ( n416 & n426 ) | ( n416 & ~n430 ) | ( n426 & ~n430 ) ;
  assign n432 = ( n416 & ~n426 ) | ( n416 & n430 ) | ( ~n426 & n430 ) ;
  assign n433 = ( ~n416 & n431 ) | ( ~n416 & n432 ) | ( n431 & n432 ) ;
  assign n434 = n296 & n433 ;
  assign n435 = ( ~n211 & n261 ) | ( ~n211 & n264 ) | ( n261 & n264 ) ;
  assign n436 = ( n370 & n430 ) | ( n370 & ~n435 ) | ( n430 & ~n435 ) ;
  assign n437 = ( n370 & ~n430 ) | ( n370 & n435 ) | ( ~n430 & n435 ) ;
  assign n438 = ( ~n370 & n436 ) | ( ~n370 & n437 ) | ( n436 & n437 ) ;
  assign n439 = n22 & ~n438 ;
  assign n440 = x8 | n419 ;
  assign n441 = x2 & ~n440 ;
  assign n442 = x6 | n441 ;
  assign n443 = ( n86 & n441 ) | ( n86 & n442 ) | ( n441 & n442 ) ;
  assign n444 = ( n284 & n291 ) | ( n284 & n370 ) | ( n291 & n370 ) ;
  assign n445 = n393 & n444 ;
  assign n446 = ( n284 & ~n393 ) | ( n284 & n445 ) | ( ~n393 & n445 ) ;
  assign n447 = x2 | n446 ;
  assign n448 = n57 & n211 ;
  assign n449 = ( n317 & ~n370 ) | ( n317 & n448 ) | ( ~n370 & n448 ) ;
  assign n450 = ~x11 & n145 ;
  assign n451 = ~n370 & n450 ;
  assign n452 = ( ~n448 & n449 ) | ( ~n448 & n451 ) | ( n449 & n451 ) ;
  assign n453 = x2 & n274 ;
  assign n454 = ( x2 & x11 ) | ( x2 & n274 ) | ( x11 & n274 ) ;
  assign n455 = n125 | n248 ;
  assign n456 = n416 & ~n455 ;
  assign n457 = n416 & n455 ;
  assign n458 = ( n455 & n456 ) | ( n455 & ~n457 ) | ( n456 & ~n457 ) ;
  assign n459 = ~x11 & n458 ;
  assign n460 = ( ~n453 & n454 ) | ( ~n453 & n459 ) | ( n454 & n459 ) ;
  assign n461 = n150 & ~n460 ;
  assign n462 = n370 & n448 ;
  assign n463 = n461 | n462 ;
  assign n464 = ( n136 & n461 ) | ( n136 & n463 ) | ( n461 & n463 ) ;
  assign n465 = n452 | n464 ;
  assign n466 = ( ~n446 & n447 ) | ( ~n446 & n465 ) | ( n447 & n465 ) ;
  assign n467 = ( ~n439 & n443 ) | ( ~n439 & n466 ) | ( n443 & n466 ) ;
  assign n468 = n112 & ~n466 ;
  assign n469 = ( n439 & n467 ) | ( n439 & ~n468 ) | ( n467 & ~n468 ) ;
  assign n470 = n434 | n469 ;
  assign n471 = ( n424 & ~n425 ) | ( n424 & n470 ) | ( ~n425 & n470 ) ;
  assign n472 = n276 | n471 ;
  assign n473 = ( n405 & n471 ) | ( n405 & n472 ) | ( n471 & n472 ) ;
  assign n474 = x13 & n473 ;
  assign n475 = ( n398 & n399 ) | ( n398 & n474 ) | ( n399 & n474 ) ;
  assign n476 = n392 | n475 ;
  assign n477 = ( ~x13 & n392 ) | ( ~x13 & n475 ) | ( n392 & n475 ) ;
  assign n478 = ( n391 & ~n476 ) | ( n391 & n477 ) | ( ~n476 & n477 ) ;
  assign n479 = ( x7 & n77 ) | ( x7 & n331 ) | ( n77 & n331 ) ;
  assign n480 = x11 & ~n479 ;
  assign n481 = x3 & n480 ;
  assign n482 = ~x3 & n336 ;
  assign n483 = x9 | n482 ;
  assign n484 = ~n335 & n483 ;
  assign n485 = ~x7 & n484 ;
  assign n486 = ( ~x2 & x6 ) | ( ~x2 & n341 ) | ( x6 & n341 ) ;
  assign n487 = x9 & ~n486 ;
  assign n488 = x3 & n487 ;
  assign n489 = ( ~x8 & n27 ) | ( ~x8 & n488 ) | ( n27 & n488 ) ;
  assign n490 = x13 & ~n489 ;
  assign n491 = ( x13 & n27 ) | ( x13 & ~n490 ) | ( n27 & ~n490 ) ;
  assign n492 = x7 & n491 ;
  assign n493 = ( x13 & n16 ) | ( x13 & ~n486 ) | ( n16 & ~n486 ) ;
  assign n494 = ~x9 & n16 ;
  assign n495 = ( n486 & n493 ) | ( n486 & n494 ) | ( n493 & n494 ) ;
  assign n496 = x3 & x7 ;
  assign n497 = ( x8 & n495 ) | ( x8 & ~n496 ) | ( n495 & ~n496 ) ;
  assign n498 = x2 & x11 ;
  assign n499 = ( x9 & x10 ) | ( x9 & n498 ) | ( x10 & n498 ) ;
  assign n500 = ~x9 & n499 ;
  assign n501 = x3 | x7 ;
  assign n502 = ( n486 & n500 ) | ( n486 & ~n501 ) | ( n500 & ~n501 ) ;
  assign n503 = x9 & ~n502 ;
  assign n504 = ( x9 & n500 ) | ( x9 & ~n503 ) | ( n500 & ~n503 ) ;
  assign n505 = ( x9 & x10 ) | ( x9 & n64 ) | ( x10 & n64 ) ;
  assign n506 = ~x13 & n505 ;
  assign n507 = n16 & n487 ;
  assign n508 = x7 & n507 ;
  assign n509 = x13 & ~n508 ;
  assign n510 = n506 | n509 ;
  assign n511 = x3 | n510 ;
  assign n512 = ~x13 & n511 ;
  assign n513 = ( ~n504 & n511 ) | ( ~n504 & n512 ) | ( n511 & n512 ) ;
  assign n514 = x8 | n513 ;
  assign n515 = ( ~n495 & n497 ) | ( ~n495 & n514 ) | ( n497 & n514 ) ;
  assign n516 = ( ~x3 & x7 ) | ( ~x3 & n44 ) | ( x7 & n44 ) ;
  assign n517 = ( x9 & x13 ) | ( x9 & n16 ) | ( x13 & n16 ) ;
  assign n518 = x13 & n48 ;
  assign n519 = ( ~x9 & n517 ) | ( ~x9 & n518 ) | ( n517 & n518 ) ;
  assign n520 = ( x3 & n44 ) | ( x3 & n519 ) | ( n44 & n519 ) ;
  assign n521 = ~n516 & n520 ;
  assign n522 = ( x7 & n44 ) | ( x7 & n521 ) | ( n44 & n521 ) ;
  assign n523 = n515 & ~n522 ;
  assign n524 = ( ~n491 & n492 ) | ( ~n491 & n523 ) | ( n492 & n523 ) ;
  assign n525 = ( x7 & n15 ) | ( x7 & ~n524 ) | ( n15 & ~n524 ) ;
  assign n526 = n61 | n524 ;
  assign n527 = ( n15 & ~n525 ) | ( n15 & n526 ) | ( ~n525 & n526 ) ;
  assign n528 = x3 & ~n524 ;
  assign n529 = ~x3 & x7 ;
  assign n530 = x7 & ~n529 ;
  assign n531 = n65 & n530 ;
  assign n532 = ( n49 & ~n529 ) | ( n49 & n530 ) | ( ~n529 & n530 ) ;
  assign n533 = ( ~x3 & n531 ) | ( ~x3 & n532 ) | ( n531 & n532 ) ;
  assign n534 = n22 | n533 ;
  assign n535 = ( n528 & n533 ) | ( n528 & n534 ) | ( n533 & n534 ) ;
  assign n536 = x9 & n535 ;
  assign n537 = n79 & n524 ;
  assign n538 = n81 | n537 ;
  assign n539 = ( ~x7 & n537 ) | ( ~x7 & n538 ) | ( n537 & n538 ) ;
  assign n540 = x9 | n539 ;
  assign n541 = ( ~x9 & n536 ) | ( ~x9 & n540 ) | ( n536 & n540 ) ;
  assign n542 = n527 & ~n541 ;
  assign n543 = ( ~n484 & n485 ) | ( ~n484 & n542 ) | ( n485 & n542 ) ;
  assign n544 = ( ~n103 & n481 ) | ( ~n103 & n543 ) | ( n481 & n543 ) ;
  assign n545 = ( n105 & ~n481 ) | ( n105 & n544 ) | ( ~n481 & n544 ) ;
  assign n546 = n392 & n475 ;
  assign n547 = n317 | n450 ;
  assign n548 = ( n450 & ~n462 ) | ( n450 & n547 ) | ( ~n462 & n547 ) ;
  assign n549 = ( ~x13 & n524 ) | ( ~x13 & n548 ) | ( n524 & n548 ) ;
  assign n550 = ( n76 & ~n116 ) | ( n76 & n524 ) | ( ~n116 & n524 ) ;
  assign n551 = ( x8 & ~x9 ) | ( x8 & n528 ) | ( ~x9 & n528 ) ;
  assign n552 = ( x8 & x9 ) | ( x8 & n496 ) | ( x9 & n496 ) ;
  assign n553 = n551 & n552 ;
  assign n554 = n116 & n553 ;
  assign n555 = ( n524 & ~n550 ) | ( n524 & n554 ) | ( ~n550 & n554 ) ;
  assign n556 = ( x3 & n524 ) | ( x3 & ~n555 ) | ( n524 & ~n555 ) ;
  assign n557 = n114 | n555 ;
  assign n558 = ( x3 & ~n556 ) | ( x3 & n557 ) | ( ~n556 & n557 ) ;
  assign n559 = n127 & ~n558 ;
  assign n560 = n496 | n559 ;
  assign n561 = ( n115 & n559 ) | ( n115 & n560 ) | ( n559 & n560 ) ;
  assign n562 = ( ~n370 & n430 ) | ( ~n370 & n435 ) | ( n430 & n435 ) ;
  assign n563 = ( n524 & ~n561 ) | ( n524 & n562 ) | ( ~n561 & n562 ) ;
  assign n564 = ( n524 & n561 ) | ( n524 & ~n562 ) | ( n561 & ~n562 ) ;
  assign n565 = ( ~n524 & n563 ) | ( ~n524 & n564 ) | ( n563 & n564 ) ;
  assign n566 = x8 & ~n565 ;
  assign n567 = ( x2 & n406 ) | ( x2 & n416 ) | ( n406 & n416 ) ;
  assign n568 = ( x3 & n558 ) | ( x3 & n567 ) | ( n558 & n567 ) ;
  assign n569 = ( ~x8 & n558 ) | ( ~x8 & n567 ) | ( n558 & n567 ) ;
  assign n570 = ~n568 & n569 ;
  assign n571 = ~n566 & n570 ;
  assign n572 = ( n494 & n566 ) | ( n494 & n571 ) | ( n566 & n571 ) ;
  assign n573 = ( x2 & ~n370 ) | ( x2 & n393 ) | ( ~n370 & n393 ) ;
  assign n574 = n524 | n573 ;
  assign n575 = ~n524 & n573 ;
  assign n576 = ( ~n573 & n574 ) | ( ~n573 & n575 ) | ( n574 & n575 ) ;
  assign n577 = ( ~x3 & n256 ) | ( ~x3 & n576 ) | ( n256 & n576 ) ;
  assign n578 = ( x2 & x6 ) | ( x2 & n400 ) | ( x6 & n400 ) ;
  assign n579 = x7 & ~n578 ;
  assign n580 = n276 & n579 ;
  assign n581 = ~x3 & n580 ;
  assign n582 = ( ~n576 & n577 ) | ( ~n576 & n581 ) | ( n577 & n581 ) ;
  assign n583 = ( n416 & n426 ) | ( n416 & n430 ) | ( n426 & n430 ) ;
  assign n584 = ( n558 & n561 ) | ( n558 & ~n583 ) | ( n561 & ~n583 ) ;
  assign n585 = ( n558 & ~n561 ) | ( n558 & n583 ) | ( ~n561 & n583 ) ;
  assign n586 = ( ~n558 & n584 ) | ( ~n558 & n585 ) | ( n584 & n585 ) ;
  assign n587 = n145 & n586 ;
  assign n588 = ~n501 & n578 ;
  assign n589 = n276 & n588 ;
  assign n590 = x2 | n274 ;
  assign n591 = ~x3 & n150 ;
  assign n592 = ~n590 & n591 ;
  assign n593 = ( x11 & n589 ) | ( x11 & n592 ) | ( n589 & n592 ) ;
  assign n594 = ~n587 & n593 ;
  assign n595 = ( x11 & n587 ) | ( x11 & n594 ) | ( n587 & n594 ) ;
  assign n596 = ( n76 & ~n558 ) | ( n76 & n567 ) | ( ~n558 & n567 ) ;
  assign n597 = n567 & ~n596 ;
  assign n598 = ( n558 & n596 ) | ( n558 & ~n597 ) | ( n596 & ~n597 ) ;
  assign n599 = x3 & ~n598 ;
  assign n600 = x7 | n599 ;
  assign n601 = ( n276 & n599 ) | ( n276 & n600 ) | ( n599 & n600 ) ;
  assign n602 = n416 | n455 ;
  assign n603 = ~n558 & n602 ;
  assign n604 = ( n150 & ~n558 ) | ( n150 & n602 ) | ( ~n558 & n602 ) ;
  assign n605 = ( n601 & ~n603 ) | ( n601 & n604 ) | ( ~n603 & n604 ) ;
  assign n606 = x11 & n605 ;
  assign n607 = ( x3 & x7 ) | ( x3 & ~n578 ) | ( x7 & ~n578 ) ;
  assign n608 = ( ~x7 & n276 ) | ( ~x7 & n578 ) | ( n276 & n578 ) ;
  assign n609 = n607 & n608 ;
  assign n610 = n462 & n524 ;
  assign n611 = ~n136 & n610 ;
  assign n612 = x11 & n150 ;
  assign n613 = ( x3 & ~n590 ) | ( x3 & n612 ) | ( ~n590 & n612 ) ;
  assign n614 = n590 & n613 ;
  assign n615 = ( x3 & n291 ) | ( x3 & n576 ) | ( n291 & n576 ) ;
  assign n616 = x3 & ~n284 ;
  assign n617 = ( ~n291 & n615 ) | ( ~n291 & n616 ) | ( n615 & n616 ) ;
  assign n618 = n614 | n617 ;
  assign n619 = ( n610 & ~n611 ) | ( n610 & n618 ) | ( ~n611 & n618 ) ;
  assign n620 = n609 | n619 ;
  assign n621 = ( n605 & ~n606 ) | ( n605 & n620 ) | ( ~n606 & n620 ) ;
  assign n622 = n595 | n621 ;
  assign n623 = ( ~n572 & n582 ) | ( ~n572 & n622 ) | ( n582 & n622 ) ;
  assign n624 = n572 | n623 ;
  assign n625 = x13 & n624 ;
  assign n626 = ( n548 & ~n549 ) | ( n548 & n625 ) | ( ~n549 & n625 ) ;
  assign n627 = n546 | n626 ;
  assign n628 = ( ~x13 & n546 ) | ( ~x13 & n626 ) | ( n546 & n626 ) ;
  assign n629 = ( n545 & ~n627 ) | ( n545 & n628 ) | ( ~n627 & n628 ) ;
  assign n630 = x3 & ~x7 ;
  assign n631 = ( ~x3 & n501 ) | ( ~x3 & n630 ) | ( n501 & n630 ) ;
  assign n632 = x8 & ~n133 ;
  assign n633 = ( x10 & ~x11 ) | ( x10 & n632 ) | ( ~x11 & n632 ) ;
  assign n634 = ( ~n133 & n632 ) | ( ~n133 & n633 ) | ( n632 & n633 ) ;
  assign n635 = ( x13 & n610 ) | ( x13 & ~n634 ) | ( n610 & ~n634 ) ;
  assign n636 = ( n558 & n561 ) | ( n558 & n583 ) | ( n561 & n583 ) ;
  assign n637 = n145 & n636 ;
  assign n638 = ( x3 & ~n524 ) | ( x3 & n573 ) | ( ~n524 & n573 ) ;
  assign n639 = n59 & n638 ;
  assign n640 = ( x3 & x7 ) | ( x3 & n578 ) | ( x7 & n578 ) ;
  assign n641 = n276 & n640 ;
  assign n642 = n592 | n641 ;
  assign n643 = ( n638 & ~n639 ) | ( n638 & n642 ) | ( ~n639 & n642 ) ;
  assign n644 = ( n17 & n558 ) | ( n17 & ~n602 ) | ( n558 & ~n602 ) ;
  assign n645 = ( n97 & ~n558 ) | ( n97 & n644 ) | ( ~n558 & n644 ) ;
  assign n646 = ( ~n524 & n561 ) | ( ~n524 & n562 ) | ( n561 & n562 ) ;
  assign n647 = x8 & n646 ;
  assign n648 = x8 | n568 ;
  assign n649 = ( ~x8 & n647 ) | ( ~x8 & n648 ) | ( n647 & n648 ) ;
  assign n650 = ( ~x9 & n645 ) | ( ~x9 & n649 ) | ( n645 & n649 ) ;
  assign n651 = x10 & ~n650 ;
  assign n652 = ( x10 & n645 ) | ( x10 & ~n651 ) | ( n645 & ~n651 ) ;
  assign n653 = n546 & n626 ;
  assign n654 = x11 & ~n653 ;
  assign n655 = ( n652 & n653 ) | ( n652 & ~n654 ) | ( n653 & ~n654 ) ;
  assign n656 = ( ~n637 & n643 ) | ( ~n637 & n655 ) | ( n643 & n655 ) ;
  assign n657 = x11 | n655 ;
  assign n658 = ( n637 & n656 ) | ( n637 & n657 ) | ( n656 & n657 ) ;
  assign n659 = x13 & n658 ;
  assign n660 = ( n634 & n635 ) | ( n634 & n659 ) | ( n635 & n659 ) ;
  assign n661 = ( ~x2 & x6 ) | ( ~x2 & n274 ) | ( x6 & n274 ) ;
  assign n662 = ( x2 & x5 ) | ( x2 & ~x6 ) | ( x5 & ~x6 ) ;
  assign n663 = n661 | n662 ;
  assign n664 = ( ~x4 & n631 ) | ( ~x4 & n663 ) | ( n631 & n663 ) ;
  assign n665 = ( x0 & ~x4 ) | ( x0 & n228 ) | ( ~x4 & n228 ) ;
  assign n666 = ( x1 & x4 ) | ( x1 & n228 ) | ( x4 & n228 ) ;
  assign n667 = ( x0 & x5 ) | ( x0 & ~n666 ) | ( x5 & ~n666 ) ;
  assign n668 = ~n665 & n667 ;
  assign n669 = ( x2 & ~x6 ) | ( x2 & n668 ) | ( ~x6 & n668 ) ;
  assign n670 = ~x2 & n669 ;
  assign n671 = ( x6 & n669 ) | ( x6 & n670 ) | ( n669 & n670 ) ;
  assign n672 = ~n631 & n671 ;
  assign n673 = ( x4 & n664 ) | ( x4 & ~n672 ) | ( n664 & ~n672 ) ;
  assign y0 = ~n182 ;
  assign y1 = ~n330 ;
  assign y2 = ~n478 ;
  assign y3 = ~n629 ;
  assign y4 = ~n631 ;
  assign y5 = n496 ;
  assign y6 = n660 ;
  assign y7 = ~n673 ;
endmodule
