module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 ;
  assign n9 = x5 & ~x7 ;
  assign n10 = x1 & n9 ;
  assign n11 = ( x2 & x4 ) | ( x2 & n10 ) | ( x4 & n10 ) ;
  assign n12 = ~x4 & n11 ;
  assign n13 = ( x1 & x2 ) | ( x1 & x5 ) | ( x2 & x5 ) ;
  assign n14 = ( ~x2 & x4 ) | ( ~x2 & n13 ) | ( x4 & n13 ) ;
  assign n15 = ( x1 & x5 ) | ( x1 & n14 ) | ( x5 & n14 ) ;
  assign n16 = ~n13 & n15 ;
  assign n17 = ( ~n14 & n15 ) | ( ~n14 & n16 ) | ( n15 & n16 ) ;
  assign n22 = ( x6 & ~x7 ) | ( x6 & n17 ) | ( ~x7 & n17 ) ;
  assign n19 = ~x1 & x2 ;
  assign n18 = ~x5 & x6 ;
  assign n20 = x4 & n18 ;
  assign n21 = n19 & n20 ;
  assign n23 = x7 & n21 ;
  assign n24 = ( n17 & ~n22 ) | ( n17 & n23 ) | ( ~n22 & n23 ) ;
  assign n25 = ~x0 & x2 ;
  assign n26 = x1 & n25 ;
  assign n27 = x6 & ~x7 ;
  assign n28 = x5 & n27 ;
  assign n29 = ( x4 & ~n26 ) | ( x4 & n28 ) | ( ~n26 & n28 ) ;
  assign n30 = n26 & n29 ;
  assign n31 = ( ~n12 & n24 ) | ( ~n12 & n30 ) | ( n24 & n30 ) ;
  assign n32 = x0 | n30 ;
  assign n33 = ( n12 & n31 ) | ( n12 & n32 ) | ( n31 & n32 ) ;
  assign n52 = ~x3 & n33 ;
  assign n34 = x0 & x2 ;
  assign n35 = x1 & n34 ;
  assign n36 = x5 & x7 ;
  assign n37 = ( x4 & x6 ) | ( x4 & n36 ) | ( x6 & n36 ) ;
  assign n38 = ~x4 & n37 ;
  assign n39 = n35 & n38 ;
  assign n40 = ( x1 & ~x2 ) | ( x1 & x5 ) | ( ~x2 & x5 ) ;
  assign n41 = ( x1 & x5 ) | ( x1 & ~x6 ) | ( x5 & ~x6 ) ;
  assign n42 = ~n40 & n41 ;
  assign n49 = ( x0 & x4 ) | ( x0 & ~n42 ) | ( x4 & ~n42 ) ;
  assign n44 = ( x1 & x5 ) | ( x1 & x6 ) | ( x5 & x6 ) ;
  assign n45 = x0 & ~n44 ;
  assign n43 = x6 & n36 ;
  assign n46 = x1 & n43 ;
  assign n47 = x0 | n46 ;
  assign n48 = ~n45 & n47 ;
  assign n50 = x4 & n48 ;
  assign n51 = ( n42 & n49 ) | ( n42 & n50 ) | ( n49 & n50 ) ;
  assign n53 = n39 | n51 ;
  assign n54 = ( n33 & ~n52 ) | ( n33 & n53 ) | ( ~n52 & n53 ) ;
  assign n57 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n58 = ( x2 & ~x5 ) | ( x2 & n57 ) | ( ~x5 & n57 ) ;
  assign n59 = ( x2 & x4 ) | ( x2 & ~n57 ) | ( x4 & ~n57 ) ;
  assign n60 = n58 & ~n59 ;
  assign n61 = x0 & ~n60 ;
  assign n55 = ~x4 & x5 ;
  assign n56 = x3 & n55 ;
  assign n62 = x2 & n56 ;
  assign n63 = x0 | n62 ;
  assign n64 = ~n61 & n63 ;
  assign n70 = ( ~x1 & x6 ) | ( ~x1 & n64 ) | ( x6 & n64 ) ;
  assign n65 = ~x0 & x3 ;
  assign n66 = ~x2 & n65 ;
  assign n67 = x5 & x6 ;
  assign n68 = ~x4 & n67 ;
  assign n69 = n66 & n68 ;
  assign n71 = x1 & n69 ;
  assign n72 = ( n64 & ~n70 ) | ( n64 & n71 ) | ( ~n70 & n71 ) ;
  assign n80 = ~x4 & n35 ;
  assign n81 = ( x3 & n67 ) | ( x3 & n80 ) | ( n67 & n80 ) ;
  assign n82 = ~x3 & n81 ;
  assign n84 = ( ~x0 & x1 ) | ( ~x0 & x5 ) | ( x1 & x5 ) ;
  assign n85 = ( x0 & ~x6 ) | ( x0 & n84 ) | ( ~x6 & n84 ) ;
  assign n86 = ( x1 & x5 ) | ( x1 & n85 ) | ( x5 & n85 ) ;
  assign n87 = ~n84 & n86 ;
  assign n88 = ( ~n85 & n86 ) | ( ~n85 & n87 ) | ( n86 & n87 ) ;
  assign n89 = x2 | n88 ;
  assign n83 = x0 & ~x1 ;
  assign n90 = n18 & n83 ;
  assign n91 = x2 & ~n90 ;
  assign n92 = n89 & ~n91 ;
  assign n96 = ( x3 & x4 ) | ( x3 & ~n92 ) | ( x4 & ~n92 ) ;
  assign n93 = ~x3 & n67 ;
  assign n94 = ~x0 & x1 ;
  assign n95 = n93 & n94 ;
  assign n97 = x4 & n95 ;
  assign n98 = ( n92 & n96 ) | ( n92 & n97 ) | ( n96 & n97 ) ;
  assign n99 = ( x3 & x6 ) | ( x3 & n41 ) | ( x6 & n41 ) ;
  assign n100 = ( x1 & x5 ) | ( x1 & n99 ) | ( x5 & n99 ) ;
  assign n101 = ~n41 & n100 ;
  assign n102 = ( ~n99 & n100 ) | ( ~n99 & n101 ) | ( n100 & n101 ) ;
  assign n103 = x2 & ~n102 ;
  assign n104 = x1 & n93 ;
  assign n105 = x2 | n104 ;
  assign n106 = ~n103 & n105 ;
  assign n107 = ~x0 & x7 ;
  assign n108 = ( x4 & n106 ) | ( x4 & ~n107 ) | ( n106 & ~n107 ) ;
  assign n109 = n106 & ~n108 ;
  assign n110 = ( ~n82 & n98 ) | ( ~n82 & n109 ) | ( n98 & n109 ) ;
  assign n111 = x7 & ~n109 ;
  assign n112 = ( n82 & n110 ) | ( n82 & ~n111 ) | ( n110 & ~n111 ) ;
  assign n73 = ( x2 & ~x4 ) | ( x2 & x5 ) | ( ~x4 & x5 ) ;
  assign n74 = ( x5 & x6 ) | ( x5 & ~n73 ) | ( x6 & ~n73 ) ;
  assign n75 = ( ~x2 & x6 ) | ( ~x2 & n73 ) | ( x6 & n73 ) ;
  assign n76 = n74 & ~n75 ;
  assign n77 = x0 & ~x3 ;
  assign n78 = ( x1 & n76 ) | ( x1 & n77 ) | ( n76 & n77 ) ;
  assign n79 = ~x1 & n78 ;
  assign n113 = ( ~x2 & x4 ) | ( ~x2 & x5 ) | ( x4 & x5 ) ;
  assign n114 = ( x1 & ~x5 ) | ( x1 & n113 ) | ( ~x5 & n113 ) ;
  assign n115 = ( x1 & x4 ) | ( x1 & ~n113 ) | ( x4 & ~n113 ) ;
  assign n116 = n114 & ~n115 ;
  assign n132 = ~x0 & n116 ;
  assign n117 = x0 & ~x4 ;
  assign n118 = x1 & x5 ;
  assign n119 = ( ~x0 & x4 ) | ( ~x0 & n118 ) | ( x4 & n118 ) ;
  assign n120 = ( n117 & ~n118 ) | ( n117 & n119 ) | ( ~n118 & n119 ) ;
  assign n123 = ( x4 & ~x5 ) | ( x4 & x6 ) | ( ~x5 & x6 ) ;
  assign n124 = x4 & ~n123 ;
  assign n125 = ( x2 & x6 ) | ( x2 & n124 ) | ( x6 & n124 ) ;
  assign n126 = ( ~n123 & n124 ) | ( ~n123 & n125 ) | ( n124 & n125 ) ;
  assign n127 = x1 & n126 ;
  assign n128 = x0 | n127 ;
  assign n121 = x4 & ~x5 ;
  assign n122 = ~x6 & n121 ;
  assign n129 = n19 & n122 ;
  assign n130 = x0 & ~n129 ;
  assign n131 = n128 & ~n130 ;
  assign n133 = n120 | n131 ;
  assign n134 = ( n116 & ~n132 ) | ( n116 & n133 ) | ( ~n132 & n133 ) ;
  assign n135 = n79 | n134 ;
  assign n136 = ( ~n72 & n112 ) | ( ~n72 & n135 ) | ( n112 & n135 ) ;
  assign n137 = n72 | n136 ;
  assign n156 = ( x2 & ~x4 ) | ( x2 & x7 ) | ( ~x4 & x7 ) ;
  assign n157 = ( ~x3 & x7 ) | ( ~x3 & n156 ) | ( x7 & n156 ) ;
  assign n158 = x7 & ~n157 ;
  assign n159 = n157 | n158 ;
  assign n160 = ( ~x7 & n158 ) | ( ~x7 & n159 ) | ( n158 & n159 ) ;
  assign n161 = ( ~x0 & x5 ) | ( ~x0 & n160 ) | ( x5 & n160 ) ;
  assign n153 = x2 & x4 ;
  assign n154 = x3 | x7 ;
  assign n155 = ( x2 & ~n153 ) | ( x2 & n154 ) | ( ~n153 & n154 ) ;
  assign n162 = ( x0 & x5 ) | ( x0 & ~n155 ) | ( x5 & ~n155 ) ;
  assign n163 = n161 & n162 ;
  assign n149 = ( x2 & ~x5 ) | ( x2 & x7 ) | ( ~x5 & x7 ) ;
  assign n150 = ( x4 & ~x7 ) | ( x4 & n149 ) | ( ~x7 & n149 ) ;
  assign n151 = ( x2 & x4 ) | ( x2 & ~n149 ) | ( x4 & ~n149 ) ;
  assign n152 = n150 & ~n151 ;
  assign n164 = ( ~x0 & n152 ) | ( ~x0 & n163 ) | ( n152 & n163 ) ;
  assign n165 = x3 & ~n164 ;
  assign n166 = ( x3 & n163 ) | ( x3 & ~n165 ) | ( n163 & ~n165 ) ;
  assign n167 = ( x1 & ~x6 ) | ( x1 & n166 ) | ( ~x6 & n166 ) ;
  assign n142 = x2 & ~x3 ;
  assign n143 = ~x4 & n142 ;
  assign n144 = ( x0 & n9 ) | ( x0 & n143 ) | ( n9 & n143 ) ;
  assign n145 = ~x0 & n144 ;
  assign n138 = ( x2 & x4 ) | ( x2 & ~x7 ) | ( x4 & ~x7 ) ;
  assign n139 = ( ~x2 & x5 ) | ( ~x2 & n138 ) | ( x5 & n138 ) ;
  assign n140 = ( ~x5 & x7 ) | ( ~x5 & n138 ) | ( x7 & n138 ) ;
  assign n141 = n139 & n140 ;
  assign n146 = ( x0 & n141 ) | ( x0 & n145 ) | ( n141 & n145 ) ;
  assign n147 = x3 & ~n146 ;
  assign n148 = ( x3 & n145 ) | ( x3 & ~n147 ) | ( n145 & ~n147 ) ;
  assign n168 = ( x1 & x6 ) | ( x1 & n148 ) | ( x6 & n148 ) ;
  assign n169 = n167 & n168 ;
  assign n184 = x3 & n83 ;
  assign n185 = x2 & n184 ;
  assign n186 = n27 & n185 ;
  assign n187 = ( x4 & x5 ) | ( x4 & n186 ) | ( x5 & n186 ) ;
  assign n188 = ~x5 & n187 ;
  assign n172 = ( x1 & x2 ) | ( x1 & ~x6 ) | ( x2 & ~x6 ) ;
  assign n173 = ( x2 & x4 ) | ( x2 & ~n172 ) | ( x4 & ~n172 ) ;
  assign n174 = ( ~x1 & x4 ) | ( ~x1 & n172 ) | ( x4 & n172 ) ;
  assign n175 = n173 & ~n174 ;
  assign n176 = x0 | n175 ;
  assign n170 = ~x2 & x4 ;
  assign n171 = ~x6 & n170 ;
  assign n177 = ~x1 & n171 ;
  assign n178 = x0 & ~n177 ;
  assign n179 = n176 & ~n178 ;
  assign n180 = ( x5 & x7 ) | ( x5 & n179 ) | ( x7 & n179 ) ;
  assign n181 = ( x3 & ~x5 ) | ( x3 & n180 ) | ( ~x5 & n180 ) ;
  assign n182 = ( x3 & x7 ) | ( x3 & ~n180 ) | ( x7 & ~n180 ) ;
  assign n183 = n181 & ~n182 ;
  assign n194 = ( x1 & x4 ) | ( x1 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n195 = ( x1 & x4 ) | ( x1 & ~n194 ) | ( x4 & ~n194 ) ;
  assign n196 = ( x4 & x6 ) | ( x4 & n195 ) | ( x6 & n195 ) ;
  assign n197 = ( n67 & n194 ) | ( n67 & ~n196 ) | ( n194 & ~n196 ) ;
  assign n198 = x0 & n197 ;
  assign n189 = ( x1 & ~x4 ) | ( x1 & x6 ) | ( ~x4 & x6 ) ;
  assign n190 = ( ~x4 & x5 ) | ( ~x4 & x6 ) | ( x5 & x6 ) ;
  assign n191 = n189 & n190 ;
  assign n192 = x5 & ~n191 ;
  assign n193 = ( n189 & ~n191 ) | ( n189 & n192 ) | ( ~n191 & n192 ) ;
  assign n199 = x0 | n193 ;
  assign n200 = ( ~x0 & n198 ) | ( ~x0 & n199 ) | ( n198 & n199 ) ;
  assign n232 = ( x1 & x3 ) | ( x1 & x5 ) | ( x3 & x5 ) ;
  assign n227 = ( x0 & x4 ) | ( x0 & x6 ) | ( x4 & x6 ) ;
  assign n228 = ( ~x2 & x6 ) | ( ~x2 & n227 ) | ( x6 & n227 ) ;
  assign n229 = x6 & ~n228 ;
  assign n230 = n228 | n229 ;
  assign n231 = ( ~x6 & n229 ) | ( ~x6 & n230 ) | ( n229 & n230 ) ;
  assign n233 = x1 | x3 ;
  assign n234 = ( x5 & n231 ) | ( x5 & n233 ) | ( n231 & n233 ) ;
  assign n235 = ~n232 & n234 ;
  assign n218 = ( x3 & x5 ) | ( x3 & x6 ) | ( x5 & x6 ) ;
  assign n219 = ( ~x4 & x6 ) | ( ~x4 & n218 ) | ( x6 & n218 ) ;
  assign n220 = x6 & ~n219 ;
  assign n221 = n219 | n220 ;
  assign n222 = ( ~x6 & n220 ) | ( ~x6 & n221 ) | ( n220 & n221 ) ;
  assign n223 = x1 | n222 ;
  assign n217 = ~x6 & n55 ;
  assign n224 = ~x3 & n217 ;
  assign n225 = x1 & ~n224 ;
  assign n226 = n223 & ~n225 ;
  assign n236 = ( x0 & n226 ) | ( x0 & n235 ) | ( n226 & n235 ) ;
  assign n237 = x2 & ~n236 ;
  assign n238 = ( x2 & n235 ) | ( x2 & ~n237 ) | ( n235 & ~n237 ) ;
  assign n239 = ( x2 & n200 ) | ( x2 & n238 ) | ( n200 & n238 ) ;
  assign n203 = ~x1 & x5 ;
  assign n204 = ( x1 & ~x4 ) | ( x1 & x5 ) | ( ~x4 & x5 ) ;
  assign n205 = ( ~x4 & x5 ) | ( ~x4 & n67 ) | ( x5 & n67 ) ;
  assign n206 = ( n203 & n204 ) | ( n203 & ~n205 ) | ( n204 & ~n205 ) ;
  assign n207 = x1 & ~x6 ;
  assign n208 = ~x1 & x4 ;
  assign n209 = x4 & ~x6 ;
  assign n210 = ( n207 & n208 ) | ( n207 & ~n209 ) | ( n208 & ~n209 ) ;
  assign n211 = ( x0 & x5 ) | ( x0 & ~n210 ) | ( x5 & ~n210 ) ;
  assign n212 = x0 & ~n211 ;
  assign n213 = ( x5 & ~n211 ) | ( x5 & n212 ) | ( ~n211 & n212 ) ;
  assign n214 = ( ~x0 & n206 ) | ( ~x0 & n213 ) | ( n206 & n213 ) ;
  assign n201 = x1 & ~x4 ;
  assign n202 = ( x5 & n18 ) | ( x5 & n201 ) | ( n18 & n201 ) ;
  assign n215 = ( x0 & n202 ) | ( x0 & n213 ) | ( n202 & n213 ) ;
  assign n216 = n214 | n215 ;
  assign n240 = ( ~x2 & n216 ) | ( ~x2 & n238 ) | ( n216 & n238 ) ;
  assign n241 = n239 | n240 ;
  assign n242 = n183 | n241 ;
  assign n243 = ( ~n169 & n188 ) | ( ~n169 & n242 ) | ( n188 & n242 ) ;
  assign n244 = n169 | n243 ;
  assign n261 = ( x2 & x3 ) | ( x2 & x7 ) | ( x3 & x7 ) ;
  assign n262 = ( x3 & ~x5 ) | ( x3 & n261 ) | ( ~x5 & n261 ) ;
  assign n263 = x3 & ~n262 ;
  assign n264 = n262 | n263 ;
  assign n265 = ( ~x3 & n263 ) | ( ~x3 & n264 ) | ( n263 & n264 ) ;
  assign n266 = ( ~x1 & x4 ) | ( ~x1 & n265 ) | ( x4 & n265 ) ;
  assign n259 = ( x2 & x3 ) | ( x2 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n260 = n149 & ~n259 ;
  assign n267 = ( x1 & x4 ) | ( x1 & n260 ) | ( x4 & n260 ) ;
  assign n268 = n266 & n267 ;
  assign n269 = x2 | x7 ;
  assign n255 = ( x3 & ~x4 ) | ( x3 & n232 ) | ( ~x4 & n232 ) ;
  assign n256 = x3 & ~n255 ;
  assign n257 = n255 | n256 ;
  assign n258 = ( ~x3 & n256 ) | ( ~x3 & n257 ) | ( n256 & n257 ) ;
  assign n270 = ( x2 & x7 ) | ( x2 & ~n258 ) | ( x7 & ~n258 ) ;
  assign n271 = ( n268 & n269 ) | ( n268 & ~n270 ) | ( n269 & ~n270 ) ;
  assign n272 = x6 & ~n271 ;
  assign n246 = ( x3 & x5 ) | ( x3 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n247 = ( ~x1 & x5 ) | ( ~x1 & n246 ) | ( x5 & n246 ) ;
  assign n248 = ( x1 & ~x3 ) | ( x1 & n247 ) | ( ~x3 & n247 ) ;
  assign n249 = x7 | n248 ;
  assign n250 = ( ~x5 & n247 ) | ( ~x5 & n249 ) | ( n247 & n249 ) ;
  assign n251 = ~x2 & n250 ;
  assign n245 = x3 & n9 ;
  assign n252 = x1 & n245 ;
  assign n253 = x2 & ~n252 ;
  assign n254 = n251 | n253 ;
  assign n273 = x4 & ~n254 ;
  assign n274 = x6 | n273 ;
  assign n275 = ~n272 & n274 ;
  assign n306 = ( x0 & x5 ) | ( x0 & ~n218 ) | ( x5 & ~n218 ) ;
  assign n307 = ( ~x5 & x6 ) | ( ~x5 & n306 ) | ( x6 & n306 ) ;
  assign n308 = n218 | n307 ;
  assign n309 = ( ~x0 & n306 ) | ( ~x0 & n308 ) | ( n306 & n308 ) ;
  assign n310 = x2 & n309 ;
  assign n304 = x3 & ~x6 ;
  assign n305 = x5 & n304 ;
  assign n311 = x0 & n305 ;
  assign n312 = x2 | n311 ;
  assign n313 = ~n310 & n312 ;
  assign n341 = ( x1 & x2 ) | ( x1 & x6 ) | ( x2 & x6 ) ;
  assign n342 = ~x2 & x5 ;
  assign n343 = x6 & n341 ;
  assign n344 = ( x1 & x5 ) | ( x1 & n343 ) | ( x5 & n343 ) ;
  assign n345 = ( n341 & n342 ) | ( n341 & ~n344 ) | ( n342 & ~n344 ) ;
  assign n346 = x4 | n345 ;
  assign n347 = n19 & n67 ;
  assign n348 = x4 & ~n347 ;
  assign n349 = n346 & ~n348 ;
  assign n361 = x3 & n349 ;
  assign n354 = x2 | x6 ;
  assign n355 = ( ~x2 & x5 ) | ( ~x2 & n354 ) | ( x5 & n354 ) ;
  assign n356 = ( ~x4 & x5 ) | ( ~x4 & n354 ) | ( x5 & n354 ) ;
  assign n357 = ( n170 & ~n355 ) | ( n170 & n356 ) | ( ~n355 & n356 ) ;
  assign n358 = x1 & n357 ;
  assign n350 = ( x2 & x4 ) | ( x2 & x6 ) | ( x4 & x6 ) ;
  assign n351 = ( x4 & x5 ) | ( x4 & x6 ) | ( x5 & x6 ) ;
  assign n352 = x2 | n351 ;
  assign n353 = ~n350 & n352 ;
  assign n359 = x1 | n353 ;
  assign n360 = ( ~x1 & n358 ) | ( ~x1 & n359 ) | ( n358 & n359 ) ;
  assign n362 = x3 | n360 ;
  assign n363 = ( ~x3 & n361 ) | ( ~x3 & n362 ) | ( n361 & n362 ) ;
  assign n364 = x0 & n363 ;
  assign n323 = ( x3 & ~x4 ) | ( x3 & x6 ) | ( ~x4 & x6 ) ;
  assign n324 = ( x3 & ~x5 ) | ( x3 & n323 ) | ( ~x5 & n323 ) ;
  assign n325 = x3 & ~n324 ;
  assign n326 = n324 | n325 ;
  assign n327 = ( ~x3 & n325 ) | ( ~x3 & n326 ) | ( n325 & n326 ) ;
  assign n331 = ( x1 & x2 ) | ( x1 & ~n327 ) | ( x2 & ~n327 ) ;
  assign n328 = x4 & n67 ;
  assign n329 = ( x1 & x3 ) | ( x1 & n328 ) | ( x3 & n328 ) ;
  assign n330 = ~x1 & n329 ;
  assign n332 = x2 & n330 ;
  assign n333 = ( n327 & n331 ) | ( n327 & n332 ) | ( n331 & n332 ) ;
  assign n334 = x4 | n190 ;
  assign n335 = ( ~x6 & n190 ) | ( ~x6 & n334 ) | ( n190 & n334 ) ;
  assign n336 = x1 & x2 ;
  assign n337 = x2 & ~n336 ;
  assign n338 = ~n335 & n337 ;
  assign n339 = ( n217 & ~n336 ) | ( n217 & n337 ) | ( ~n336 & n337 ) ;
  assign n340 = ( x1 & n338 ) | ( x1 & n339 ) | ( n338 & n339 ) ;
  assign n365 = n333 | n340 ;
  assign n366 = ~x0 & n365 ;
  assign n367 = n364 | n366 ;
  assign n368 = ( x1 & n313 ) | ( x1 & n367 ) | ( n313 & n367 ) ;
  assign n316 = ( ~x2 & x6 ) | ( ~x2 & n142 ) | ( x6 & n142 ) ;
  assign n317 = ( x0 & x6 ) | ( x0 & n142 ) | ( x6 & n142 ) ;
  assign n318 = ( n34 & n316 ) | ( n34 & ~n317 ) | ( n316 & ~n317 ) ;
  assign n319 = x5 | n318 ;
  assign n314 = ~x3 & x6 ;
  assign n315 = ( ~x2 & x6 ) | ( ~x2 & n314 ) | ( x6 & n314 ) ;
  assign n320 = ~x0 & n315 ;
  assign n321 = x5 & ~n320 ;
  assign n322 = n319 & ~n321 ;
  assign n369 = ( ~x1 & n322 ) | ( ~x1 & n367 ) | ( n322 & n367 ) ;
  assign n370 = n368 | n369 ;
  assign n371 = ( x0 & n275 ) | ( x0 & n370 ) | ( n275 & n370 ) ;
  assign n286 = ( ~x2 & x3 ) | ( ~x2 & x7 ) | ( x3 & x7 ) ;
  assign n287 = ( x2 & x5 ) | ( x2 & ~n286 ) | ( x5 & ~n286 ) ;
  assign n288 = ( ~x5 & x7 ) | ( ~x5 & n287 ) | ( x7 & n287 ) ;
  assign n289 = x3 & n288 ;
  assign n290 = ( ~x2 & n287 ) | ( ~x2 & n289 ) | ( n287 & n289 ) ;
  assign n291 = ( x6 & n9 ) | ( x6 & n142 ) | ( n9 & n142 ) ;
  assign n292 = ~x6 & n291 ;
  assign n293 = x6 | n292 ;
  assign n294 = ( n290 & n292 ) | ( n290 & n293 ) | ( n292 & n293 ) ;
  assign n298 = ( ~x1 & x4 ) | ( ~x1 & n294 ) | ( x4 & n294 ) ;
  assign n295 = ~x5 & n142 ;
  assign n296 = ( x1 & n27 ) | ( x1 & n295 ) | ( n27 & n295 ) ;
  assign n297 = ~x1 & n296 ;
  assign n299 = ~x4 & n297 ;
  assign n300 = ( n294 & ~n298 ) | ( n294 & n299 ) | ( ~n298 & n299 ) ;
  assign n301 = x6 | x7 ;
  assign n276 = x2 & x3 ;
  assign n277 = ( ~x1 & x4 ) | ( ~x1 & n276 ) | ( x4 & n276 ) ;
  assign n278 = x4 | n277 ;
  assign n279 = x4 & n277 ;
  assign n280 = n278 & ~n279 ;
  assign n281 = x1 & ~x5 ;
  assign n282 = ( x2 & x4 ) | ( x2 & n281 ) | ( x4 & n281 ) ;
  assign n283 = ~x2 & n282 ;
  assign n284 = x5 | n283 ;
  assign n285 = ( n280 & n283 ) | ( n280 & n284 ) | ( n283 & n284 ) ;
  assign n302 = ( x6 & x7 ) | ( x6 & ~n285 ) | ( x7 & ~n285 ) ;
  assign n303 = ( n300 & n301 ) | ( n300 & ~n302 ) | ( n301 & ~n302 ) ;
  assign n372 = ( ~x0 & n303 ) | ( ~x0 & n370 ) | ( n303 & n370 ) ;
  assign n373 = n371 | n372 ;
  assign n375 = ( x1 & ~x4 ) | ( x1 & x7 ) | ( ~x4 & x7 ) ;
  assign n376 = ( x2 & x4 ) | ( x2 & n375 ) | ( x4 & n375 ) ;
  assign n377 = ( x4 & x7 ) | ( x4 & ~n376 ) | ( x7 & ~n376 ) ;
  assign n378 = n375 & n377 ;
  assign n379 = ( x2 & ~n376 ) | ( x2 & n378 ) | ( ~n376 & n378 ) ;
  assign n380 = x3 & ~n379 ;
  assign n374 = x4 & x7 ;
  assign n381 = n19 & n374 ;
  assign n382 = x3 | n381 ;
  assign n383 = ~n380 & n382 ;
  assign n384 = ( x0 & x5 ) | ( x0 & ~n383 ) | ( x5 & ~n383 ) ;
  assign n385 = x0 & ~n384 ;
  assign n386 = ( x5 & ~n384 ) | ( x5 & n385 ) | ( ~n384 & n385 ) ;
  assign n397 = ( ~x2 & x5 ) | ( ~x2 & x7 ) | ( x5 & x7 ) ;
  assign n398 = ( x1 & x7 ) | ( x1 & ~n397 ) | ( x7 & ~n397 ) ;
  assign n399 = ( x2 & ~x5 ) | ( x2 & n398 ) | ( ~x5 & n398 ) ;
  assign n400 = n397 & n399 ;
  assign n401 = ( ~n398 & n399 ) | ( ~n398 & n400 ) | ( n399 & n400 ) ;
  assign n402 = ~x4 & n401 ;
  assign n403 = ~x0 & n402 ;
  assign n396 = ~x7 & n121 ;
  assign n404 = n396 | n403 ;
  assign n405 = ( n35 & n403 ) | ( n35 & n404 ) | ( n403 & n404 ) ;
  assign n406 = ( x3 & x6 ) | ( x3 & ~n405 ) | ( x6 & ~n405 ) ;
  assign n407 = x3 & ~n406 ;
  assign n408 = ( x6 & ~n406 ) | ( x6 & n407 ) | ( ~n406 & n407 ) ;
  assign n388 = x1 & ~x2 ;
  assign n457 = x0 & ~x2 ;
  assign n458 = ( n94 & ~n388 ) | ( n94 & n457 ) | ( ~n388 & n457 ) ;
  assign n459 = ( x5 & x7 ) | ( x5 & n458 ) | ( x7 & n458 ) ;
  assign n460 = ( x6 & ~x7 ) | ( x6 & n459 ) | ( ~x7 & n459 ) ;
  assign n461 = ( x5 & x6 ) | ( x5 & ~n459 ) | ( x6 & ~n459 ) ;
  assign n462 = n460 & ~n461 ;
  assign n453 = ( x2 & ~x6 ) | ( x2 & x7 ) | ( ~x6 & x7 ) ;
  assign n454 = ( x1 & ~x7 ) | ( x1 & n453 ) | ( ~x7 & n453 ) ;
  assign n455 = ( x1 & x2 ) | ( x1 & ~n453 ) | ( x2 & ~n453 ) ;
  assign n456 = n454 & ~n455 ;
  assign n463 = ( x0 & n456 ) | ( x0 & n462 ) | ( n456 & n462 ) ;
  assign n464 = x5 & ~n463 ;
  assign n465 = ( x5 & n462 ) | ( x5 & ~n464 ) | ( n462 & ~n464 ) ;
  assign n466 = x4 | n465 ;
  assign n444 = ~x1 & x7 ;
  assign n445 = ( ~x5 & x6 ) | ( ~x5 & n444 ) | ( x6 & n444 ) ;
  assign n446 = ( x6 & x7 ) | ( x6 & ~n444 ) | ( x7 & ~n444 ) ;
  assign n447 = ( x1 & x5 ) | ( x1 & ~n446 ) | ( x5 & ~n446 ) ;
  assign n448 = n445 | n447 ;
  assign n449 = x2 & n448 ;
  assign n441 = ( x5 & x6 ) | ( x5 & x7 ) | ( x6 & x7 ) ;
  assign n442 = x5 & ~n441 ;
  assign n443 = ( x7 & ~n441 ) | ( x7 & n442 ) | ( ~n441 & n442 ) ;
  assign n450 = x1 & n443 ;
  assign n451 = x2 | n450 ;
  assign n452 = ~n449 & n451 ;
  assign n467 = x0 & n452 ;
  assign n468 = x4 & ~n467 ;
  assign n469 = n466 & ~n468 ;
  assign n470 = x3 | n469 ;
  assign n425 = ( x5 & x7 ) | ( x5 & ~n208 ) | ( x7 & ~n208 ) ;
  assign n426 = x4 & n425 ;
  assign n427 = ( ~x5 & n208 ) | ( ~x5 & n426 ) | ( n208 & n426 ) ;
  assign n428 = ( ~x1 & n425 ) | ( ~x1 & n427 ) | ( n425 & n427 ) ;
  assign n429 = ( ~x7 & n426 ) | ( ~x7 & n428 ) | ( n426 & n428 ) ;
  assign n430 = x2 | n429 ;
  assign n422 = ( x4 & x5 ) | ( x4 & x7 ) | ( x5 & x7 ) ;
  assign n423 = x4 & ~n422 ;
  assign n424 = ( x5 & ~n422 ) | ( x5 & n423 ) | ( ~n422 & n423 ) ;
  assign n431 = ~x1 & n424 ;
  assign n432 = x2 & ~n431 ;
  assign n433 = n430 & ~n432 ;
  assign n434 = x5 | x7 ;
  assign n435 = x6 | n434 ;
  assign n436 = x1 & x4 ;
  assign n437 = ( x2 & ~n435 ) | ( x2 & n436 ) | ( ~n435 & n436 ) ;
  assign n438 = ~x2 & n437 ;
  assign n439 = x6 | n438 ;
  assign n440 = ( n433 & n438 ) | ( n433 & n439 ) | ( n438 & n439 ) ;
  assign n471 = x0 & n440 ;
  assign n472 = x3 & ~n471 ;
  assign n473 = n470 & ~n472 ;
  assign n411 = ( ~x2 & x3 ) | ( ~x2 & x5 ) | ( x3 & x5 ) ;
  assign n412 = ( x2 & ~x3 ) | ( x2 & x6 ) | ( ~x3 & x6 ) ;
  assign n413 = n411 & n412 ;
  assign n414 = x1 & ~n413 ;
  assign n409 = x3 & ~x5 ;
  assign n410 = ~x6 & n409 ;
  assign n415 = ~x2 & n410 ;
  assign n416 = x1 | n415 ;
  assign n417 = ~n414 & n416 ;
  assign n418 = ( ~x0 & x7 ) | ( ~x0 & n417 ) | ( x7 & n417 ) ;
  assign n419 = ( x4 & ~x7 ) | ( x4 & n418 ) | ( ~x7 & n418 ) ;
  assign n420 = ( x0 & ~x4 ) | ( x0 & n418 ) | ( ~x4 & n418 ) ;
  assign n421 = n419 & n420 ;
  assign n479 = x4 & ~n435 ;
  assign n480 = ( x0 & x3 ) | ( x0 & n479 ) | ( x3 & n479 ) ;
  assign n481 = ~x0 & n480 ;
  assign n474 = ( x0 & ~x3 ) | ( x0 & x6 ) | ( ~x3 & x6 ) ;
  assign n475 = ( x0 & x5 ) | ( x0 & ~n474 ) | ( x5 & ~n474 ) ;
  assign n476 = ( x3 & ~x6 ) | ( x3 & n475 ) | ( ~x6 & n475 ) ;
  assign n477 = n474 & n476 ;
  assign n478 = ( ~n475 & n476 ) | ( ~n475 & n477 ) | ( n476 & n477 ) ;
  assign n482 = ( ~x4 & n478 ) | ( ~x4 & n481 ) | ( n478 & n481 ) ;
  assign n483 = x7 & ~n482 ;
  assign n484 = ( x7 & n481 ) | ( x7 & ~n483 ) | ( n481 & ~n483 ) ;
  assign n485 = x0 & x3 ;
  assign n486 = ( x2 & n38 ) | ( x2 & n485 ) | ( n38 & n485 ) ;
  assign n487 = ~x2 & n486 ;
  assign n488 = x2 | n487 ;
  assign n489 = ( n484 & n487 ) | ( n484 & n488 ) | ( n487 & n488 ) ;
  assign n490 = n421 | n489 ;
  assign n491 = ( ~n408 & n473 ) | ( ~n408 & n490 ) | ( n473 & n490 ) ;
  assign n492 = n408 | n491 ;
  assign n387 = ~x7 & n201 ;
  assign n389 = ( ~x1 & x2 ) | ( ~x1 & n201 ) | ( x2 & n201 ) ;
  assign n390 = ( x7 & n388 ) | ( x7 & n389 ) | ( n388 & n389 ) ;
  assign n391 = ( x7 & n387 ) | ( x7 & ~n390 ) | ( n387 & ~n390 ) ;
  assign n392 = ( x3 & x5 ) | ( x3 & n391 ) | ( x5 & n391 ) ;
  assign n393 = ( x0 & ~x5 ) | ( x0 & n392 ) | ( ~x5 & n392 ) ;
  assign n394 = ( x0 & x3 ) | ( x0 & ~n392 ) | ( x3 & ~n392 ) ;
  assign n395 = n393 & ~n394 ;
  assign n510 = ( x1 & ~x2 ) | ( x1 & x7 ) | ( ~x2 & x7 ) ;
  assign n511 = x2 & ~x7 ;
  assign n512 = ( x1 & x5 ) | ( x1 & ~n511 ) | ( x5 & ~n511 ) ;
  assign n513 = ~n510 & n512 ;
  assign n518 = x0 & n513 ;
  assign n514 = x2 & x7 ;
  assign n515 = x1 | x5 ;
  assign n516 = x7 & n515 ;
  assign n517 = ( n388 & n514 ) | ( n388 & ~n516 ) | ( n514 & ~n516 ) ;
  assign n519 = x0 | n517 ;
  assign n520 = ( ~x0 & n518 ) | ( ~x0 & n519 ) | ( n518 & n519 ) ;
  assign n521 = x4 & ~n520 ;
  assign n507 = x7 & ~n397 ;
  assign n508 = ( x1 & x2 ) | ( x1 & ~n507 ) | ( x2 & ~n507 ) ;
  assign n509 = ( n397 & ~n507 ) | ( n397 & n508 ) | ( ~n507 & n508 ) ;
  assign n522 = x0 & ~n509 ;
  assign n523 = x4 | n522 ;
  assign n524 = ~n521 & n523 ;
  assign n528 = ( x0 & x3 ) | ( x0 & x5 ) | ( x3 & x5 ) ;
  assign n529 = ( ~x4 & x5 ) | ( ~x4 & n528 ) | ( x5 & n528 ) ;
  assign n530 = x5 & ~n529 ;
  assign n531 = n529 | n530 ;
  assign n532 = ( ~x5 & n530 ) | ( ~x5 & n531 ) | ( n530 & n531 ) ;
  assign n533 = ~x7 & n532 ;
  assign n534 = x1 & ~n533 ;
  assign n525 = x4 & x5 ;
  assign n526 = ( x3 & x7 ) | ( x3 & ~n525 ) | ( x7 & ~n525 ) ;
  assign n527 = n57 & n526 ;
  assign n535 = ~x0 & n527 ;
  assign n536 = x1 | n535 ;
  assign n537 = ~n534 & n536 ;
  assign n538 = ( x3 & n524 ) | ( x3 & n537 ) | ( n524 & n537 ) ;
  assign n495 = ( x1 & ~x5 ) | ( x1 & n397 ) | ( ~x5 & n397 ) ;
  assign n496 = ( ~x2 & x7 ) | ( ~x2 & n495 ) | ( x7 & n495 ) ;
  assign n497 = ~n397 & n496 ;
  assign n498 = ( ~n495 & n496 ) | ( ~n495 & n497 ) | ( n496 & n497 ) ;
  assign n499 = x4 & ~n498 ;
  assign n493 = x1 | x2 ;
  assign n494 = ~x5 & x7 ;
  assign n500 = ~n493 & n494 ;
  assign n501 = x4 | n500 ;
  assign n502 = ~n499 & n501 ;
  assign n503 = x0 | n502 ;
  assign n504 = n396 & ~n493 ;
  assign n505 = x0 & ~n504 ;
  assign n506 = n503 & ~n505 ;
  assign n539 = ( ~x3 & n506 ) | ( ~x3 & n537 ) | ( n506 & n537 ) ;
  assign n540 = n538 | n539 ;
  assign n541 = n395 | n540 ;
  assign n542 = ( ~n386 & n492 ) | ( ~n386 & n541 ) | ( n492 & n541 ) ;
  assign n543 = n386 | n542 ;
  assign y0 = n54 ;
  assign y1 = n137 ;
  assign y2 = n244 ;
  assign y3 = n373 ;
  assign y4 = n543 ;
endmodule
