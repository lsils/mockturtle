module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 , G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G4 , G5 , G6 , G7 , G8 , G9 ;
  output G1884 , G1885 , G1886 , G1887 , G1888 , G1889 , G1890 , G1891 , G1892 , G1893 , G1894 , G1895 , G1896 , G1897 , G1898 , G1899 , G1900 , G1901 , G1902 , G1903 , G1904 , G1905 , G1906 , G1907 , G1908 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 ;
  assign n34 = G24 | G31 ;
  assign n35 = G18 & n34 ;
  assign n36 = G6 | G7 ;
  assign n37 = G6 & G7 ;
  assign n38 = n36 & ~n37 ;
  assign n39 = G5 & n38 ;
  assign n40 = G5 | n38 ;
  assign n41 = ~n39 & n40 ;
  assign n42 = G4 | G8 ;
  assign n43 = G4 & G8 ;
  assign n44 = n42 & ~n43 ;
  assign n45 = G2 | G3 ;
  assign n46 = G2 & G3 ;
  assign n47 = n45 & ~n46 ;
  assign n48 = G1 & n47 ;
  assign n49 = G1 | n47 ;
  assign n50 = ~n48 & n49 ;
  assign n51 = ~n44 & n50 ;
  assign n52 = n44 & ~n50 ;
  assign n53 = n51 | n52 ;
  assign n54 = n41 | n53 ;
  assign n55 = n41 & n53 ;
  assign n56 = n54 & ~n55 ;
  assign n57 = G21 & ~G33 ;
  assign n58 = ~G9 & n57 ;
  assign n59 = G9 & ~n57 ;
  assign n60 = n58 | n59 ;
  assign n61 = G10 & ~G15 ;
  assign n62 = ~G10 & G15 ;
  assign n63 = n61 | n62 ;
  assign n64 = ~G16 & n63 ;
  assign n65 = G16 & ~n63 ;
  assign n66 = n64 | n65 ;
  assign n67 = ~n60 & n66 ;
  assign n68 = n60 & ~n66 ;
  assign n69 = n67 | n68 ;
  assign n70 = n56 & ~n69 ;
  assign n71 = ~n56 & n69 ;
  assign n72 = n70 | n71 ;
  assign n73 = G31 | n72 ;
  assign n74 = G17 & n34 ;
  assign n75 = n73 & ~n74 ;
  assign n76 = ~n73 & n74 ;
  assign n77 = n75 | n76 ;
  assign n78 = n35 & ~n77 ;
  assign n79 = ~G11 & G13 ;
  assign n80 = G11 & ~G13 ;
  assign n81 = n79 | n80 ;
  assign n82 = G12 & ~n81 ;
  assign n83 = ~G12 & n81 ;
  assign n84 = n82 | n83 ;
  assign n85 = ~n66 & n84 ;
  assign n86 = n66 & ~n84 ;
  assign n87 = n85 | n86 ;
  assign n88 = G24 | G33 ;
  assign n89 = G17 & ~n88 ;
  assign n90 = ~G1 & n89 ;
  assign n91 = G1 & ~n89 ;
  assign n92 = n90 | n91 ;
  assign n93 = n41 | n92 ;
  assign n94 = n41 & n92 ;
  assign n95 = n93 & ~n94 ;
  assign n96 = n87 | n95 ;
  assign n97 = n87 & n95 ;
  assign n98 = n96 & ~n97 ;
  assign n99 = G31 | n98 ;
  assign n100 = G26 | n99 ;
  assign n101 = G26 & n99 ;
  assign n102 = n100 & ~n101 ;
  assign n103 = ~G14 & G9 ;
  assign n104 = G14 & ~G9 ;
  assign n105 = n103 | n104 ;
  assign n106 = ~G16 & n105 ;
  assign n107 = G16 & ~n105 ;
  assign n108 = n106 | n107 ;
  assign n109 = G23 | G33 ;
  assign n110 = G20 & ~n109 ;
  assign n111 = ~G13 & n110 ;
  assign n112 = G13 & ~n110 ;
  assign n113 = n111 | n112 ;
  assign n114 = ~n108 & n113 ;
  assign n115 = n108 & ~n113 ;
  assign n116 = n114 | n115 ;
  assign n117 = G4 & ~G7 ;
  assign n118 = ~G4 & G7 ;
  assign n119 = n117 | n118 ;
  assign n120 = G10 & ~n119 ;
  assign n121 = ~G10 & n119 ;
  assign n122 = n120 | n121 ;
  assign n123 = n116 & n122 ;
  assign n124 = n116 | n122 ;
  assign n125 = ~n123 & n124 ;
  assign n126 = G31 | n125 ;
  assign n127 = G23 | G31 ;
  assign n128 = G19 & n127 ;
  assign n129 = n126 & n128 ;
  assign n130 = n126 | n128 ;
  assign n131 = ~n129 & n130 ;
  assign n132 = n102 & n131 ;
  assign n133 = G18 & ~n88 ;
  assign n134 = G11 | G15 ;
  assign n135 = G11 & G15 ;
  assign n136 = n134 & ~n135 ;
  assign n137 = n133 | n136 ;
  assign n138 = n133 & n136 ;
  assign n139 = n137 & ~n138 ;
  assign n140 = n108 & n139 ;
  assign n141 = n108 | n139 ;
  assign n142 = ~n140 & n141 ;
  assign n143 = G5 & ~G8 ;
  assign n144 = ~G5 & G8 ;
  assign n145 = n143 | n144 ;
  assign n146 = G2 & ~n145 ;
  assign n147 = ~G2 & n145 ;
  assign n148 = n146 | n147 ;
  assign n149 = ~n142 & n148 ;
  assign n150 = n142 & ~n148 ;
  assign n151 = n149 | n150 ;
  assign n152 = ~G31 & n151 ;
  assign n153 = G27 & n152 ;
  assign n154 = G27 | n152 ;
  assign n155 = ~n153 & n154 ;
  assign n156 = G3 | G6 ;
  assign n157 = G3 & G6 ;
  assign n158 = n156 & ~n157 ;
  assign n159 = G8 & n158 ;
  assign n160 = G8 | n158 ;
  assign n161 = ~n159 & n160 ;
  assign n162 = G19 & ~n109 ;
  assign n163 = G12 & n63 ;
  assign n164 = G12 | n63 ;
  assign n165 = ~n163 & n164 ;
  assign n166 = n162 & ~n165 ;
  assign n167 = ~n162 & n165 ;
  assign n168 = n166 | n167 ;
  assign n169 = n161 | n168 ;
  assign n170 = n161 & n168 ;
  assign n171 = n169 & ~n170 ;
  assign n172 = ~G31 & n171 ;
  assign n173 = G28 & n172 ;
  assign n174 = G28 | n172 ;
  assign n175 = ~n173 & n174 ;
  assign n176 = n155 | n175 ;
  assign n177 = n132 & ~n176 ;
  assign n178 = G20 & n127 ;
  assign n179 = G22 & ~G33 ;
  assign n180 = ~G14 & G4 ;
  assign n181 = G14 & ~G4 ;
  assign n182 = n180 | n181 ;
  assign n183 = n179 & ~n182 ;
  assign n184 = ~n179 & n182 ;
  assign n185 = n183 | n184 ;
  assign n186 = n50 | n185 ;
  assign n187 = n50 & n185 ;
  assign n188 = n186 & ~n187 ;
  assign n189 = n87 | n188 ;
  assign n190 = n87 & n188 ;
  assign n191 = n189 & ~n190 ;
  assign n192 = ~G31 & n191 ;
  assign n193 = G25 | n192 ;
  assign n194 = G25 & n192 ;
  assign n195 = n193 & ~n194 ;
  assign n196 = n178 & n195 ;
  assign n197 = n177 & ~n196 ;
  assign n198 = ~n78 & n197 ;
  assign n199 = G29 | G33 ;
  assign n200 = ~G23 & G24 ;
  assign n201 = G31 | n200 ;
  assign n202 = n199 | n201 ;
  assign n203 = G32 | G33 ;
  assign n204 = n200 | n203 ;
  assign n205 = n202 & n204 ;
  assign n206 = n198 & ~n205 ;
  assign n207 = G1 | n206 ;
  assign n208 = G1 & n206 ;
  assign n209 = n207 & ~n208 ;
  assign n210 = G2 | n206 ;
  assign n211 = G2 & n206 ;
  assign n212 = n210 & ~n211 ;
  assign n213 = G3 | n206 ;
  assign n214 = G3 & n206 ;
  assign n215 = n213 & ~n214 ;
  assign n216 = G4 | n206 ;
  assign n217 = G4 & n206 ;
  assign n218 = n216 & ~n217 ;
  assign n219 = G30 | G33 ;
  assign n220 = n201 | n219 ;
  assign n221 = n204 & n220 ;
  assign n222 = n198 & ~n221 ;
  assign n223 = G10 | n222 ;
  assign n224 = G10 & n222 ;
  assign n225 = n223 & ~n224 ;
  assign n226 = G15 | n222 ;
  assign n227 = G15 & n222 ;
  assign n228 = n226 & ~n227 ;
  assign n229 = G16 | n222 ;
  assign n230 = G16 & n222 ;
  assign n231 = n229 & ~n230 ;
  assign n232 = n178 & ~n195 ;
  assign n233 = n177 & n232 ;
  assign n234 = ~n78 & n233 ;
  assign n235 = ~n205 & n234 ;
  assign n236 = G5 | n235 ;
  assign n237 = G5 & n235 ;
  assign n238 = n236 & ~n237 ;
  assign n239 = G6 | n235 ;
  assign n240 = G6 & n235 ;
  assign n241 = n239 & ~n240 ;
  assign n242 = G7 | n235 ;
  assign n243 = G7 & n235 ;
  assign n244 = n242 & ~n243 ;
  assign n245 = G8 | n235 ;
  assign n246 = G8 & n235 ;
  assign n247 = n245 & ~n246 ;
  assign n248 = ~n221 & n234 ;
  assign n249 = G9 & ~n248 ;
  assign n250 = ~G9 & n248 ;
  assign n251 = n249 | n250 ;
  assign n252 = n35 & n197 ;
  assign n253 = n77 & n252 ;
  assign n254 = ~n221 & n253 ;
  assign n255 = G11 | n254 ;
  assign n256 = G11 & n254 ;
  assign n257 = n255 & ~n256 ;
  assign n258 = G12 | n254 ;
  assign n259 = G12 & n254 ;
  assign n260 = n258 & ~n259 ;
  assign n261 = G13 | n254 ;
  assign n262 = G13 & n254 ;
  assign n263 = n261 & ~n262 ;
  assign n264 = G14 | n254 ;
  assign n265 = G14 & n254 ;
  assign n266 = n264 & ~n265 ;
  assign n267 = n206 | n222 ;
  assign n268 = G32 & n267 ;
  assign n269 = n35 | n178 ;
  assign n270 = n195 | n269 ;
  assign n271 = n77 & ~n270 ;
  assign n272 = n177 & n271 ;
  assign n273 = G33 | n272 ;
  assign n274 = n268 | n273 ;
  assign n275 = n74 & n267 ;
  assign n276 = ~G31 & n275 ;
  assign n277 = n72 & ~n276 ;
  assign n278 = ~n73 & n275 ;
  assign n279 = n203 & ~n278 ;
  assign n280 = ~n277 & n279 ;
  assign n281 = G25 & n267 ;
  assign n282 = ~G31 & n281 ;
  assign n283 = n191 | n282 ;
  assign n284 = n192 & n281 ;
  assign n285 = n203 & ~n284 ;
  assign n286 = n283 & n285 ;
  assign n287 = G27 & ~G31 ;
  assign n288 = n267 & n287 ;
  assign n289 = n151 & ~n288 ;
  assign n290 = n203 & ~n289 ;
  assign n291 = G28 & ~G31 ;
  assign n292 = n267 & n291 ;
  assign n293 = n171 & ~n292 ;
  assign n294 = n203 & ~n293 ;
  assign n295 = ~G31 & n128 ;
  assign n296 = n267 & n295 ;
  assign n297 = n125 | n296 ;
  assign n298 = n203 & n297 ;
  assign n299 = n56 & n199 ;
  assign n300 = G21 & G29 ;
  assign n301 = n206 | n300 ;
  assign n302 = n206 & n300 ;
  assign n303 = n301 & ~n302 ;
  assign n304 = G33 | n303 ;
  assign n305 = n299 & n304 ;
  assign n306 = n299 | n304 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = n87 | n105 ;
  assign n309 = n87 & n105 ;
  assign n310 = n219 & ~n309 ;
  assign n311 = n308 & n310 ;
  assign n312 = G22 & G30 ;
  assign n313 = n222 | n312 ;
  assign n314 = n222 & n312 ;
  assign n315 = n313 & ~n314 ;
  assign n316 = G33 | n315 ;
  assign n317 = n311 & ~n316 ;
  assign n318 = ~n311 & n316 ;
  assign n319 = n317 | n318 ;
  assign n320 = G26 & n267 ;
  assign n321 = ~n98 & n203 ;
  assign n322 = ~n320 & n321 ;
  assign G1884 = ~n209 ;
  assign G1885 = ~n212 ;
  assign G1886 = ~n215 ;
  assign G1887 = ~n218 ;
  assign G1888 = ~n225 ;
  assign G1889 = ~n228 ;
  assign G1890 = ~n231 ;
  assign G1891 = ~n238 ;
  assign G1892 = ~n241 ;
  assign G1893 = ~n244 ;
  assign G1894 = ~n247 ;
  assign G1895 = ~n251 ;
  assign G1896 = ~n257 ;
  assign G1897 = ~n260 ;
  assign G1898 = ~n263 ;
  assign G1899 = ~n266 ;
  assign G1900 = n274 ;
  assign G1901 = n280 ;
  assign G1902 = n286 ;
  assign G1903 = n290 ;
  assign G1904 = n294 ;
  assign G1905 = n298 ;
  assign G1906 = ~n307 ;
  assign G1907 = ~n319 ;
  assign G1908 = n322 ;
endmodule
