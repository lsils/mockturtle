module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 ;
  wire n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 ;
  assign n27 = ( x12 & x14 ) | ( x12 & ~x15 ) | ( x14 & ~x15 ) ;
  assign n28 = ~x12 & x13 ;
  assign n29 = ( x14 & ~n27 ) | ( x14 & n28 ) | ( ~n27 & n28 ) ;
  assign n30 = ~x10 & n29 ;
  assign n31 = ( x9 & ~x11 ) | ( x9 & n30 ) | ( ~x11 & n30 ) ;
  assign n32 = ~x9 & n31 ;
  assign n33 = x16 | n32 ;
  assign n48 = x0 & ~x19 ;
  assign n49 = x15 & ~x22 ;
  assign n50 = ( ~x0 & n48 ) | ( ~x0 & n49 ) | ( n48 & n49 ) ;
  assign n51 = ( x19 & x24 ) | ( x19 & n50 ) | ( x24 & n50 ) ;
  assign n42 = x0 & x8 ;
  assign n43 = x3 & n42 ;
  assign n52 = n43 & n50 ;
  assign n53 = ( ~x24 & n51 ) | ( ~x24 & n52 ) | ( n51 & n52 ) ;
  assign n70 = x18 & ~n53 ;
  assign n54 = x0 | x21 ;
  assign n55 = ~x19 & n54 ;
  assign n56 = ( x18 & n54 ) | ( x18 & n55 ) | ( n54 & n55 ) ;
  assign n34 = ~x1 & x9 ;
  assign n35 = ( ~x2 & x10 ) | ( ~x2 & x11 ) | ( x10 & x11 ) ;
  assign n36 = ~x12 & n35 ;
  assign n37 = ( ~x2 & x12 ) | ( ~x2 & n36 ) | ( x12 & n36 ) ;
  assign n38 = x9 | n37 ;
  assign n57 = ( ~n34 & n38 ) | ( ~n34 & n56 ) | ( n38 & n56 ) ;
  assign n58 = x24 | n57 ;
  assign n59 = ( ~x24 & n56 ) | ( ~x24 & n58 ) | ( n56 & n58 ) ;
  assign n60 = ~x3 & x25 ;
  assign n61 = x8 & ~x19 ;
  assign n62 = ( x3 & n60 ) | ( x3 & n61 ) | ( n60 & n61 ) ;
  assign n63 = x0 & ~x8 ;
  assign n64 = ( x0 & ~x3 ) | ( x0 & n63 ) | ( ~x3 & n63 ) ;
  assign n65 = x24 | n64 ;
  assign n66 = ( ~n62 & n64 ) | ( ~n62 & n65 ) | ( n64 & n65 ) ;
  assign n67 = ~x21 & n66 ;
  assign n68 = x25 | n67 ;
  assign n69 = ( x22 & n67 ) | ( x22 & n68 ) | ( n67 & n68 ) ;
  assign n71 = n59 & ~n69 ;
  assign n72 = ( n53 & n70 ) | ( n53 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ( x21 & x25 ) | ( x21 & n72 ) | ( x25 & n72 ) ;
  assign n39 = ( x0 & x19 ) | ( x0 & n34 ) | ( x19 & n34 ) ;
  assign n40 = n38 & n39 ;
  assign n41 = ( x19 & ~n38 ) | ( x19 & n40 ) | ( ~n38 & n40 ) ;
  assign n44 = x19 | n43 ;
  assign n45 = x15 & n44 ;
  assign n46 = ( ~x18 & n41 ) | ( ~x18 & n45 ) | ( n41 & n45 ) ;
  assign n47 = ~n41 & n46 ;
  assign n74 = n47 & n72 ;
  assign n75 = ( ~x25 & n73 ) | ( ~x25 & n74 ) | ( n73 & n74 ) ;
  assign n76 = x5 | x7 ;
  assign n77 = ( ~x4 & x6 ) | ( ~x4 & n76 ) | ( x6 & n76 ) ;
  assign n78 = x4 | n77 ;
  assign n79 = x10 | x15 ;
  assign n80 = ( x12 & n78 ) | ( x12 & n79 ) | ( n78 & n79 ) ;
  assign n81 = n78 & ~n80 ;
  assign n82 = ~x10 & x12 ;
  assign n83 = ~x2 & x15 ;
  assign n84 = ( x10 & n82 ) | ( x10 & n83 ) | ( n82 & n83 ) ;
  assign n85 = n81 | n84 ;
  assign n86 = x11 | n85 ;
  assign n87 = x11 & ~n83 ;
  assign n88 = n86 & ~n87 ;
  assign n89 = x19 & ~x22 ;
  assign n90 = ( x24 & n88 ) | ( x24 & ~n89 ) | ( n88 & ~n89 ) ;
  assign n91 = n88 & ~n90 ;
  assign n92 = ~x9 & n91 ;
  assign n93 = ( x0 & ~x18 ) | ( x0 & n92 ) | ( ~x18 & n92 ) ;
  assign n94 = ~x0 & n93 ;
  assign n95 = x25 & ~n94 ;
  assign n96 = ( x18 & n94 ) | ( x18 & ~n95 ) | ( n94 & ~n95 ) ;
  assign n120 = x18 & x25 ;
  assign n112 = ( ~x3 & x15 ) | ( ~x3 & x19 ) | ( x15 & x19 ) ;
  assign n113 = x19 & ~n112 ;
  assign n114 = ( x8 & x15 ) | ( x8 & n113 ) | ( x15 & n113 ) ;
  assign n115 = ( ~n112 & n113 ) | ( ~n112 & n114 ) | ( n113 & n114 ) ;
  assign n116 = x0 & ~n115 ;
  assign n97 = ~x6 & x7 ;
  assign n98 = x12 | x15 ;
  assign n99 = ( x6 & n97 ) | ( x6 & ~n98 ) | ( n97 & ~n98 ) ;
  assign n102 = ( ~x10 & x11 ) | ( ~x10 & n99 ) | ( x11 & n99 ) ;
  assign n100 = ~x11 & x12 ;
  assign n101 = ( x11 & n83 ) | ( x11 & n100 ) | ( n83 & n100 ) ;
  assign n103 = ~x10 & n101 ;
  assign n104 = ( ~x11 & n102 ) | ( ~x11 & n103 ) | ( n102 & n103 ) ;
  assign n109 = ( x9 & ~x24 ) | ( x9 & n104 ) | ( ~x24 & n104 ) ;
  assign n105 = x1 & x15 ;
  assign n106 = x9 & n105 ;
  assign n107 = x15 & ~n106 ;
  assign n108 = ( x2 & n106 ) | ( x2 & ~n107 ) | ( n106 & ~n107 ) ;
  assign n110 = ~x24 & n108 ;
  assign n111 = ( ~x9 & n109 ) | ( ~x9 & n110 ) | ( n109 & n110 ) ;
  assign n117 = x19 & n111 ;
  assign n118 = x0 | n117 ;
  assign n119 = ~n116 & n118 ;
  assign n121 = ~x22 & n119 ;
  assign n122 = x18 | n121 ;
  assign n123 = ~n120 & n122 ;
  assign n124 = ~x5 & x7 ;
  assign n125 = ( x5 & ~n98 ) | ( x5 & n124 ) | ( ~n98 & n124 ) ;
  assign n126 = ( x10 & ~x11 ) | ( x10 & n125 ) | ( ~x11 & n125 ) ;
  assign n127 = ~x11 & n84 ;
  assign n128 = ( ~x10 & n126 ) | ( ~x10 & n127 ) | ( n126 & n127 ) ;
  assign n129 = ( x9 & ~x24 ) | ( x9 & n128 ) | ( ~x24 & n128 ) ;
  assign n130 = ( ~x9 & n110 ) | ( ~x9 & n129 ) | ( n110 & n129 ) ;
  assign n131 = x19 & n130 ;
  assign n132 = x0 | n131 ;
  assign n133 = ~n116 & n132 ;
  assign n134 = ~x22 & n133 ;
  assign n135 = x18 | n134 ;
  assign n136 = x17 & ~x25 ;
  assign n137 = x18 & ~n136 ;
  assign n138 = n135 & ~n137 ;
  assign n139 = ~x22 & n45 ;
  assign n140 = x23 & ~n139 ;
  assign n149 = ( x11 & x12 ) | ( x11 & x15 ) | ( x12 & x15 ) ;
  assign n150 = ~x10 & n149 ;
  assign n151 = ( x10 & x15 ) | ( x10 & n150 ) | ( x15 & n150 ) ;
  assign n157 = ( x2 & ~x9 ) | ( x2 & n151 ) | ( ~x9 & n151 ) ;
  assign n152 = x12 | x23 ;
  assign n153 = ( x15 & n78 ) | ( x15 & n152 ) | ( n78 & n152 ) ;
  assign n154 = n78 & ~n153 ;
  assign n155 = ~x10 & n154 ;
  assign n156 = ~x11 & n155 ;
  assign n158 = ~x9 & n156 ;
  assign n159 = ( ~x2 & n157 ) | ( ~x2 & n158 ) | ( n157 & n158 ) ;
  assign n146 = ( x15 & x23 ) | ( x15 & ~n106 ) | ( x23 & ~n106 ) ;
  assign n147 = x2 & n146 ;
  assign n148 = ( x2 & n106 ) | ( x2 & ~n147 ) | ( n106 & ~n147 ) ;
  assign n160 = n148 & ~n159 ;
  assign n161 = x19 & ~x24 ;
  assign n162 = ( n159 & n160 ) | ( n159 & n161 ) | ( n160 & n161 ) ;
  assign n163 = x0 | n162 ;
  assign n141 = x15 & x19 ;
  assign n142 = x19 & ~n141 ;
  assign n143 = ~x23 & n142 ;
  assign n144 = ( x8 & ~n141 ) | ( x8 & n142 ) | ( ~n141 & n142 ) ;
  assign n145 = ( x15 & n143 ) | ( x15 & n144 ) | ( n143 & n144 ) ;
  assign n164 = x3 & n145 ;
  assign n165 = x0 & ~n164 ;
  assign n166 = n163 & ~n165 ;
  assign n167 = ~x22 & n166 ;
  assign n168 = ~x20 & n167 ;
  assign n169 = ( x18 & x23 ) | ( x18 & ~x25 ) | ( x23 & ~x25 ) ;
  assign n170 = ( x18 & ~x20 ) | ( x18 & x25 ) | ( ~x20 & x25 ) ;
  assign n171 = n169 & n170 ;
  assign n172 = ( ~x19 & x20 ) | ( ~x19 & n171 ) | ( x20 & n171 ) ;
  assign n173 = x23 | n171 ;
  assign n174 = ( x19 & n172 ) | ( x19 & n173 ) | ( n172 & n173 ) ;
  assign n175 = ( ~n140 & n168 ) | ( ~n140 & n174 ) | ( n168 & n174 ) ;
  assign n176 = x18 & ~n174 ;
  assign n177 = ( n140 & n175 ) | ( n140 & ~n176 ) | ( n175 & ~n176 ) ;
  assign n178 = ~x18 & n168 ;
  assign n179 = x18 & ~x20 ;
  assign n180 = ~x25 & n179 ;
  assign n181 = x24 | n34 ;
  assign n182 = x0 | n181 ;
  assign n183 = ( n38 & ~n139 ) | ( n38 & n182 ) | ( ~n139 & n182 ) ;
  assign n184 = ~x19 & n139 ;
  assign n185 = ( n38 & ~n183 ) | ( n38 & n184 ) | ( ~n183 & n184 ) ;
  assign n186 = ( x18 & ~x20 ) | ( x18 & n185 ) | ( ~x20 & n185 ) ;
  assign n187 = ( x18 & x20 ) | ( x18 & x25 ) | ( x20 & x25 ) ;
  assign n188 = n186 & ~n187 ;
  assign n189 = x23 & ~n188 ;
  assign n190 = ( x9 & ~x11 ) | ( x9 & n82 ) | ( ~x11 & n82 ) ;
  assign n191 = ~x9 & n190 ;
  assign y0 = n33 ;
  assign y1 = ~n75 ;
  assign y2 = n96 ;
  assign y3 = n123 ;
  assign y4 = n138 ;
  assign y5 = n177 ;
  assign y6 = n178 ;
  assign y7 = n180 ;
  assign y8 = n189 ;
  assign y9 = n191 ;
endmodule
