module top( in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ , out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ );
  input in_6_ , in_15_ , in_13_ , in_14_ , in_2_ , in_10_ , in_24_ , in_8_ , in_22_ , in_20_ , in_7_ , in_25_ , in_5_ , in_4_ , in_23_ , in_27_ , in_1_ , in_0_ , in_16_ , in_30_ , in_26_ , in_12_ , in_11_ , in_17_ , in_19_ , in_18_ , in_21_ , in_31_ , in_29_ , in_28_ , in_9_ , in_3_ ;
  output out_2_ , out_1_ , out_3_ , out_0_ , out_5_ , out_4_ ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ;
  assign n33 = in_29_ | in_28_ ;
  assign n34 = in_20_ | in_21_ ;
  assign n35 = in_16_ | in_17_ ;
  assign n36 = in_19_ & in_18_ ;
  assign n37 = ( n34 & n35 ) | ( n34 & n36 ) | ( n35 & n36 ) ;
  assign n38 = ( ~n34 & n35 ) | ( ~n34 & n36 ) | ( n35 & n36 ) ;
  assign n39 = ( n34 & ~n37 ) | ( n34 & n38 ) | ( ~n37 & n38 ) ;
  assign n40 = in_27_ & in_26_ ;
  assign n41 = in_22_ & in_23_ ;
  assign n42 = in_24_ | in_25_ ;
  assign n43 = ( n40 & n41 ) | ( n40 & n42 ) | ( n41 & n42 ) ;
  assign n44 = ( ~n40 & n41 ) | ( ~n40 & n42 ) | ( n41 & n42 ) ;
  assign n45 = ( n40 & ~n43 ) | ( n40 & n44 ) | ( ~n43 & n44 ) ;
  assign n46 = ( n33 & n39 ) | ( n33 & n45 ) | ( n39 & n45 ) ;
  assign n47 = ( n37 & n43 ) | ( n37 & n46 ) | ( n43 & n46 ) ;
  assign n48 = ( n37 & n43 ) | ( n37 & ~n46 ) | ( n43 & ~n46 ) ;
  assign n49 = ( n46 & ~n47 ) | ( n46 & n48 ) | ( ~n47 & n48 ) ;
  assign n50 = in_30_ & in_31_ ;
  assign n51 = ( ~n33 & n39 ) | ( ~n33 & n45 ) | ( n39 & n45 ) ;
  assign n52 = ( n33 & ~n46 ) | ( n33 & n51 ) | ( ~n46 & n51 ) ;
  assign n53 = n50 & n52 ;
  assign n54 = n49 & n53 ;
  assign n55 = n49 | n53 ;
  assign n56 = ~n54 & n55 ;
  assign n57 = in_13_ | in_12_ ;
  assign n58 = in_5_ | in_4_ ;
  assign n59 = in_1_ | in_0_ ;
  assign n60 = in_2_ & in_3_ ;
  assign n61 = ( n58 & n59 ) | ( n58 & n60 ) | ( n59 & n60 ) ;
  assign n62 = ( ~n58 & n59 ) | ( ~n58 & n60 ) | ( n59 & n60 ) ;
  assign n63 = ( n58 & ~n61 ) | ( n58 & n62 ) | ( ~n61 & n62 ) ;
  assign n64 = in_10_ & in_11_ ;
  assign n65 = in_6_ & in_7_ ;
  assign n66 = in_8_ | in_9_ ;
  assign n67 = ( n64 & n65 ) | ( n64 & n66 ) | ( n65 & n66 ) ;
  assign n68 = ( ~n64 & n65 ) | ( ~n64 & n66 ) | ( n65 & n66 ) ;
  assign n69 = ( n64 & ~n67 ) | ( n64 & n68 ) | ( ~n67 & n68 ) ;
  assign n70 = ( n57 & n63 ) | ( n57 & n69 ) | ( n63 & n69 ) ;
  assign n71 = ( n61 & n67 ) | ( n61 & n70 ) | ( n67 & n70 ) ;
  assign n72 = ( n61 & n67 ) | ( n61 & ~n70 ) | ( n67 & ~n70 ) ;
  assign n73 = ( n70 & ~n71 ) | ( n70 & n72 ) | ( ~n71 & n72 ) ;
  assign n74 = in_15_ & in_14_ ;
  assign n75 = ( ~n57 & n63 ) | ( ~n57 & n69 ) | ( n63 & n69 ) ;
  assign n76 = ( n57 & ~n70 ) | ( n57 & n75 ) | ( ~n70 & n75 ) ;
  assign n77 = n74 & n76 ;
  assign n78 = n73 & n77 ;
  assign n79 = n73 | n77 ;
  assign n80 = ~n78 & n79 ;
  assign n81 = n56 & n80 ;
  assign n82 = n56 | n80 ;
  assign n83 = ~n81 & n82 ;
  assign n84 = n50 | n52 ;
  assign n85 = ~n53 & n84 ;
  assign n86 = n74 | n76 ;
  assign n87 = ~n77 & n86 ;
  assign n88 = n85 & n87 ;
  assign n89 = n83 & n88 ;
  assign n90 = n83 | n88 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = n85 | n87 ;
  assign n93 = ~n88 & n92 ;
  assign n94 = n47 & n54 ;
  assign n95 = n47 | n54 ;
  assign n96 = ~n94 & n95 ;
  assign n97 = n71 & n78 ;
  assign n98 = n71 | n78 ;
  assign n99 = ~n97 & n98 ;
  assign n100 = n96 & n99 ;
  assign n101 = n96 | n99 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = ( n56 & n80 ) | ( n56 & n88 ) | ( n80 & n88 ) ;
  assign n104 = n102 & n103 ;
  assign n105 = n102 | n103 ;
  assign n106 = ~n104 & n105 ;
  assign n107 = ( n96 & n99 ) | ( n96 & n103 ) | ( n99 & n103 ) ;
  assign n108 = ( n94 & n97 ) | ( n94 & n107 ) | ( n97 & n107 ) ;
  assign n109 = n94 | n97 ;
  assign n110 = n94 & n97 ;
  assign n111 = n109 & ~n110 ;
  assign n112 = n107 & n111 ;
  assign n113 = n107 | n111 ;
  assign n114 = ~n112 & n113 ;
  assign out_2_ = n91 ;
  assign out_1_ = n93 ;
  assign out_3_ = n106 ;
  assign out_0_ = 1'b0 ;
  assign out_5_ = n108 ;
  assign out_4_ = n114 ;
endmodule
