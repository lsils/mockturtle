module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , y0 , y1 , y2 , y3 , y4 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 ;
  output y0 , y1 , y2 , y3 , y4 ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 ;
  assign n17 = ( x4 & ~x6 ) | ( x4 & x12 ) | ( ~x6 & x12 ) ;
  assign n18 = ( ~x5 & x6 ) | ( ~x5 & x12 ) | ( x6 & x12 ) ;
  assign n19 = ~n17 & n18 ;
  assign n20 = ( x4 & ~x7 ) | ( x4 & x12 ) | ( ~x7 & x12 ) ;
  assign n21 = ( x5 & x7 ) | ( x5 & ~x12 ) | ( x7 & ~x12 ) ;
  assign n22 = n20 & n21 ;
  assign n23 = n19 | n22 ;
  assign n24 = x8 & ~n23 ;
  assign n25 = ~x7 & x12 ;
  assign n26 = ( x5 & x7 ) | ( x5 & x12 ) | ( x7 & x12 ) ;
  assign n27 = ~x6 & x12 ;
  assign n28 = ( x5 & x12 ) | ( x5 & n27 ) | ( x12 & n27 ) ;
  assign n29 = ( n25 & n26 ) | ( n25 & ~n28 ) | ( n26 & ~n28 ) ;
  assign n30 = x4 & n29 ;
  assign n31 = x8 | n30 ;
  assign n32 = ~n24 & n31 ;
  assign n33 = x4 & x5 ;
  assign n34 = x5 & ~n33 ;
  assign n35 = x12 & n34 ;
  assign n36 = ( x0 & ~n33 ) | ( x0 & n34 ) | ( ~n33 & n34 ) ;
  assign n37 = ( x4 & n35 ) | ( x4 & n36 ) | ( n35 & n36 ) ;
  assign n38 = n32 | n37 ;
  assign n39 = ( ~x6 & n32 ) | ( ~x6 & n38 ) | ( n32 & n38 ) ;
  assign n40 = x6 & ~x9 ;
  assign n41 = ( x5 & ~x13 ) | ( x5 & n40 ) | ( ~x13 & n40 ) ;
  assign n42 = ( x5 & x6 ) | ( x5 & ~n40 ) | ( x6 & ~n40 ) ;
  assign n43 = ~n41 & n42 ;
  assign n44 = ~x4 & n43 ;
  assign n45 = ~x9 & x13 ;
  assign n46 = ( x6 & ~x9 ) | ( x6 & x13 ) | ( ~x9 & x13 ) ;
  assign n47 = x1 | x6 ;
  assign n48 = ( n45 & ~n46 ) | ( n45 & n47 ) | ( ~n46 & n47 ) ;
  assign n49 = ~x5 & n48 ;
  assign n50 = x0 & x7 ;
  assign n51 = x12 | n50 ;
  assign n52 = ( x8 & n50 ) | ( x8 & n51 ) | ( n50 & n51 ) ;
  assign n53 = ( x9 & ~x13 ) | ( x9 & n52 ) | ( ~x13 & n52 ) ;
  assign n54 = ( x9 & x13 ) | ( x9 & n52 ) | ( x13 & n52 ) ;
  assign n55 = ( x13 & n53 ) | ( x13 & ~n54 ) | ( n53 & ~n54 ) ;
  assign n56 = x5 & n55 ;
  assign n57 = n49 | n56 ;
  assign n58 = x4 & n57 ;
  assign n59 = n44 | n58 ;
  assign n60 = x6 & ~x10 ;
  assign n61 = ( x5 & ~x14 ) | ( x5 & n60 ) | ( ~x14 & n60 ) ;
  assign n62 = ( x5 & x6 ) | ( x5 & ~n60 ) | ( x6 & ~n60 ) ;
  assign n63 = ~n61 & n62 ;
  assign n64 = ~x4 & n63 ;
  assign n65 = ~x10 & x14 ;
  assign n66 = ( x6 & ~x10 ) | ( x6 & x14 ) | ( ~x10 & x14 ) ;
  assign n67 = x2 | x6 ;
  assign n68 = ( n65 & ~n66 ) | ( n65 & n67 ) | ( ~n66 & n67 ) ;
  assign n69 = ~x5 & n68 ;
  assign n70 = x1 & n52 ;
  assign n71 = x13 | n70 ;
  assign n72 = ( x9 & n70 ) | ( x9 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ( x10 & ~x14 ) | ( x10 & n72 ) | ( ~x14 & n72 ) ;
  assign n74 = ( x10 & x14 ) | ( x10 & n72 ) | ( x14 & n72 ) ;
  assign n75 = ( x14 & n73 ) | ( x14 & ~n74 ) | ( n73 & ~n74 ) ;
  assign n76 = x5 & n75 ;
  assign n77 = n69 | n76 ;
  assign n78 = x4 & n77 ;
  assign n79 = n64 | n78 ;
  assign n80 = x2 & n72 ;
  assign n81 = x14 | n80 ;
  assign n82 = ( x10 & n80 ) | ( x10 & n81 ) | ( n80 & n81 ) ;
  assign n83 = ( x11 & ~x15 ) | ( x11 & n82 ) | ( ~x15 & n82 ) ;
  assign n84 = ( x11 & n82 ) | ( x11 & ~n83 ) | ( n82 & ~n83 ) ;
  assign n85 = ( x15 & n83 ) | ( x15 & ~n84 ) | ( n83 & ~n84 ) ;
  assign n86 = x5 & n85 ;
  assign n87 = ~x11 & x15 ;
  assign n88 = ( x6 & ~x11 ) | ( x6 & x15 ) | ( ~x11 & x15 ) ;
  assign n89 = x3 | x6 ;
  assign n90 = ( n87 & ~n88 ) | ( n87 & n89 ) | ( ~n88 & n89 ) ;
  assign n91 = x5 | n90 ;
  assign n92 = ( ~x5 & n86 ) | ( ~x5 & n91 ) | ( n86 & n91 ) ;
  assign n93 = x4 & n92 ;
  assign n94 = x6 & ~x11 ;
  assign n95 = ( x5 & ~x15 ) | ( x5 & n94 ) | ( ~x15 & n94 ) ;
  assign n96 = ( x5 & x6 ) | ( x5 & ~n94 ) | ( x6 & ~n94 ) ;
  assign n97 = ~n95 & n96 ;
  assign n98 = x4 | n97 ;
  assign n99 = ( ~x4 & n93 ) | ( ~x4 & n98 ) | ( n93 & n98 ) ;
  assign n100 = ( ~x0 & x2 ) | ( ~x0 & x7 ) | ( x2 & x7 ) ;
  assign n101 = x1 & x12 ;
  assign n102 = x8 & n101 ;
  assign n103 = x13 | n102 ;
  assign n104 = ( x9 & n102 ) | ( x9 & n103 ) | ( n102 & n103 ) ;
  assign n105 = x2 & n104 ;
  assign n106 = ( x0 & n100 ) | ( x0 & n105 ) | ( n100 & n105 ) ;
  assign n107 = x14 | n106 ;
  assign n108 = ( x10 & n106 ) | ( x10 & n107 ) | ( n106 & n107 ) ;
  assign n109 = x3 & n108 ;
  assign n110 = x15 | n109 ;
  assign n111 = ( x11 & n109 ) | ( x11 & n110 ) | ( n109 & n110 ) ;
  assign y0 = n39 ;
  assign y1 = n59 ;
  assign y2 = n79 ;
  assign y3 = n99 ;
  assign y4 = n111 ;
endmodule
