module top( a_11_ , a_18_ , a_15_ , a_3_ , a_9_ , a_6_ , a_28_ , a_7_ , a_25_ , a_29_ , a_22_ , a_26_ , a_1_ , a_8_ , a_16_ , a_10_ , a_30_ , a_12_ , a_24_ , a_5_ , a_0_ , a_17_ , a_4_ , a_14_ , a_20_ , a_27_ , a_23_ , a_13_ , a_31_ , a_2_ , a_19_ , a_21_ , b_9_ , b_1_ , b_17_ , b_11_ , b_31_ , b_26_ , b_29_ , b_24_ , b_23_ , b_8_ , b_4_ , b_25_ , b_7_ , b_5_ , b_18_ , b_12_ , b_16_ , b_22_ , b_14_ , b_20_ , b_15_ , b_3_ , b_30_ , b_27_ , b_21_ , b_19_ , b_13_ , b_6_ , b_0_ , b_10_ , b_28_ , b_2_ );
  input a_11_ , a_18_ , a_15_ , a_3_ , a_9_ , a_6_ , a_28_ , a_7_ , a_25_ , a_29_ , a_22_ , a_26_ , a_1_ , a_8_ , a_16_ , a_10_ , a_30_ , a_12_ , a_24_ , a_5_ , a_0_ , a_17_ , a_4_ , a_14_ , a_20_ , a_27_ , a_23_ , a_13_ , a_31_ , a_2_ , a_19_ , a_21_ ;
  output b_9_ , b_1_ , b_17_ , b_11_ , b_31_ , b_26_ , b_29_ , b_24_ , b_23_ , b_8_ , b_4_ , b_25_ , b_7_ , b_5_ , b_18_ , b_12_ , b_16_ , b_22_ , b_14_ , b_20_ , b_15_ , b_3_ , b_30_ , b_27_ , b_21_ , b_19_ , b_13_ , b_6_ , b_0_ , b_10_ , b_28_ , b_2_ ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 ;
  assign n33 = a_15_ | a_14_ ;
  assign n34 = a_12_ & a_13_ ;
  assign n35 = n33 & n34 ;
  assign n36 = a_15_ & a_14_ ;
  assign n37 = a_12_ | a_13_ ;
  assign n38 = n36 & n37 ;
  assign n39 = n35 | n38 ;
  assign n40 = a_11_ | a_10_ ;
  assign n41 = a_9_ & a_8_ ;
  assign n42 = n40 | n41 ;
  assign n43 = a_11_ & a_10_ ;
  assign n44 = a_9_ | a_8_ ;
  assign n45 = n43 | n44 ;
  assign n46 = n42 & n45 ;
  assign n47 = n39 & n46 ;
  assign n48 = n33 | n34 ;
  assign n49 = n36 | n37 ;
  assign n50 = n48 | n49 ;
  assign n51 = n40 & n41 ;
  assign n52 = n43 & n44 ;
  assign n53 = n51 & n52 ;
  assign n54 = n50 & n53 ;
  assign n55 = n47 & n54 ;
  assign n56 = n35 & n38 ;
  assign n57 = n42 | n45 ;
  assign n58 = n56 & n57 ;
  assign n59 = n48 & n49 ;
  assign n60 = n51 | n52 ;
  assign n61 = n59 & n60 ;
  assign n62 = n58 & n61 ;
  assign n63 = n55 | n62 ;
  assign n64 = a_3_ | a_2_ ;
  assign n65 = a_1_ & a_0_ ;
  assign n66 = n64 | n65 ;
  assign n67 = a_3_ & a_2_ ;
  assign n68 = a_1_ | a_0_ ;
  assign n69 = n67 | n68 ;
  assign n70 = n66 | n69 ;
  assign n71 = a_6_ | a_7_ ;
  assign n72 = a_5_ & a_4_ ;
  assign n73 = n71 & n72 ;
  assign n74 = a_6_ & a_7_ ;
  assign n75 = a_5_ | a_4_ ;
  assign n76 = n74 & n75 ;
  assign n77 = n73 & n76 ;
  assign n78 = n70 | n77 ;
  assign n79 = n64 & n65 ;
  assign n80 = n67 & n68 ;
  assign n81 = n79 | n80 ;
  assign n82 = n71 | n72 ;
  assign n83 = n74 | n75 ;
  assign n84 = n82 & n83 ;
  assign n85 = n81 | n84 ;
  assign n86 = n78 | n85 ;
  assign n87 = n79 & n80 ;
  assign n88 = n82 | n83 ;
  assign n89 = n87 | n88 ;
  assign n90 = n66 & n69 ;
  assign n91 = n73 | n76 ;
  assign n92 = n90 | n91 ;
  assign n93 = n89 | n92 ;
  assign n94 = n86 & n93 ;
  assign n95 = n63 | n94 ;
  assign n96 = n39 | n46 ;
  assign n97 = n50 | n53 ;
  assign n98 = n96 & n97 ;
  assign n99 = n56 | n57 ;
  assign n100 = n59 | n60 ;
  assign n101 = n99 & n100 ;
  assign n102 = n98 | n101 ;
  assign n103 = n70 & n77 ;
  assign n104 = n81 & n84 ;
  assign n105 = n103 | n104 ;
  assign n106 = n87 & n88 ;
  assign n107 = n90 & n91 ;
  assign n108 = n106 | n107 ;
  assign n109 = n105 & n108 ;
  assign n110 = n102 | n109 ;
  assign n111 = n95 | n110 ;
  assign n112 = n47 | n54 ;
  assign n113 = n58 | n61 ;
  assign n114 = n112 | n113 ;
  assign n115 = n78 & n85 ;
  assign n116 = n89 & n92 ;
  assign n117 = n115 & n116 ;
  assign n118 = n114 | n117 ;
  assign n119 = n96 | n97 ;
  assign n120 = n99 | n100 ;
  assign n121 = n119 | n120 ;
  assign n122 = n103 & n104 ;
  assign n123 = n106 & n107 ;
  assign n124 = n122 & n123 ;
  assign n125 = n121 | n124 ;
  assign n126 = n118 | n125 ;
  assign n127 = n111 & n126 ;
  assign n128 = n55 & n62 ;
  assign n129 = n86 | n93 ;
  assign n130 = n128 | n129 ;
  assign n131 = n98 & n101 ;
  assign n132 = n105 | n108 ;
  assign n133 = n131 | n132 ;
  assign n134 = n130 | n133 ;
  assign n135 = n119 & n120 ;
  assign n136 = n122 | n123 ;
  assign n137 = n135 | n136 ;
  assign n138 = n112 & n113 ;
  assign n139 = n115 | n116 ;
  assign n140 = n138 | n139 ;
  assign n141 = n137 | n140 ;
  assign n142 = n134 & n141 ;
  assign n143 = n127 & n142 ;
  assign n144 = a_26_ | a_27_ ;
  assign n145 = a_25_ & a_24_ ;
  assign n146 = n144 & n145 ;
  assign n147 = a_26_ & a_27_ ;
  assign n148 = a_25_ | a_24_ ;
  assign n149 = n147 & n148 ;
  assign n150 = n146 & n149 ;
  assign n151 = a_30_ & a_31_ ;
  assign n152 = a_28_ | a_29_ ;
  assign n153 = n151 | n152 ;
  assign n154 = a_28_ & a_29_ ;
  assign n155 = a_30_ | a_31_ ;
  assign n156 = n154 | n155 ;
  assign n157 = n153 | n156 ;
  assign n158 = n150 & n157 ;
  assign n159 = n144 | n145 ;
  assign n160 = n147 | n148 ;
  assign n161 = n159 & n160 ;
  assign n162 = n151 & n152 ;
  assign n163 = n154 & n155 ;
  assign n164 = n162 | n163 ;
  assign n165 = n161 & n164 ;
  assign n166 = n158 & n165 ;
  assign n167 = n146 | n149 ;
  assign n168 = n153 & n156 ;
  assign n169 = n167 & n168 ;
  assign n170 = n159 | n160 ;
  assign n171 = n162 & n163 ;
  assign n172 = n170 & n171 ;
  assign n173 = n169 & n172 ;
  assign n174 = n166 & n173 ;
  assign n175 = a_22_ | a_23_ ;
  assign n176 = a_20_ & a_21_ ;
  assign n177 = n175 & n176 ;
  assign n178 = a_22_ & a_23_ ;
  assign n179 = a_20_ | a_21_ ;
  assign n180 = n178 & n179 ;
  assign n181 = n177 | n180 ;
  assign n182 = a_18_ | a_19_ ;
  assign n183 = a_16_ & a_17_ ;
  assign n184 = n182 | n183 ;
  assign n185 = a_18_ & a_19_ ;
  assign n186 = a_16_ | a_17_ ;
  assign n187 = n185 | n186 ;
  assign n188 = n184 & n187 ;
  assign n189 = n181 | n188 ;
  assign n190 = n175 | n176 ;
  assign n191 = n178 | n179 ;
  assign n192 = n190 | n191 ;
  assign n193 = n182 & n183 ;
  assign n194 = n185 & n186 ;
  assign n195 = n193 & n194 ;
  assign n196 = n192 | n195 ;
  assign n197 = n189 | n196 ;
  assign n198 = n177 & n180 ;
  assign n199 = n184 | n187 ;
  assign n200 = n198 | n199 ;
  assign n201 = n190 & n191 ;
  assign n202 = n193 | n194 ;
  assign n203 = n201 | n202 ;
  assign n204 = n200 | n203 ;
  assign n205 = n197 | n204 ;
  assign n206 = n174 & n205 ;
  assign n207 = n181 & n188 ;
  assign n208 = n192 & n195 ;
  assign n209 = n207 | n208 ;
  assign n210 = n198 & n199 ;
  assign n211 = n201 & n202 ;
  assign n212 = n210 | n211 ;
  assign n213 = n209 | n212 ;
  assign n214 = n150 | n157 ;
  assign n215 = n161 | n164 ;
  assign n216 = n214 & n215 ;
  assign n217 = n167 | n168 ;
  assign n218 = n170 | n171 ;
  assign n219 = n217 & n218 ;
  assign n220 = n216 & n219 ;
  assign n221 = n213 & n220 ;
  assign n222 = n206 & n221 ;
  assign n223 = n158 | n165 ;
  assign n224 = n169 | n172 ;
  assign n225 = n223 & n224 ;
  assign n226 = n189 & n196 ;
  assign n227 = n200 & n203 ;
  assign n228 = n226 | n227 ;
  assign n229 = n225 & n228 ;
  assign n230 = n207 & n208 ;
  assign n231 = n210 & n211 ;
  assign n232 = n230 | n231 ;
  assign n233 = n214 | n215 ;
  assign n234 = n217 | n218 ;
  assign n235 = n233 & n234 ;
  assign n236 = n232 & n235 ;
  assign n237 = n229 & n236 ;
  assign n238 = n222 | n237 ;
  assign n239 = n166 | n173 ;
  assign n240 = n197 & n204 ;
  assign n241 = n239 & n240 ;
  assign n242 = n209 & n212 ;
  assign n243 = n216 | n219 ;
  assign n244 = n242 & n243 ;
  assign n245 = n241 & n244 ;
  assign n246 = n223 | n224 ;
  assign n247 = n226 & n227 ;
  assign n248 = n246 & n247 ;
  assign n249 = n230 & n231 ;
  assign n250 = n233 | n234 ;
  assign n251 = n249 & n250 ;
  assign n252 = n248 & n251 ;
  assign n253 = n245 | n252 ;
  assign n254 = n238 | n253 ;
  assign n255 = n143 & n254 ;
  assign n256 = n63 & n94 ;
  assign n257 = n102 & n109 ;
  assign n258 = n256 | n257 ;
  assign n259 = n114 & n117 ;
  assign n260 = n121 & n124 ;
  assign n261 = n259 | n260 ;
  assign n262 = n258 & n261 ;
  assign n263 = n128 & n129 ;
  assign n264 = n131 & n132 ;
  assign n265 = n263 | n264 ;
  assign n266 = n138 & n139 ;
  assign n267 = n135 & n136 ;
  assign n268 = n266 | n267 ;
  assign n269 = n265 & n268 ;
  assign n270 = n262 & n269 ;
  assign n271 = n239 | n240 ;
  assign n272 = n242 | n243 ;
  assign n273 = n271 & n272 ;
  assign n274 = n246 | n247 ;
  assign n275 = n249 | n250 ;
  assign n276 = n274 & n275 ;
  assign n277 = n273 | n276 ;
  assign n278 = n174 | n205 ;
  assign n279 = n213 | n220 ;
  assign n280 = n278 & n279 ;
  assign n281 = n225 | n228 ;
  assign n282 = n232 | n235 ;
  assign n283 = n281 & n282 ;
  assign n284 = n280 | n283 ;
  assign n285 = n277 | n284 ;
  assign n286 = n270 & n285 ;
  assign n287 = n255 | n286 ;
  assign n288 = n95 & n110 ;
  assign n289 = n118 & n125 ;
  assign n290 = n288 & n289 ;
  assign n291 = n130 & n133 ;
  assign n292 = n137 & n140 ;
  assign n293 = n291 & n292 ;
  assign n294 = n290 & n293 ;
  assign n295 = n206 | n221 ;
  assign n296 = n229 | n236 ;
  assign n297 = n295 | n296 ;
  assign n298 = n241 | n244 ;
  assign n299 = n248 | n251 ;
  assign n300 = n298 | n299 ;
  assign n301 = n297 | n300 ;
  assign n302 = n294 & n301 ;
  assign n303 = n256 & n257 ;
  assign n304 = n259 & n260 ;
  assign n305 = n303 & n304 ;
  assign n306 = n263 & n264 ;
  assign n307 = n266 & n267 ;
  assign n308 = n306 & n307 ;
  assign n309 = n305 & n308 ;
  assign n310 = n271 | n272 ;
  assign n311 = n274 | n275 ;
  assign n312 = n310 | n311 ;
  assign n313 = n278 | n279 ;
  assign n314 = n281 | n282 ;
  assign n315 = n313 | n314 ;
  assign n316 = n312 | n315 ;
  assign n317 = n309 & n316 ;
  assign n318 = n302 | n317 ;
  assign n319 = n287 & n318 ;
  assign n320 = n111 | n126 ;
  assign n321 = n134 | n141 ;
  assign n322 = n320 & n321 ;
  assign n323 = n222 & n237 ;
  assign n324 = n245 & n252 ;
  assign n325 = n323 | n324 ;
  assign n326 = n322 & n325 ;
  assign n327 = n258 | n261 ;
  assign n328 = n265 | n268 ;
  assign n329 = n327 & n328 ;
  assign n330 = n273 & n276 ;
  assign n331 = n280 & n283 ;
  assign n332 = n330 | n331 ;
  assign n333 = n329 & n332 ;
  assign n334 = n326 | n333 ;
  assign n335 = n288 | n289 ;
  assign n336 = n291 | n292 ;
  assign n337 = n335 & n336 ;
  assign n338 = n295 & n296 ;
  assign n339 = n298 & n299 ;
  assign n340 = n338 | n339 ;
  assign n341 = n337 & n340 ;
  assign n342 = n303 | n304 ;
  assign n343 = n306 | n307 ;
  assign n344 = n342 & n343 ;
  assign n345 = n310 & n311 ;
  assign n346 = n313 & n314 ;
  assign n347 = n345 | n346 ;
  assign n348 = n344 & n347 ;
  assign n349 = n341 | n348 ;
  assign n350 = n334 & n349 ;
  assign n351 = n319 & n350 ;
  assign n352 = n127 | n142 ;
  assign n353 = n238 & n253 ;
  assign n354 = n352 & n353 ;
  assign n355 = n262 | n269 ;
  assign n356 = n277 & n284 ;
  assign n357 = n355 & n356 ;
  assign n358 = n354 | n357 ;
  assign n359 = n290 | n293 ;
  assign n360 = n297 & n300 ;
  assign n361 = n359 & n360 ;
  assign n362 = n305 | n308 ;
  assign n363 = n312 & n315 ;
  assign n364 = n362 & n363 ;
  assign n365 = n361 | n364 ;
  assign n366 = n358 & n365 ;
  assign n367 = n320 | n321 ;
  assign n368 = n323 & n324 ;
  assign n369 = n367 & n368 ;
  assign n370 = n327 | n328 ;
  assign n371 = n330 & n331 ;
  assign n372 = n370 & n371 ;
  assign n373 = n369 | n372 ;
  assign n374 = n335 | n336 ;
  assign n375 = n338 & n339 ;
  assign n376 = n374 & n375 ;
  assign n377 = n342 | n343 ;
  assign n378 = n345 & n346 ;
  assign n379 = n377 & n378 ;
  assign n380 = n376 | n379 ;
  assign n381 = n373 & n380 ;
  assign n382 = n366 & n381 ;
  assign n383 = n351 | n382 ;
  assign n384 = n255 & n286 ;
  assign n385 = n302 & n317 ;
  assign n386 = n384 & n385 ;
  assign n387 = n326 & n333 ;
  assign n388 = n341 & n348 ;
  assign n389 = n387 & n388 ;
  assign n390 = n386 & n389 ;
  assign n391 = n354 & n357 ;
  assign n392 = n361 & n364 ;
  assign n393 = n391 & n392 ;
  assign n394 = n369 & n372 ;
  assign n395 = n376 & n379 ;
  assign n396 = n394 & n395 ;
  assign n397 = n393 & n396 ;
  assign n398 = n390 | n397 ;
  assign n399 = n143 | n254 ;
  assign n400 = n270 | n285 ;
  assign n401 = n399 & n400 ;
  assign n402 = n294 | n301 ;
  assign n403 = n309 | n316 ;
  assign n404 = n402 & n403 ;
  assign n405 = n401 & n404 ;
  assign n406 = n322 | n325 ;
  assign n407 = n329 | n332 ;
  assign n408 = n406 & n407 ;
  assign n409 = n337 | n340 ;
  assign n410 = n344 | n347 ;
  assign n411 = n409 & n410 ;
  assign n412 = n408 & n411 ;
  assign n413 = n405 & n412 ;
  assign n414 = n352 | n353 ;
  assign n415 = n355 | n356 ;
  assign n416 = n414 & n415 ;
  assign n417 = n359 | n360 ;
  assign n418 = n362 | n363 ;
  assign n419 = n417 & n418 ;
  assign n420 = n416 & n419 ;
  assign n421 = n367 | n368 ;
  assign n422 = n370 | n371 ;
  assign n423 = n421 & n422 ;
  assign n424 = n374 | n375 ;
  assign n425 = n377 | n378 ;
  assign n426 = n424 & n425 ;
  assign n427 = n423 & n426 ;
  assign n428 = n420 & n427 ;
  assign n429 = n413 | n428 ;
  assign n430 = n319 | n350 ;
  assign n431 = n366 | n381 ;
  assign n432 = n430 | n431 ;
  assign n433 = n399 | n400 ;
  assign n434 = n402 | n403 ;
  assign n435 = n433 | n434 ;
  assign n436 = n406 | n407 ;
  assign n437 = n409 | n410 ;
  assign n438 = n436 | n437 ;
  assign n439 = n435 | n438 ;
  assign n440 = n414 | n415 ;
  assign n441 = n417 | n418 ;
  assign n442 = n440 | n441 ;
  assign n443 = n421 | n422 ;
  assign n444 = n424 | n425 ;
  assign n445 = n443 | n444 ;
  assign n446 = n442 | n445 ;
  assign n447 = n439 | n446 ;
  assign n448 = n433 & n434 ;
  assign n449 = n436 & n437 ;
  assign n450 = n448 | n449 ;
  assign n451 = n440 & n441 ;
  assign n452 = n443 & n444 ;
  assign n453 = n451 | n452 ;
  assign n454 = n450 & n453 ;
  assign n455 = n435 & n438 ;
  assign n456 = n442 & n445 ;
  assign n457 = n455 | n456 ;
  assign n458 = n448 & n449 ;
  assign n459 = n451 & n452 ;
  assign n460 = n458 & n459 ;
  assign n461 = n401 | n404 ;
  assign n462 = n408 | n411 ;
  assign n463 = n461 | n462 ;
  assign n464 = n416 | n419 ;
  assign n465 = n423 | n426 ;
  assign n466 = n464 | n465 ;
  assign n467 = n463 | n466 ;
  assign n468 = n351 & n382 ;
  assign n469 = n384 | n385 ;
  assign n470 = n387 | n388 ;
  assign n471 = n469 & n470 ;
  assign n472 = n391 | n392 ;
  assign n473 = n394 | n395 ;
  assign n474 = n472 & n473 ;
  assign n475 = n471 & n474 ;
  assign n476 = n458 | n459 ;
  assign n477 = n469 | n470 ;
  assign n478 = n472 | n473 ;
  assign n479 = n477 | n478 ;
  assign n480 = n471 | n474 ;
  assign n481 = n405 | n412 ;
  assign n482 = n420 | n427 ;
  assign n483 = n481 & n482 ;
  assign n484 = n287 | n318 ;
  assign n485 = n334 | n349 ;
  assign n486 = n484 & n485 ;
  assign n487 = n358 | n365 ;
  assign n488 = n373 | n380 ;
  assign n489 = n487 & n488 ;
  assign n490 = n486 & n489 ;
  assign n491 = n413 & n428 ;
  assign n492 = n463 & n466 ;
  assign n493 = n484 | n485 ;
  assign n494 = n487 | n488 ;
  assign n495 = n493 & n494 ;
  assign n496 = n461 & n462 ;
  assign n497 = n464 & n465 ;
  assign n498 = n496 & n497 ;
  assign n499 = n493 | n494 ;
  assign n500 = n386 | n389 ;
  assign n501 = n393 | n396 ;
  assign n502 = n500 | n501 ;
  assign n503 = n439 & n446 ;
  assign n504 = n450 | n453 ;
  assign n505 = n496 | n497 ;
  assign n506 = n481 | n482 ;
  assign n507 = n486 | n489 ;
  assign n508 = n477 & n478 ;
  assign n509 = n390 & n397 ;
  assign n510 = n430 & n431 ;
  assign n511 = n455 & n456 ;
  assign n512 = n500 & n501 ;
  assign b_9_ = n383 ;
  assign b_1_ = n398 ;
  assign b_17_ = n429 ;
  assign b_11_ = n432 ;
  assign b_31_ = n447 ;
  assign b_26_ = n454 ;
  assign b_29_ = n457 ;
  assign b_24_ = n460 ;
  assign b_23_ = n467 ;
  assign b_8_ = n468 ;
  assign b_4_ = n475 ;
  assign b_25_ = n476 ;
  assign b_7_ = n479 ;
  assign b_5_ = n480 ;
  assign b_18_ = n483 ;
  assign b_12_ = n490 ;
  assign b_16_ = n491 ;
  assign b_22_ = n492 ;
  assign b_14_ = n495 ;
  assign b_20_ = n498 ;
  assign b_15_ = n499 ;
  assign b_3_ = n502 ;
  assign b_30_ = n503 ;
  assign b_27_ = n504 ;
  assign b_21_ = n505 ;
  assign b_19_ = n506 ;
  assign b_13_ = n507 ;
  assign b_6_ = n508 ;
  assign b_0_ = n509 ;
  assign b_10_ = n510 ;
  assign b_28_ = n511 ;
  assign b_2_ = n512 ;
endmodule
