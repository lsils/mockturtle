module top( N1 , N103 , N120 , N137 , N154 , N171 , N18 , N188 , N205 , N222 , N239 , N256 , N273 , N290 , N307 , N324 , N341 , N35 , N358 , N375 , N392 , N409 , N426 , N443 , N460 , N477 , N494 , N511 , N52 , N528 , N69 , N86 , N1581 , N1901 , N2223 , N2548 , N2877 , N3211 , N3552 , N3895 , N4241 , N4591 , N4946 , N5308 , N545 , N5672 , N5971 , N6123 , N6150 , N6160 , N6170 , N6180 , N6190 , N6200 , N6210 , N6220 , N6230 , N6240 , N6250 , N6260 , N6270 , N6280 , N6287 , N6288 );
  input N1 , N103 , N120 , N137 , N154 , N171 , N18 , N188 , N205 , N222 , N239 , N256 , N273 , N290 , N307 , N324 , N341 , N35 , N358 , N375 , N392 , N409 , N426 , N443 , N460 , N477 , N494 , N511 , N52 , N528 , N69 , N86 ;
  output N1581 , N1901 , N2223 , N2548 , N2877 , N3211 , N3552 , N3895 , N4241 , N4591 , N4946 , N5308 , N545 , N5672 , N5971 , N6123 , N6150 , N6160 , N6170 , N6180 , N6190 , N6200 , N6210 , N6220 , N6230 , N6240 , N6250 , N6260 , N6270 , N6280 , N6287 , N6288 ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 ;
  assign n33 = N18 & N290 ;
  assign n34 = N1 & N273 ;
  assign n35 = n33 & n34 ;
  assign n36 = N18 & N273 ;
  assign n37 = N1 & N290 ;
  assign n38 = n36 | n37 ;
  assign n39 = ~n35 & n38 ;
  assign n40 = N1 & N307 ;
  assign n41 = N290 & N35 ;
  assign n42 = n36 & n41 ;
  assign n43 = N273 & N35 ;
  assign n44 = n33 | n43 ;
  assign n45 = ~n42 & n44 ;
  assign n46 = n35 | n45 ;
  assign n47 = n35 & n45 ;
  assign n48 = n46 & ~n47 ;
  assign n49 = ~n40 & n48 ;
  assign n50 = n40 & ~n48 ;
  assign n51 = n49 | n50 ;
  assign n52 = N1 & N324 ;
  assign n53 = n46 & ~n49 ;
  assign n54 = N18 & N307 ;
  assign n55 = N290 & N52 ;
  assign n56 = n43 & n55 ;
  assign n57 = N273 & N52 ;
  assign n58 = n41 | n57 ;
  assign n59 = ~n56 & n58 ;
  assign n60 = n42 | n59 ;
  assign n61 = n42 & n59 ;
  assign n62 = n60 & ~n61 ;
  assign n63 = ~n54 & n62 ;
  assign n64 = n54 & ~n62 ;
  assign n65 = n63 | n64 ;
  assign n66 = n53 | n65 ;
  assign n67 = n53 & n65 ;
  assign n68 = n66 & ~n67 ;
  assign n69 = ~n52 & n68 ;
  assign n70 = n52 & ~n68 ;
  assign n71 = n69 | n70 ;
  assign n72 = N1 & N341 ;
  assign n73 = n66 & ~n69 ;
  assign n74 = N18 & N324 ;
  assign n75 = n60 & ~n63 ;
  assign n76 = N307 & N35 ;
  assign n77 = N290 & N69 ;
  assign n78 = n57 & n77 ;
  assign n79 = N273 & N69 ;
  assign n80 = n55 | n79 ;
  assign n81 = ~n78 & n80 ;
  assign n82 = n56 | n81 ;
  assign n83 = n56 & n81 ;
  assign n84 = n82 & ~n83 ;
  assign n85 = ~n76 & n84 ;
  assign n86 = n76 & ~n84 ;
  assign n87 = n85 | n86 ;
  assign n88 = n75 | n87 ;
  assign n89 = n75 & n87 ;
  assign n90 = n88 & ~n89 ;
  assign n91 = ~n74 & n90 ;
  assign n92 = n74 & ~n90 ;
  assign n93 = n91 | n92 ;
  assign n94 = n73 | n93 ;
  assign n95 = n73 & n93 ;
  assign n96 = n94 & ~n95 ;
  assign n97 = ~n72 & n96 ;
  assign n98 = n72 & ~n96 ;
  assign n99 = n97 | n98 ;
  assign n100 = N1 & N358 ;
  assign n101 = n94 & ~n97 ;
  assign n102 = N18 & N341 ;
  assign n103 = n88 & ~n91 ;
  assign n104 = N324 & N35 ;
  assign n105 = n82 & ~n85 ;
  assign n106 = N307 & N52 ;
  assign n107 = N290 & N86 ;
  assign n108 = n79 & n107 ;
  assign n109 = N273 & N86 ;
  assign n110 = n77 | n109 ;
  assign n111 = ~n108 & n110 ;
  assign n112 = n78 | n111 ;
  assign n113 = n78 & n111 ;
  assign n114 = n112 & ~n113 ;
  assign n115 = ~n106 & n114 ;
  assign n116 = n106 & ~n114 ;
  assign n117 = n115 | n116 ;
  assign n118 = n105 | n117 ;
  assign n119 = n105 & n117 ;
  assign n120 = n118 & ~n119 ;
  assign n121 = ~n104 & n120 ;
  assign n122 = n104 & ~n120 ;
  assign n123 = n121 | n122 ;
  assign n124 = n103 | n123 ;
  assign n125 = n103 & n123 ;
  assign n126 = n124 & ~n125 ;
  assign n127 = ~n102 & n126 ;
  assign n128 = n102 & ~n126 ;
  assign n129 = n127 | n128 ;
  assign n130 = n101 | n129 ;
  assign n131 = n101 & n129 ;
  assign n132 = n130 & ~n131 ;
  assign n133 = ~n100 & n132 ;
  assign n134 = n100 & ~n132 ;
  assign n135 = n133 | n134 ;
  assign n136 = N1 & N375 ;
  assign n137 = n130 & ~n133 ;
  assign n138 = N18 & N358 ;
  assign n139 = n124 & ~n127 ;
  assign n140 = N341 & N35 ;
  assign n141 = n118 & ~n121 ;
  assign n142 = N324 & N52 ;
  assign n143 = n112 & ~n115 ;
  assign n144 = N307 & N69 ;
  assign n145 = N103 & N290 ;
  assign n146 = n109 & n145 ;
  assign n147 = N103 & N273 ;
  assign n148 = n107 | n147 ;
  assign n149 = ~n146 & n148 ;
  assign n150 = n108 | n149 ;
  assign n151 = n108 & n149 ;
  assign n152 = n150 & ~n151 ;
  assign n153 = ~n144 & n152 ;
  assign n154 = n144 & ~n152 ;
  assign n155 = n153 | n154 ;
  assign n156 = n143 | n155 ;
  assign n157 = n143 & n155 ;
  assign n158 = n156 & ~n157 ;
  assign n159 = ~n142 & n158 ;
  assign n160 = n142 & ~n158 ;
  assign n161 = n159 | n160 ;
  assign n162 = n141 | n161 ;
  assign n163 = n141 & n161 ;
  assign n164 = n162 & ~n163 ;
  assign n165 = ~n140 & n164 ;
  assign n166 = n140 & ~n164 ;
  assign n167 = n165 | n166 ;
  assign n168 = n139 | n167 ;
  assign n169 = n139 & n167 ;
  assign n170 = n168 & ~n169 ;
  assign n171 = ~n138 & n170 ;
  assign n172 = n138 & ~n170 ;
  assign n173 = n171 | n172 ;
  assign n174 = n137 | n173 ;
  assign n175 = n137 & n173 ;
  assign n176 = n174 & ~n175 ;
  assign n177 = ~n136 & n176 ;
  assign n178 = n136 & ~n176 ;
  assign n179 = n177 | n178 ;
  assign n180 = N1 & N392 ;
  assign n181 = n174 & ~n177 ;
  assign n182 = N18 & N375 ;
  assign n183 = n168 & ~n171 ;
  assign n184 = N35 & N358 ;
  assign n185 = n162 & ~n165 ;
  assign n186 = N341 & N52 ;
  assign n187 = n156 & ~n159 ;
  assign n188 = N324 & N69 ;
  assign n189 = n150 & ~n153 ;
  assign n190 = N307 & N86 ;
  assign n191 = N120 & N290 ;
  assign n192 = n147 & n191 ;
  assign n193 = N120 & N273 ;
  assign n194 = n145 | n193 ;
  assign n195 = ~n192 & n194 ;
  assign n196 = n146 | n195 ;
  assign n197 = n146 & n195 ;
  assign n198 = n196 & ~n197 ;
  assign n199 = ~n190 & n198 ;
  assign n200 = n190 & ~n198 ;
  assign n201 = n199 | n200 ;
  assign n202 = n189 | n201 ;
  assign n203 = n189 & n201 ;
  assign n204 = n202 & ~n203 ;
  assign n205 = ~n188 & n204 ;
  assign n206 = n188 & ~n204 ;
  assign n207 = n205 | n206 ;
  assign n208 = n187 | n207 ;
  assign n209 = n187 & n207 ;
  assign n210 = n208 & ~n209 ;
  assign n211 = ~n186 & n210 ;
  assign n212 = n186 & ~n210 ;
  assign n213 = n211 | n212 ;
  assign n214 = n185 | n213 ;
  assign n215 = n185 & n213 ;
  assign n216 = n214 & ~n215 ;
  assign n217 = ~n184 & n216 ;
  assign n218 = n184 & ~n216 ;
  assign n219 = n217 | n218 ;
  assign n220 = n183 | n219 ;
  assign n221 = n183 & n219 ;
  assign n222 = n220 & ~n221 ;
  assign n223 = ~n182 & n222 ;
  assign n224 = n182 & ~n222 ;
  assign n225 = n223 | n224 ;
  assign n226 = n181 | n225 ;
  assign n227 = n181 & n225 ;
  assign n228 = n226 & ~n227 ;
  assign n229 = ~n180 & n228 ;
  assign n230 = n180 & ~n228 ;
  assign n231 = n229 | n230 ;
  assign n232 = N1 & N409 ;
  assign n233 = n226 & ~n229 ;
  assign n234 = N18 & N392 ;
  assign n235 = n220 & ~n223 ;
  assign n236 = N35 & N375 ;
  assign n237 = n214 & ~n217 ;
  assign n238 = N358 & N52 ;
  assign n239 = n208 & ~n211 ;
  assign n240 = N341 & N69 ;
  assign n241 = n202 & ~n205 ;
  assign n242 = N324 & N86 ;
  assign n243 = n196 & ~n199 ;
  assign n244 = N103 & N307 ;
  assign n245 = N137 & N290 ;
  assign n246 = n193 & n245 ;
  assign n247 = N137 & N273 ;
  assign n248 = n191 | n247 ;
  assign n249 = ~n246 & n248 ;
  assign n250 = n192 | n249 ;
  assign n251 = n192 & n249 ;
  assign n252 = n250 & ~n251 ;
  assign n253 = ~n244 & n252 ;
  assign n254 = n244 & ~n252 ;
  assign n255 = n253 | n254 ;
  assign n256 = n243 | n255 ;
  assign n257 = n243 & n255 ;
  assign n258 = n256 & ~n257 ;
  assign n259 = ~n242 & n258 ;
  assign n260 = n242 & ~n258 ;
  assign n261 = n259 | n260 ;
  assign n262 = n241 | n261 ;
  assign n263 = n241 & n261 ;
  assign n264 = n262 & ~n263 ;
  assign n265 = ~n240 & n264 ;
  assign n266 = n240 & ~n264 ;
  assign n267 = n265 | n266 ;
  assign n268 = n239 | n267 ;
  assign n269 = n239 & n267 ;
  assign n270 = n268 & ~n269 ;
  assign n271 = ~n238 & n270 ;
  assign n272 = n238 & ~n270 ;
  assign n273 = n271 | n272 ;
  assign n274 = n237 | n273 ;
  assign n275 = n237 & n273 ;
  assign n276 = n274 & ~n275 ;
  assign n277 = ~n236 & n276 ;
  assign n278 = n236 & ~n276 ;
  assign n279 = n277 | n278 ;
  assign n280 = n235 | n279 ;
  assign n281 = n235 & n279 ;
  assign n282 = n280 & ~n281 ;
  assign n283 = ~n234 & n282 ;
  assign n284 = n234 & ~n282 ;
  assign n285 = n283 | n284 ;
  assign n286 = n233 | n285 ;
  assign n287 = n233 & n285 ;
  assign n288 = n286 & ~n287 ;
  assign n289 = ~n232 & n288 ;
  assign n290 = n232 & ~n288 ;
  assign n291 = n289 | n290 ;
  assign n292 = N1 & N426 ;
  assign n293 = n286 & ~n289 ;
  assign n294 = N18 & N409 ;
  assign n295 = n280 & ~n283 ;
  assign n296 = N35 & N392 ;
  assign n297 = n274 & ~n277 ;
  assign n298 = N375 & N52 ;
  assign n299 = n268 & ~n271 ;
  assign n300 = N358 & N69 ;
  assign n301 = n262 & ~n265 ;
  assign n302 = N341 & N86 ;
  assign n303 = n256 & ~n259 ;
  assign n304 = N103 & N324 ;
  assign n305 = n250 & ~n253 ;
  assign n306 = N120 & N307 ;
  assign n307 = N154 & N290 ;
  assign n308 = n247 & n307 ;
  assign n309 = N154 & N273 ;
  assign n310 = n245 | n309 ;
  assign n311 = ~n308 & n310 ;
  assign n312 = n246 | n311 ;
  assign n313 = n246 & n311 ;
  assign n314 = n312 & ~n313 ;
  assign n315 = ~n306 & n314 ;
  assign n316 = n306 & ~n314 ;
  assign n317 = n315 | n316 ;
  assign n318 = n305 | n317 ;
  assign n319 = n305 & n317 ;
  assign n320 = n318 & ~n319 ;
  assign n321 = ~n304 & n320 ;
  assign n322 = n304 & ~n320 ;
  assign n323 = n321 | n322 ;
  assign n324 = n303 | n323 ;
  assign n325 = n303 & n323 ;
  assign n326 = n324 & ~n325 ;
  assign n327 = ~n302 & n326 ;
  assign n328 = n302 & ~n326 ;
  assign n329 = n327 | n328 ;
  assign n330 = n301 | n329 ;
  assign n331 = n301 & n329 ;
  assign n332 = n330 & ~n331 ;
  assign n333 = ~n300 & n332 ;
  assign n334 = n300 & ~n332 ;
  assign n335 = n333 | n334 ;
  assign n336 = n299 | n335 ;
  assign n337 = n299 & n335 ;
  assign n338 = n336 & ~n337 ;
  assign n339 = ~n298 & n338 ;
  assign n340 = n298 & ~n338 ;
  assign n341 = n339 | n340 ;
  assign n342 = n297 | n341 ;
  assign n343 = n297 & n341 ;
  assign n344 = n342 & ~n343 ;
  assign n345 = ~n296 & n344 ;
  assign n346 = n296 & ~n344 ;
  assign n347 = n345 | n346 ;
  assign n348 = n295 | n347 ;
  assign n349 = n295 & n347 ;
  assign n350 = n348 & ~n349 ;
  assign n351 = ~n294 & n350 ;
  assign n352 = n294 & ~n350 ;
  assign n353 = n351 | n352 ;
  assign n354 = n293 | n353 ;
  assign n355 = n293 & n353 ;
  assign n356 = n354 & ~n355 ;
  assign n357 = ~n292 & n356 ;
  assign n358 = n292 & ~n356 ;
  assign n359 = n357 | n358 ;
  assign n360 = N1 & N443 ;
  assign n361 = n354 & ~n357 ;
  assign n362 = N18 & N426 ;
  assign n363 = n348 & ~n351 ;
  assign n364 = N35 & N409 ;
  assign n365 = n342 & ~n345 ;
  assign n366 = N392 & N52 ;
  assign n367 = n336 & ~n339 ;
  assign n368 = N375 & N69 ;
  assign n369 = n330 & ~n333 ;
  assign n370 = N358 & N86 ;
  assign n371 = n324 & ~n327 ;
  assign n372 = N103 & N341 ;
  assign n373 = n318 & ~n321 ;
  assign n374 = N120 & N324 ;
  assign n375 = n312 & ~n315 ;
  assign n376 = N137 & N307 ;
  assign n377 = N171 & N290 ;
  assign n378 = n309 & n377 ;
  assign n379 = N171 & N273 ;
  assign n380 = n307 | n379 ;
  assign n381 = ~n378 & n380 ;
  assign n382 = n308 | n381 ;
  assign n383 = n308 & n381 ;
  assign n384 = n382 & ~n383 ;
  assign n385 = ~n376 & n384 ;
  assign n386 = n376 & ~n384 ;
  assign n387 = n385 | n386 ;
  assign n388 = n375 | n387 ;
  assign n389 = n375 & n387 ;
  assign n390 = n388 & ~n389 ;
  assign n391 = ~n374 & n390 ;
  assign n392 = n374 & ~n390 ;
  assign n393 = n391 | n392 ;
  assign n394 = n373 | n393 ;
  assign n395 = n373 & n393 ;
  assign n396 = n394 & ~n395 ;
  assign n397 = ~n372 & n396 ;
  assign n398 = n372 & ~n396 ;
  assign n399 = n397 | n398 ;
  assign n400 = n371 | n399 ;
  assign n401 = n371 & n399 ;
  assign n402 = n400 & ~n401 ;
  assign n403 = ~n370 & n402 ;
  assign n404 = n370 & ~n402 ;
  assign n405 = n403 | n404 ;
  assign n406 = n369 | n405 ;
  assign n407 = n369 & n405 ;
  assign n408 = n406 & ~n407 ;
  assign n409 = ~n368 & n408 ;
  assign n410 = n368 & ~n408 ;
  assign n411 = n409 | n410 ;
  assign n412 = n367 | n411 ;
  assign n413 = n367 & n411 ;
  assign n414 = n412 & ~n413 ;
  assign n415 = ~n366 & n414 ;
  assign n416 = n366 & ~n414 ;
  assign n417 = n415 | n416 ;
  assign n418 = n365 | n417 ;
  assign n419 = n365 & n417 ;
  assign n420 = n418 & ~n419 ;
  assign n421 = ~n364 & n420 ;
  assign n422 = n364 & ~n420 ;
  assign n423 = n421 | n422 ;
  assign n424 = n363 | n423 ;
  assign n425 = n363 & n423 ;
  assign n426 = n424 & ~n425 ;
  assign n427 = ~n362 & n426 ;
  assign n428 = n362 & ~n426 ;
  assign n429 = n427 | n428 ;
  assign n430 = n361 | n429 ;
  assign n431 = n361 & n429 ;
  assign n432 = n430 & ~n431 ;
  assign n433 = ~n360 & n432 ;
  assign n434 = n360 & ~n432 ;
  assign n435 = n433 | n434 ;
  assign n436 = N1 & N460 ;
  assign n437 = n430 & ~n433 ;
  assign n438 = N18 & N443 ;
  assign n439 = n424 & ~n427 ;
  assign n440 = N35 & N426 ;
  assign n441 = n418 & ~n421 ;
  assign n442 = N409 & N52 ;
  assign n443 = n412 & ~n415 ;
  assign n444 = N392 & N69 ;
  assign n445 = n406 & ~n409 ;
  assign n446 = N375 & N86 ;
  assign n447 = n400 & ~n403 ;
  assign n448 = N103 & N358 ;
  assign n449 = n394 & ~n397 ;
  assign n450 = N120 & N341 ;
  assign n451 = n388 & ~n391 ;
  assign n452 = N137 & N324 ;
  assign n453 = n382 & ~n385 ;
  assign n454 = N154 & N307 ;
  assign n455 = N188 & N290 ;
  assign n456 = n379 & n455 ;
  assign n457 = N188 & N273 ;
  assign n458 = n377 | n457 ;
  assign n459 = ~n456 & n458 ;
  assign n460 = n378 | n459 ;
  assign n461 = n378 & n459 ;
  assign n462 = n460 & ~n461 ;
  assign n463 = ~n454 & n462 ;
  assign n464 = n454 & ~n462 ;
  assign n465 = n463 | n464 ;
  assign n466 = n453 | n465 ;
  assign n467 = n453 & n465 ;
  assign n468 = n466 & ~n467 ;
  assign n469 = ~n452 & n468 ;
  assign n470 = n452 & ~n468 ;
  assign n471 = n469 | n470 ;
  assign n472 = n451 | n471 ;
  assign n473 = n451 & n471 ;
  assign n474 = n472 & ~n473 ;
  assign n475 = ~n450 & n474 ;
  assign n476 = n450 & ~n474 ;
  assign n477 = n475 | n476 ;
  assign n478 = n449 | n477 ;
  assign n479 = n449 & n477 ;
  assign n480 = n478 & ~n479 ;
  assign n481 = ~n448 & n480 ;
  assign n482 = n448 & ~n480 ;
  assign n483 = n481 | n482 ;
  assign n484 = n447 | n483 ;
  assign n485 = n447 & n483 ;
  assign n486 = n484 & ~n485 ;
  assign n487 = ~n446 & n486 ;
  assign n488 = n446 & ~n486 ;
  assign n489 = n487 | n488 ;
  assign n490 = n445 | n489 ;
  assign n491 = n445 & n489 ;
  assign n492 = n490 & ~n491 ;
  assign n493 = ~n444 & n492 ;
  assign n494 = n444 & ~n492 ;
  assign n495 = n493 | n494 ;
  assign n496 = n443 | n495 ;
  assign n497 = n443 & n495 ;
  assign n498 = n496 & ~n497 ;
  assign n499 = ~n442 & n498 ;
  assign n500 = n442 & ~n498 ;
  assign n501 = n499 | n500 ;
  assign n502 = n441 | n501 ;
  assign n503 = n441 & n501 ;
  assign n504 = n502 & ~n503 ;
  assign n505 = ~n440 & n504 ;
  assign n506 = n440 & ~n504 ;
  assign n507 = n505 | n506 ;
  assign n508 = n439 | n507 ;
  assign n509 = n439 & n507 ;
  assign n510 = n508 & ~n509 ;
  assign n511 = ~n438 & n510 ;
  assign n512 = n438 & ~n510 ;
  assign n513 = n511 | n512 ;
  assign n514 = n437 | n513 ;
  assign n515 = n437 & n513 ;
  assign n516 = n514 & ~n515 ;
  assign n517 = ~n436 & n516 ;
  assign n518 = n436 & ~n516 ;
  assign n519 = n517 | n518 ;
  assign n520 = N1 & N477 ;
  assign n521 = n514 & ~n517 ;
  assign n522 = N18 & N460 ;
  assign n523 = n508 & ~n511 ;
  assign n524 = N35 & N443 ;
  assign n525 = n502 & ~n505 ;
  assign n526 = N426 & N52 ;
  assign n527 = n496 & ~n499 ;
  assign n528 = N409 & N69 ;
  assign n529 = n490 & ~n493 ;
  assign n530 = N392 & N86 ;
  assign n531 = n484 & ~n487 ;
  assign n532 = N103 & N375 ;
  assign n533 = n478 & ~n481 ;
  assign n534 = N120 & N358 ;
  assign n535 = n472 & ~n475 ;
  assign n536 = N137 & N341 ;
  assign n537 = n466 & ~n469 ;
  assign n538 = N154 & N324 ;
  assign n539 = n460 & ~n463 ;
  assign n540 = N171 & N307 ;
  assign n541 = N205 & N290 ;
  assign n542 = n457 & n541 ;
  assign n543 = N205 & N273 ;
  assign n544 = n455 | n543 ;
  assign n545 = ~n542 & n544 ;
  assign n546 = n456 | n545 ;
  assign n547 = n456 & n545 ;
  assign n548 = n546 & ~n547 ;
  assign n549 = ~n540 & n548 ;
  assign n550 = n540 & ~n548 ;
  assign n551 = n549 | n550 ;
  assign n552 = n539 | n551 ;
  assign n553 = n539 & n551 ;
  assign n554 = n552 & ~n553 ;
  assign n555 = ~n538 & n554 ;
  assign n556 = n538 & ~n554 ;
  assign n557 = n555 | n556 ;
  assign n558 = n537 | n557 ;
  assign n559 = n537 & n557 ;
  assign n560 = n558 & ~n559 ;
  assign n561 = ~n536 & n560 ;
  assign n562 = n536 & ~n560 ;
  assign n563 = n561 | n562 ;
  assign n564 = n535 | n563 ;
  assign n565 = n535 & n563 ;
  assign n566 = n564 & ~n565 ;
  assign n567 = ~n534 & n566 ;
  assign n568 = n534 & ~n566 ;
  assign n569 = n567 | n568 ;
  assign n570 = n533 | n569 ;
  assign n571 = n533 & n569 ;
  assign n572 = n570 & ~n571 ;
  assign n573 = ~n532 & n572 ;
  assign n574 = n532 & ~n572 ;
  assign n575 = n573 | n574 ;
  assign n576 = n531 | n575 ;
  assign n577 = n531 & n575 ;
  assign n578 = n576 & ~n577 ;
  assign n579 = ~n530 & n578 ;
  assign n580 = n530 & ~n578 ;
  assign n581 = n579 | n580 ;
  assign n582 = n529 | n581 ;
  assign n583 = n529 & n581 ;
  assign n584 = n582 & ~n583 ;
  assign n585 = ~n528 & n584 ;
  assign n586 = n528 & ~n584 ;
  assign n587 = n585 | n586 ;
  assign n588 = n527 | n587 ;
  assign n589 = n527 & n587 ;
  assign n590 = n588 & ~n589 ;
  assign n591 = ~n526 & n590 ;
  assign n592 = n526 & ~n590 ;
  assign n593 = n591 | n592 ;
  assign n594 = n525 | n593 ;
  assign n595 = n525 & n593 ;
  assign n596 = n594 & ~n595 ;
  assign n597 = ~n524 & n596 ;
  assign n598 = n524 & ~n596 ;
  assign n599 = n597 | n598 ;
  assign n600 = n523 | n599 ;
  assign n601 = n523 & n599 ;
  assign n602 = n600 & ~n601 ;
  assign n603 = ~n522 & n602 ;
  assign n604 = n522 & ~n602 ;
  assign n605 = n603 | n604 ;
  assign n606 = n521 | n605 ;
  assign n607 = n521 & n605 ;
  assign n608 = n606 & ~n607 ;
  assign n609 = ~n520 & n608 ;
  assign n610 = n520 & ~n608 ;
  assign n611 = n609 | n610 ;
  assign n612 = N1 & N494 ;
  assign n613 = n606 & ~n609 ;
  assign n614 = N18 & N477 ;
  assign n615 = n600 & ~n603 ;
  assign n616 = N35 & N460 ;
  assign n617 = n594 & ~n597 ;
  assign n618 = N443 & N52 ;
  assign n619 = n588 & ~n591 ;
  assign n620 = N426 & N69 ;
  assign n621 = n582 & ~n585 ;
  assign n622 = N409 & N86 ;
  assign n623 = n576 & ~n579 ;
  assign n624 = N103 & N392 ;
  assign n625 = n570 & ~n573 ;
  assign n626 = N120 & N375 ;
  assign n627 = n564 & ~n567 ;
  assign n628 = N137 & N358 ;
  assign n629 = n558 & ~n561 ;
  assign n630 = N154 & N341 ;
  assign n631 = n552 & ~n555 ;
  assign n632 = N171 & N324 ;
  assign n633 = n546 & ~n549 ;
  assign n634 = N188 & N307 ;
  assign n635 = N222 & N290 ;
  assign n636 = n543 & n635 ;
  assign n637 = N222 & N273 ;
  assign n638 = n541 | n637 ;
  assign n639 = ~n636 & n638 ;
  assign n640 = n542 | n639 ;
  assign n641 = n542 & n639 ;
  assign n642 = n640 & ~n641 ;
  assign n643 = ~n634 & n642 ;
  assign n644 = n634 & ~n642 ;
  assign n645 = n643 | n644 ;
  assign n646 = n633 | n645 ;
  assign n647 = n633 & n645 ;
  assign n648 = n646 & ~n647 ;
  assign n649 = ~n632 & n648 ;
  assign n650 = n632 & ~n648 ;
  assign n651 = n649 | n650 ;
  assign n652 = n631 | n651 ;
  assign n653 = n631 & n651 ;
  assign n654 = n652 & ~n653 ;
  assign n655 = ~n630 & n654 ;
  assign n656 = n630 & ~n654 ;
  assign n657 = n655 | n656 ;
  assign n658 = n629 | n657 ;
  assign n659 = n629 & n657 ;
  assign n660 = n658 & ~n659 ;
  assign n661 = ~n628 & n660 ;
  assign n662 = n628 & ~n660 ;
  assign n663 = n661 | n662 ;
  assign n664 = n627 | n663 ;
  assign n665 = n627 & n663 ;
  assign n666 = n664 & ~n665 ;
  assign n667 = ~n626 & n666 ;
  assign n668 = n626 & ~n666 ;
  assign n669 = n667 | n668 ;
  assign n670 = n625 | n669 ;
  assign n671 = n625 & n669 ;
  assign n672 = n670 & ~n671 ;
  assign n673 = ~n624 & n672 ;
  assign n674 = n624 & ~n672 ;
  assign n675 = n673 | n674 ;
  assign n676 = n623 | n675 ;
  assign n677 = n623 & n675 ;
  assign n678 = n676 & ~n677 ;
  assign n679 = ~n622 & n678 ;
  assign n680 = n622 & ~n678 ;
  assign n681 = n679 | n680 ;
  assign n682 = n621 | n681 ;
  assign n683 = n621 & n681 ;
  assign n684 = n682 & ~n683 ;
  assign n685 = ~n620 & n684 ;
  assign n686 = n620 & ~n684 ;
  assign n687 = n685 | n686 ;
  assign n688 = n619 | n687 ;
  assign n689 = n619 & n687 ;
  assign n690 = n688 & ~n689 ;
  assign n691 = ~n618 & n690 ;
  assign n692 = n618 & ~n690 ;
  assign n693 = n691 | n692 ;
  assign n694 = n617 | n693 ;
  assign n695 = n617 & n693 ;
  assign n696 = n694 & ~n695 ;
  assign n697 = ~n616 & n696 ;
  assign n698 = n616 & ~n696 ;
  assign n699 = n697 | n698 ;
  assign n700 = n615 | n699 ;
  assign n701 = n615 & n699 ;
  assign n702 = n700 & ~n701 ;
  assign n703 = ~n614 & n702 ;
  assign n704 = n614 & ~n702 ;
  assign n705 = n703 | n704 ;
  assign n706 = n613 | n705 ;
  assign n707 = n613 & n705 ;
  assign n708 = n706 & ~n707 ;
  assign n709 = ~n612 & n708 ;
  assign n710 = n612 & ~n708 ;
  assign n711 = n709 | n710 ;
  assign n712 = N1 & N511 ;
  assign n713 = n706 & ~n709 ;
  assign n714 = N18 & N494 ;
  assign n715 = n700 & ~n703 ;
  assign n716 = N35 & N477 ;
  assign n717 = n694 & ~n697 ;
  assign n718 = N460 & N52 ;
  assign n719 = n688 & ~n691 ;
  assign n720 = N443 & N69 ;
  assign n721 = n682 & ~n685 ;
  assign n722 = N426 & N86 ;
  assign n723 = n676 & ~n679 ;
  assign n724 = N103 & N409 ;
  assign n725 = n670 & ~n673 ;
  assign n726 = N120 & N392 ;
  assign n727 = n664 & ~n667 ;
  assign n728 = N137 & N375 ;
  assign n729 = n658 & ~n661 ;
  assign n730 = N154 & N358 ;
  assign n731 = n652 & ~n655 ;
  assign n732 = N171 & N341 ;
  assign n733 = n646 & ~n649 ;
  assign n734 = N188 & N324 ;
  assign n735 = n640 & ~n643 ;
  assign n736 = N205 & N307 ;
  assign n737 = N239 & N290 ;
  assign n738 = n637 & n737 ;
  assign n739 = N239 & N273 ;
  assign n740 = n635 | n739 ;
  assign n741 = ~n738 & n740 ;
  assign n742 = n636 | n741 ;
  assign n743 = n636 & n741 ;
  assign n744 = n742 & ~n743 ;
  assign n745 = ~n736 & n744 ;
  assign n746 = n736 & ~n744 ;
  assign n747 = n745 | n746 ;
  assign n748 = n735 | n747 ;
  assign n749 = n735 & n747 ;
  assign n750 = n748 & ~n749 ;
  assign n751 = ~n734 & n750 ;
  assign n752 = n734 & ~n750 ;
  assign n753 = n751 | n752 ;
  assign n754 = n733 | n753 ;
  assign n755 = n733 & n753 ;
  assign n756 = n754 & ~n755 ;
  assign n757 = ~n732 & n756 ;
  assign n758 = n732 & ~n756 ;
  assign n759 = n757 | n758 ;
  assign n760 = n731 | n759 ;
  assign n761 = n731 & n759 ;
  assign n762 = n760 & ~n761 ;
  assign n763 = ~n730 & n762 ;
  assign n764 = n730 & ~n762 ;
  assign n765 = n763 | n764 ;
  assign n766 = n729 | n765 ;
  assign n767 = n729 & n765 ;
  assign n768 = n766 & ~n767 ;
  assign n769 = ~n728 & n768 ;
  assign n770 = n728 & ~n768 ;
  assign n771 = n769 | n770 ;
  assign n772 = n727 | n771 ;
  assign n773 = n727 & n771 ;
  assign n774 = n772 & ~n773 ;
  assign n775 = ~n726 & n774 ;
  assign n776 = n726 & ~n774 ;
  assign n777 = n775 | n776 ;
  assign n778 = n725 | n777 ;
  assign n779 = n725 & n777 ;
  assign n780 = n778 & ~n779 ;
  assign n781 = ~n724 & n780 ;
  assign n782 = n724 & ~n780 ;
  assign n783 = n781 | n782 ;
  assign n784 = n723 | n783 ;
  assign n785 = n723 & n783 ;
  assign n786 = n784 & ~n785 ;
  assign n787 = ~n722 & n786 ;
  assign n788 = n722 & ~n786 ;
  assign n789 = n787 | n788 ;
  assign n790 = n721 | n789 ;
  assign n791 = n721 & n789 ;
  assign n792 = n790 & ~n791 ;
  assign n793 = ~n720 & n792 ;
  assign n794 = n720 & ~n792 ;
  assign n795 = n793 | n794 ;
  assign n796 = n719 | n795 ;
  assign n797 = n719 & n795 ;
  assign n798 = n796 & ~n797 ;
  assign n799 = ~n718 & n798 ;
  assign n800 = n718 & ~n798 ;
  assign n801 = n799 | n800 ;
  assign n802 = n717 | n801 ;
  assign n803 = n717 & n801 ;
  assign n804 = n802 & ~n803 ;
  assign n805 = ~n716 & n804 ;
  assign n806 = n716 & ~n804 ;
  assign n807 = n805 | n806 ;
  assign n808 = n715 | n807 ;
  assign n809 = n715 & n807 ;
  assign n810 = n808 & ~n809 ;
  assign n811 = ~n714 & n810 ;
  assign n812 = n714 & ~n810 ;
  assign n813 = n811 | n812 ;
  assign n814 = n713 | n813 ;
  assign n815 = n713 & n813 ;
  assign n816 = n814 & ~n815 ;
  assign n817 = ~n712 & n816 ;
  assign n818 = n712 & ~n816 ;
  assign n819 = n817 | n818 ;
  assign n820 = N1 & N528 ;
  assign n821 = n814 & ~n817 ;
  assign n822 = N18 & N511 ;
  assign n823 = n808 & ~n811 ;
  assign n824 = N35 & N494 ;
  assign n825 = n802 & ~n805 ;
  assign n826 = N477 & N52 ;
  assign n827 = n796 & ~n799 ;
  assign n828 = N460 & N69 ;
  assign n829 = n790 & ~n793 ;
  assign n830 = N443 & N86 ;
  assign n831 = n784 & ~n787 ;
  assign n832 = N103 & N426 ;
  assign n833 = n778 & ~n781 ;
  assign n834 = N120 & N409 ;
  assign n835 = n772 & ~n775 ;
  assign n836 = N137 & N392 ;
  assign n837 = n766 & ~n769 ;
  assign n838 = N154 & N375 ;
  assign n839 = n760 & ~n763 ;
  assign n840 = N171 & N358 ;
  assign n841 = n754 & ~n757 ;
  assign n842 = N188 & N341 ;
  assign n843 = n748 & ~n751 ;
  assign n844 = N205 & N324 ;
  assign n845 = n742 & ~n745 ;
  assign n846 = N222 & N307 ;
  assign n847 = ~N256 & n738 ;
  assign n848 = N256 & N273 ;
  assign n849 = n737 | n848 ;
  assign n850 = ~N222 & n737 ;
  assign n851 = n848 & n850 ;
  assign n852 = n849 & ~n851 ;
  assign n853 = ~n847 & n852 ;
  assign n854 = ~n846 & n853 ;
  assign n855 = n846 & ~n853 ;
  assign n856 = n854 | n855 ;
  assign n857 = n845 | n856 ;
  assign n858 = n845 & n856 ;
  assign n859 = n857 & ~n858 ;
  assign n860 = ~n844 & n859 ;
  assign n861 = n844 & ~n859 ;
  assign n862 = n860 | n861 ;
  assign n863 = n843 | n862 ;
  assign n864 = n843 & n862 ;
  assign n865 = n863 & ~n864 ;
  assign n866 = ~n842 & n865 ;
  assign n867 = n842 & ~n865 ;
  assign n868 = n866 | n867 ;
  assign n869 = n841 | n868 ;
  assign n870 = n841 & n868 ;
  assign n871 = n869 & ~n870 ;
  assign n872 = ~n840 & n871 ;
  assign n873 = n840 & ~n871 ;
  assign n874 = n872 | n873 ;
  assign n875 = n839 | n874 ;
  assign n876 = n839 & n874 ;
  assign n877 = n875 & ~n876 ;
  assign n878 = ~n838 & n877 ;
  assign n879 = n838 & ~n877 ;
  assign n880 = n878 | n879 ;
  assign n881 = n837 | n880 ;
  assign n882 = n837 & n880 ;
  assign n883 = n881 & ~n882 ;
  assign n884 = ~n836 & n883 ;
  assign n885 = n836 & ~n883 ;
  assign n886 = n884 | n885 ;
  assign n887 = n835 | n886 ;
  assign n888 = n835 & n886 ;
  assign n889 = n887 & ~n888 ;
  assign n890 = ~n834 & n889 ;
  assign n891 = n834 & ~n889 ;
  assign n892 = n890 | n891 ;
  assign n893 = n833 | n892 ;
  assign n894 = n833 & n892 ;
  assign n895 = n893 & ~n894 ;
  assign n896 = ~n832 & n895 ;
  assign n897 = n832 & ~n895 ;
  assign n898 = n896 | n897 ;
  assign n899 = n831 | n898 ;
  assign n900 = n831 & n898 ;
  assign n901 = n899 & ~n900 ;
  assign n902 = ~n830 & n901 ;
  assign n903 = n830 & ~n901 ;
  assign n904 = n902 | n903 ;
  assign n905 = n829 | n904 ;
  assign n906 = n829 & n904 ;
  assign n907 = n905 & ~n906 ;
  assign n908 = ~n828 & n907 ;
  assign n909 = n828 & ~n907 ;
  assign n910 = n908 | n909 ;
  assign n911 = n827 | n910 ;
  assign n912 = n827 & n910 ;
  assign n913 = n911 & ~n912 ;
  assign n914 = ~n826 & n913 ;
  assign n915 = n826 & ~n913 ;
  assign n916 = n914 | n915 ;
  assign n917 = n825 | n916 ;
  assign n918 = n825 & n916 ;
  assign n919 = n917 & ~n918 ;
  assign n920 = ~n824 & n919 ;
  assign n921 = n824 & ~n919 ;
  assign n922 = n920 | n921 ;
  assign n923 = n823 | n922 ;
  assign n924 = n823 & n922 ;
  assign n925 = n923 & ~n924 ;
  assign n926 = ~n822 & n925 ;
  assign n927 = n822 & ~n925 ;
  assign n928 = n926 | n927 ;
  assign n929 = n821 | n928 ;
  assign n930 = n821 & n928 ;
  assign n931 = n929 & ~n930 ;
  assign n932 = ~n820 & n931 ;
  assign n933 = n820 & ~n931 ;
  assign n934 = n932 | n933 ;
  assign n935 = n929 & ~n932 ;
  assign n936 = N18 & N528 ;
  assign n937 = n923 & ~n926 ;
  assign n938 = N35 & N511 ;
  assign n939 = n917 & ~n920 ;
  assign n940 = N494 & N52 ;
  assign n941 = n911 & ~n914 ;
  assign n942 = N477 & N69 ;
  assign n943 = n905 & ~n908 ;
  assign n944 = N460 & N86 ;
  assign n945 = n899 & ~n902 ;
  assign n946 = N103 & N443 ;
  assign n947 = n893 & ~n896 ;
  assign n948 = N120 & N426 ;
  assign n949 = n887 & ~n890 ;
  assign n950 = N137 & N409 ;
  assign n951 = n881 & ~n884 ;
  assign n952 = N154 & N392 ;
  assign n953 = n875 & ~n878 ;
  assign n954 = N171 & N375 ;
  assign n955 = n869 & ~n872 ;
  assign n956 = N188 & N358 ;
  assign n957 = n863 & ~n866 ;
  assign n958 = N205 & N341 ;
  assign n959 = n857 & ~n860 ;
  assign n960 = N222 & N324 ;
  assign n961 = n852 & ~n854 ;
  assign n962 = N256 & N290 ;
  assign n963 = ~n739 & n962 ;
  assign n964 = N239 & N307 ;
  assign n965 = n963 & ~n964 ;
  assign n966 = ~n963 & n964 ;
  assign n967 = n965 | n966 ;
  assign n968 = n961 | n967 ;
  assign n969 = n961 & n967 ;
  assign n970 = n968 & ~n969 ;
  assign n971 = ~n960 & n970 ;
  assign n972 = n960 & ~n970 ;
  assign n973 = n971 | n972 ;
  assign n974 = n959 | n973 ;
  assign n975 = n959 & n973 ;
  assign n976 = n974 & ~n975 ;
  assign n977 = ~n958 & n976 ;
  assign n978 = n958 & ~n976 ;
  assign n979 = n977 | n978 ;
  assign n980 = n957 | n979 ;
  assign n981 = n957 & n979 ;
  assign n982 = n980 & ~n981 ;
  assign n983 = ~n956 & n982 ;
  assign n984 = n956 & ~n982 ;
  assign n985 = n983 | n984 ;
  assign n986 = n955 | n985 ;
  assign n987 = n955 & n985 ;
  assign n988 = n986 & ~n987 ;
  assign n989 = ~n954 & n988 ;
  assign n990 = n954 & ~n988 ;
  assign n991 = n989 | n990 ;
  assign n992 = n953 | n991 ;
  assign n993 = n953 & n991 ;
  assign n994 = n992 & ~n993 ;
  assign n995 = ~n952 & n994 ;
  assign n996 = n952 & ~n994 ;
  assign n997 = n995 | n996 ;
  assign n998 = n951 | n997 ;
  assign n999 = n951 & n997 ;
  assign n1000 = n998 & ~n999 ;
  assign n1001 = ~n950 & n1000 ;
  assign n1002 = n950 & ~n1000 ;
  assign n1003 = n1001 | n1002 ;
  assign n1004 = n949 | n1003 ;
  assign n1005 = n949 & n1003 ;
  assign n1006 = n1004 & ~n1005 ;
  assign n1007 = ~n948 & n1006 ;
  assign n1008 = n948 & ~n1006 ;
  assign n1009 = n1007 | n1008 ;
  assign n1010 = n947 | n1009 ;
  assign n1011 = n947 & n1009 ;
  assign n1012 = n1010 & ~n1011 ;
  assign n1013 = ~n946 & n1012 ;
  assign n1014 = n946 & ~n1012 ;
  assign n1015 = n1013 | n1014 ;
  assign n1016 = n945 | n1015 ;
  assign n1017 = n945 & n1015 ;
  assign n1018 = n1016 & ~n1017 ;
  assign n1019 = ~n944 & n1018 ;
  assign n1020 = n944 & ~n1018 ;
  assign n1021 = n1019 | n1020 ;
  assign n1022 = n943 | n1021 ;
  assign n1023 = n943 & n1021 ;
  assign n1024 = n1022 & ~n1023 ;
  assign n1025 = ~n942 & n1024 ;
  assign n1026 = n942 & ~n1024 ;
  assign n1027 = n1025 | n1026 ;
  assign n1028 = n941 | n1027 ;
  assign n1029 = n941 & n1027 ;
  assign n1030 = n1028 & ~n1029 ;
  assign n1031 = ~n940 & n1030 ;
  assign n1032 = n940 & ~n1030 ;
  assign n1033 = n1031 | n1032 ;
  assign n1034 = n939 | n1033 ;
  assign n1035 = n939 & n1033 ;
  assign n1036 = n1034 & ~n1035 ;
  assign n1037 = ~n938 & n1036 ;
  assign n1038 = n938 & ~n1036 ;
  assign n1039 = n1037 | n1038 ;
  assign n1040 = n937 | n1039 ;
  assign n1041 = n937 & n1039 ;
  assign n1042 = n1040 & ~n1041 ;
  assign n1043 = ~n936 & n1042 ;
  assign n1044 = n936 & ~n1042 ;
  assign n1045 = n1043 | n1044 ;
  assign n1046 = n935 & n1045 ;
  assign n1047 = n935 | n1045 ;
  assign n1048 = ~n1046 & n1047 ;
  assign n1049 = n1040 & ~n1043 ;
  assign n1050 = N35 & N528 ;
  assign n1051 = n1034 & ~n1037 ;
  assign n1052 = N511 & N52 ;
  assign n1053 = n1028 & ~n1031 ;
  assign n1054 = N494 & N69 ;
  assign n1055 = n1022 & ~n1025 ;
  assign n1056 = N477 & N86 ;
  assign n1057 = n1016 & ~n1019 ;
  assign n1058 = N103 & N460 ;
  assign n1059 = n1010 & ~n1013 ;
  assign n1060 = N120 & N443 ;
  assign n1061 = n1004 & ~n1007 ;
  assign n1062 = N137 & N426 ;
  assign n1063 = n998 & ~n1001 ;
  assign n1064 = N154 & N409 ;
  assign n1065 = n992 & ~n995 ;
  assign n1066 = N171 & N392 ;
  assign n1067 = n986 & ~n989 ;
  assign n1068 = N188 & N375 ;
  assign n1069 = n980 & ~n983 ;
  assign n1070 = N205 & N358 ;
  assign n1071 = n974 & ~n977 ;
  assign n1072 = N222 & N341 ;
  assign n1073 = n968 & ~n971 ;
  assign n1074 = N239 & N324 ;
  assign n1075 = N256 & N307 ;
  assign n1076 = n962 & ~n965 ;
  assign n1077 = n1075 | n1076 ;
  assign n1078 = n1075 & n1076 ;
  assign n1079 = n1077 & ~n1078 ;
  assign n1080 = ~n1074 & n1079 ;
  assign n1081 = n1074 & ~n1079 ;
  assign n1082 = n1080 | n1081 ;
  assign n1083 = n1073 | n1082 ;
  assign n1084 = n1073 & n1082 ;
  assign n1085 = n1083 & ~n1084 ;
  assign n1086 = ~n1072 & n1085 ;
  assign n1087 = n1072 & ~n1085 ;
  assign n1088 = n1086 | n1087 ;
  assign n1089 = n1071 | n1088 ;
  assign n1090 = n1071 & n1088 ;
  assign n1091 = n1089 & ~n1090 ;
  assign n1092 = ~n1070 & n1091 ;
  assign n1093 = n1070 & ~n1091 ;
  assign n1094 = n1092 | n1093 ;
  assign n1095 = n1069 | n1094 ;
  assign n1096 = n1069 & n1094 ;
  assign n1097 = n1095 & ~n1096 ;
  assign n1098 = ~n1068 & n1097 ;
  assign n1099 = n1068 & ~n1097 ;
  assign n1100 = n1098 | n1099 ;
  assign n1101 = n1067 | n1100 ;
  assign n1102 = n1067 & n1100 ;
  assign n1103 = n1101 & ~n1102 ;
  assign n1104 = ~n1066 & n1103 ;
  assign n1105 = n1066 & ~n1103 ;
  assign n1106 = n1104 | n1105 ;
  assign n1107 = n1065 | n1106 ;
  assign n1108 = n1065 & n1106 ;
  assign n1109 = n1107 & ~n1108 ;
  assign n1110 = ~n1064 & n1109 ;
  assign n1111 = n1064 & ~n1109 ;
  assign n1112 = n1110 | n1111 ;
  assign n1113 = n1063 | n1112 ;
  assign n1114 = n1063 & n1112 ;
  assign n1115 = n1113 & ~n1114 ;
  assign n1116 = ~n1062 & n1115 ;
  assign n1117 = n1062 & ~n1115 ;
  assign n1118 = n1116 | n1117 ;
  assign n1119 = n1061 | n1118 ;
  assign n1120 = n1061 & n1118 ;
  assign n1121 = n1119 & ~n1120 ;
  assign n1122 = ~n1060 & n1121 ;
  assign n1123 = n1060 & ~n1121 ;
  assign n1124 = n1122 | n1123 ;
  assign n1125 = n1059 | n1124 ;
  assign n1126 = n1059 & n1124 ;
  assign n1127 = n1125 & ~n1126 ;
  assign n1128 = ~n1058 & n1127 ;
  assign n1129 = n1058 & ~n1127 ;
  assign n1130 = n1128 | n1129 ;
  assign n1131 = n1057 | n1130 ;
  assign n1132 = n1057 & n1130 ;
  assign n1133 = n1131 & ~n1132 ;
  assign n1134 = ~n1056 & n1133 ;
  assign n1135 = n1056 & ~n1133 ;
  assign n1136 = n1134 | n1135 ;
  assign n1137 = n1055 | n1136 ;
  assign n1138 = n1055 & n1136 ;
  assign n1139 = n1137 & ~n1138 ;
  assign n1140 = ~n1054 & n1139 ;
  assign n1141 = n1054 & ~n1139 ;
  assign n1142 = n1140 | n1141 ;
  assign n1143 = n1053 | n1142 ;
  assign n1144 = n1053 & n1142 ;
  assign n1145 = n1143 & ~n1144 ;
  assign n1146 = ~n1052 & n1145 ;
  assign n1147 = n1052 & ~n1145 ;
  assign n1148 = n1146 | n1147 ;
  assign n1149 = n1051 | n1148 ;
  assign n1150 = n1051 & n1148 ;
  assign n1151 = n1149 & ~n1150 ;
  assign n1152 = ~n1050 & n1151 ;
  assign n1153 = n1050 & ~n1151 ;
  assign n1154 = n1152 | n1153 ;
  assign n1155 = n1049 | n1154 ;
  assign n1156 = n1049 & n1154 ;
  assign n1157 = n1155 & ~n1156 ;
  assign n1158 = ~n1046 & n1157 ;
  assign n1159 = n1046 & ~n1157 ;
  assign n1160 = n1158 | n1159 ;
  assign n1161 = n1155 & ~n1158 ;
  assign n1162 = n1149 & ~n1152 ;
  assign n1163 = N52 & N528 ;
  assign n1164 = n1143 & ~n1146 ;
  assign n1165 = N511 & N69 ;
  assign n1166 = n1137 & ~n1140 ;
  assign n1167 = N494 & N86 ;
  assign n1168 = n1131 & ~n1134 ;
  assign n1169 = N103 & N477 ;
  assign n1170 = n1125 & ~n1128 ;
  assign n1171 = N120 & N460 ;
  assign n1172 = n1119 & ~n1122 ;
  assign n1173 = N137 & N443 ;
  assign n1174 = n1113 & ~n1116 ;
  assign n1175 = N154 & N426 ;
  assign n1176 = n1107 & ~n1110 ;
  assign n1177 = N171 & N409 ;
  assign n1178 = n1101 & ~n1104 ;
  assign n1179 = N188 & N392 ;
  assign n1180 = n1095 & ~n1098 ;
  assign n1181 = N205 & N375 ;
  assign n1182 = n1089 & ~n1092 ;
  assign n1183 = N222 & N358 ;
  assign n1184 = n1083 & ~n1086 ;
  assign n1185 = N239 & N341 ;
  assign n1186 = N256 & N324 ;
  assign n1187 = n1077 & ~n1080 ;
  assign n1188 = n1186 | n1187 ;
  assign n1189 = n1186 & n1187 ;
  assign n1190 = n1188 & ~n1189 ;
  assign n1191 = ~n1185 & n1190 ;
  assign n1192 = n1185 & ~n1190 ;
  assign n1193 = n1191 | n1192 ;
  assign n1194 = n1184 | n1193 ;
  assign n1195 = n1184 & n1193 ;
  assign n1196 = n1194 & ~n1195 ;
  assign n1197 = ~n1183 & n1196 ;
  assign n1198 = n1183 & ~n1196 ;
  assign n1199 = n1197 | n1198 ;
  assign n1200 = n1182 | n1199 ;
  assign n1201 = n1182 & n1199 ;
  assign n1202 = n1200 & ~n1201 ;
  assign n1203 = ~n1181 & n1202 ;
  assign n1204 = n1181 & ~n1202 ;
  assign n1205 = n1203 | n1204 ;
  assign n1206 = n1180 | n1205 ;
  assign n1207 = n1180 & n1205 ;
  assign n1208 = n1206 & ~n1207 ;
  assign n1209 = ~n1179 & n1208 ;
  assign n1210 = n1179 & ~n1208 ;
  assign n1211 = n1209 | n1210 ;
  assign n1212 = n1178 | n1211 ;
  assign n1213 = n1178 & n1211 ;
  assign n1214 = n1212 & ~n1213 ;
  assign n1215 = ~n1177 & n1214 ;
  assign n1216 = n1177 & ~n1214 ;
  assign n1217 = n1215 | n1216 ;
  assign n1218 = n1176 | n1217 ;
  assign n1219 = n1176 & n1217 ;
  assign n1220 = n1218 & ~n1219 ;
  assign n1221 = ~n1175 & n1220 ;
  assign n1222 = n1175 & ~n1220 ;
  assign n1223 = n1221 | n1222 ;
  assign n1224 = n1174 | n1223 ;
  assign n1225 = n1174 & n1223 ;
  assign n1226 = n1224 & ~n1225 ;
  assign n1227 = ~n1173 & n1226 ;
  assign n1228 = n1173 & ~n1226 ;
  assign n1229 = n1227 | n1228 ;
  assign n1230 = n1172 | n1229 ;
  assign n1231 = n1172 & n1229 ;
  assign n1232 = n1230 & ~n1231 ;
  assign n1233 = ~n1171 & n1232 ;
  assign n1234 = n1171 & ~n1232 ;
  assign n1235 = n1233 | n1234 ;
  assign n1236 = n1170 | n1235 ;
  assign n1237 = n1170 & n1235 ;
  assign n1238 = n1236 & ~n1237 ;
  assign n1239 = ~n1169 & n1238 ;
  assign n1240 = n1169 & ~n1238 ;
  assign n1241 = n1239 | n1240 ;
  assign n1242 = n1168 | n1241 ;
  assign n1243 = n1168 & n1241 ;
  assign n1244 = n1242 & ~n1243 ;
  assign n1245 = ~n1167 & n1244 ;
  assign n1246 = n1167 & ~n1244 ;
  assign n1247 = n1245 | n1246 ;
  assign n1248 = n1166 | n1247 ;
  assign n1249 = n1166 & n1247 ;
  assign n1250 = n1248 & ~n1249 ;
  assign n1251 = ~n1165 & n1250 ;
  assign n1252 = n1165 & ~n1250 ;
  assign n1253 = n1251 | n1252 ;
  assign n1254 = n1164 | n1253 ;
  assign n1255 = n1164 & n1253 ;
  assign n1256 = n1254 & ~n1255 ;
  assign n1257 = ~n1163 & n1256 ;
  assign n1258 = n1163 & ~n1256 ;
  assign n1259 = n1257 | n1258 ;
  assign n1260 = n1162 | n1259 ;
  assign n1261 = n1162 & n1259 ;
  assign n1262 = n1260 & ~n1261 ;
  assign n1263 = ~n1161 & n1262 ;
  assign n1264 = n1161 & ~n1262 ;
  assign n1265 = n1263 | n1264 ;
  assign n1266 = n1260 & ~n1263 ;
  assign n1267 = n1254 & ~n1257 ;
  assign n1268 = N528 & N69 ;
  assign n1269 = n1248 & ~n1251 ;
  assign n1270 = N511 & N86 ;
  assign n1271 = n1242 & ~n1245 ;
  assign n1272 = N103 & N494 ;
  assign n1273 = n1236 & ~n1239 ;
  assign n1274 = N120 & N477 ;
  assign n1275 = n1230 & ~n1233 ;
  assign n1276 = N137 & N460 ;
  assign n1277 = n1224 & ~n1227 ;
  assign n1278 = N154 & N443 ;
  assign n1279 = n1218 & ~n1221 ;
  assign n1280 = N171 & N426 ;
  assign n1281 = n1212 & ~n1215 ;
  assign n1282 = N188 & N409 ;
  assign n1283 = n1206 & ~n1209 ;
  assign n1284 = N205 & N392 ;
  assign n1285 = n1200 & ~n1203 ;
  assign n1286 = N222 & N375 ;
  assign n1287 = n1194 & ~n1197 ;
  assign n1288 = N239 & N358 ;
  assign n1289 = N256 & N341 ;
  assign n1290 = n1188 & ~n1191 ;
  assign n1291 = n1289 | n1290 ;
  assign n1292 = n1289 & n1290 ;
  assign n1293 = n1291 & ~n1292 ;
  assign n1294 = ~n1288 & n1293 ;
  assign n1295 = n1288 & ~n1293 ;
  assign n1296 = n1294 | n1295 ;
  assign n1297 = n1287 | n1296 ;
  assign n1298 = n1287 & n1296 ;
  assign n1299 = n1297 & ~n1298 ;
  assign n1300 = ~n1286 & n1299 ;
  assign n1301 = n1286 & ~n1299 ;
  assign n1302 = n1300 | n1301 ;
  assign n1303 = n1285 | n1302 ;
  assign n1304 = n1285 & n1302 ;
  assign n1305 = n1303 & ~n1304 ;
  assign n1306 = ~n1284 & n1305 ;
  assign n1307 = n1284 & ~n1305 ;
  assign n1308 = n1306 | n1307 ;
  assign n1309 = n1283 | n1308 ;
  assign n1310 = n1283 & n1308 ;
  assign n1311 = n1309 & ~n1310 ;
  assign n1312 = ~n1282 & n1311 ;
  assign n1313 = n1282 & ~n1311 ;
  assign n1314 = n1312 | n1313 ;
  assign n1315 = n1281 | n1314 ;
  assign n1316 = n1281 & n1314 ;
  assign n1317 = n1315 & ~n1316 ;
  assign n1318 = ~n1280 & n1317 ;
  assign n1319 = n1280 & ~n1317 ;
  assign n1320 = n1318 | n1319 ;
  assign n1321 = n1279 | n1320 ;
  assign n1322 = n1279 & n1320 ;
  assign n1323 = n1321 & ~n1322 ;
  assign n1324 = ~n1278 & n1323 ;
  assign n1325 = n1278 & ~n1323 ;
  assign n1326 = n1324 | n1325 ;
  assign n1327 = n1277 | n1326 ;
  assign n1328 = n1277 & n1326 ;
  assign n1329 = n1327 & ~n1328 ;
  assign n1330 = ~n1276 & n1329 ;
  assign n1331 = n1276 & ~n1329 ;
  assign n1332 = n1330 | n1331 ;
  assign n1333 = n1275 | n1332 ;
  assign n1334 = n1275 & n1332 ;
  assign n1335 = n1333 & ~n1334 ;
  assign n1336 = ~n1274 & n1335 ;
  assign n1337 = n1274 & ~n1335 ;
  assign n1338 = n1336 | n1337 ;
  assign n1339 = n1273 | n1338 ;
  assign n1340 = n1273 & n1338 ;
  assign n1341 = n1339 & ~n1340 ;
  assign n1342 = ~n1272 & n1341 ;
  assign n1343 = n1272 & ~n1341 ;
  assign n1344 = n1342 | n1343 ;
  assign n1345 = n1271 | n1344 ;
  assign n1346 = n1271 & n1344 ;
  assign n1347 = n1345 & ~n1346 ;
  assign n1348 = ~n1270 & n1347 ;
  assign n1349 = n1270 & ~n1347 ;
  assign n1350 = n1348 | n1349 ;
  assign n1351 = n1269 | n1350 ;
  assign n1352 = n1269 & n1350 ;
  assign n1353 = n1351 & ~n1352 ;
  assign n1354 = ~n1268 & n1353 ;
  assign n1355 = n1268 & ~n1353 ;
  assign n1356 = n1354 | n1355 ;
  assign n1357 = n1267 | n1356 ;
  assign n1358 = n1267 & n1356 ;
  assign n1359 = n1357 & ~n1358 ;
  assign n1360 = ~n1266 & n1359 ;
  assign n1361 = n1266 & ~n1359 ;
  assign n1362 = n1360 | n1361 ;
  assign n1363 = n1357 & ~n1360 ;
  assign n1364 = n1351 & ~n1354 ;
  assign n1365 = N528 & N86 ;
  assign n1366 = n1345 & ~n1348 ;
  assign n1367 = N103 & N511 ;
  assign n1368 = n1339 & ~n1342 ;
  assign n1369 = N120 & N494 ;
  assign n1370 = n1333 & ~n1336 ;
  assign n1371 = N137 & N477 ;
  assign n1372 = n1327 & ~n1330 ;
  assign n1373 = N154 & N460 ;
  assign n1374 = n1321 & ~n1324 ;
  assign n1375 = N171 & N443 ;
  assign n1376 = n1315 & ~n1318 ;
  assign n1377 = N188 & N426 ;
  assign n1378 = n1309 & ~n1312 ;
  assign n1379 = N205 & N409 ;
  assign n1380 = n1303 & ~n1306 ;
  assign n1381 = N222 & N392 ;
  assign n1382 = n1297 & ~n1300 ;
  assign n1383 = N239 & N375 ;
  assign n1384 = N256 & N358 ;
  assign n1385 = n1291 & ~n1294 ;
  assign n1386 = n1384 | n1385 ;
  assign n1387 = n1384 & n1385 ;
  assign n1388 = n1386 & ~n1387 ;
  assign n1389 = ~n1383 & n1388 ;
  assign n1390 = n1383 & ~n1388 ;
  assign n1391 = n1389 | n1390 ;
  assign n1392 = n1382 | n1391 ;
  assign n1393 = n1382 & n1391 ;
  assign n1394 = n1392 & ~n1393 ;
  assign n1395 = ~n1381 & n1394 ;
  assign n1396 = n1381 & ~n1394 ;
  assign n1397 = n1395 | n1396 ;
  assign n1398 = n1380 | n1397 ;
  assign n1399 = n1380 & n1397 ;
  assign n1400 = n1398 & ~n1399 ;
  assign n1401 = ~n1379 & n1400 ;
  assign n1402 = n1379 & ~n1400 ;
  assign n1403 = n1401 | n1402 ;
  assign n1404 = n1378 | n1403 ;
  assign n1405 = n1378 & n1403 ;
  assign n1406 = n1404 & ~n1405 ;
  assign n1407 = ~n1377 & n1406 ;
  assign n1408 = n1377 & ~n1406 ;
  assign n1409 = n1407 | n1408 ;
  assign n1410 = n1376 | n1409 ;
  assign n1411 = n1376 & n1409 ;
  assign n1412 = n1410 & ~n1411 ;
  assign n1413 = ~n1375 & n1412 ;
  assign n1414 = n1375 & ~n1412 ;
  assign n1415 = n1413 | n1414 ;
  assign n1416 = n1374 | n1415 ;
  assign n1417 = n1374 & n1415 ;
  assign n1418 = n1416 & ~n1417 ;
  assign n1419 = ~n1373 & n1418 ;
  assign n1420 = n1373 & ~n1418 ;
  assign n1421 = n1419 | n1420 ;
  assign n1422 = n1372 | n1421 ;
  assign n1423 = n1372 & n1421 ;
  assign n1424 = n1422 & ~n1423 ;
  assign n1425 = ~n1371 & n1424 ;
  assign n1426 = n1371 & ~n1424 ;
  assign n1427 = n1425 | n1426 ;
  assign n1428 = n1370 | n1427 ;
  assign n1429 = n1370 & n1427 ;
  assign n1430 = n1428 & ~n1429 ;
  assign n1431 = ~n1369 & n1430 ;
  assign n1432 = n1369 & ~n1430 ;
  assign n1433 = n1431 | n1432 ;
  assign n1434 = n1368 | n1433 ;
  assign n1435 = n1368 & n1433 ;
  assign n1436 = n1434 & ~n1435 ;
  assign n1437 = ~n1367 & n1436 ;
  assign n1438 = n1367 & ~n1436 ;
  assign n1439 = n1437 | n1438 ;
  assign n1440 = n1366 | n1439 ;
  assign n1441 = n1366 & n1439 ;
  assign n1442 = n1440 & ~n1441 ;
  assign n1443 = ~n1365 & n1442 ;
  assign n1444 = n1365 & ~n1442 ;
  assign n1445 = n1443 | n1444 ;
  assign n1446 = n1364 | n1445 ;
  assign n1447 = n1364 & n1445 ;
  assign n1448 = n1446 & ~n1447 ;
  assign n1449 = ~n1363 & n1448 ;
  assign n1450 = n1363 & ~n1448 ;
  assign n1451 = n1449 | n1450 ;
  assign n1452 = n1446 & ~n1449 ;
  assign n1453 = n1440 & ~n1443 ;
  assign n1454 = N103 & N528 ;
  assign n1455 = n1434 & ~n1437 ;
  assign n1456 = N120 & N511 ;
  assign n1457 = n1428 & ~n1431 ;
  assign n1458 = N137 & N494 ;
  assign n1459 = n1422 & ~n1425 ;
  assign n1460 = N154 & N477 ;
  assign n1461 = n1416 & ~n1419 ;
  assign n1462 = N171 & N460 ;
  assign n1463 = n1410 & ~n1413 ;
  assign n1464 = N188 & N443 ;
  assign n1465 = n1404 & ~n1407 ;
  assign n1466 = N205 & N426 ;
  assign n1467 = n1398 & ~n1401 ;
  assign n1468 = N222 & N409 ;
  assign n1469 = n1392 & ~n1395 ;
  assign n1470 = N239 & N392 ;
  assign n1471 = N256 & N375 ;
  assign n1472 = n1386 & ~n1389 ;
  assign n1473 = n1471 | n1472 ;
  assign n1474 = n1471 & n1472 ;
  assign n1475 = n1473 & ~n1474 ;
  assign n1476 = ~n1470 & n1475 ;
  assign n1477 = n1470 & ~n1475 ;
  assign n1478 = n1476 | n1477 ;
  assign n1479 = n1469 | n1478 ;
  assign n1480 = n1469 & n1478 ;
  assign n1481 = n1479 & ~n1480 ;
  assign n1482 = ~n1468 & n1481 ;
  assign n1483 = n1468 & ~n1481 ;
  assign n1484 = n1482 | n1483 ;
  assign n1485 = n1467 | n1484 ;
  assign n1486 = n1467 & n1484 ;
  assign n1487 = n1485 & ~n1486 ;
  assign n1488 = ~n1466 & n1487 ;
  assign n1489 = n1466 & ~n1487 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = n1465 | n1490 ;
  assign n1492 = n1465 & n1490 ;
  assign n1493 = n1491 & ~n1492 ;
  assign n1494 = ~n1464 & n1493 ;
  assign n1495 = n1464 & ~n1493 ;
  assign n1496 = n1494 | n1495 ;
  assign n1497 = n1463 | n1496 ;
  assign n1498 = n1463 & n1496 ;
  assign n1499 = n1497 & ~n1498 ;
  assign n1500 = ~n1462 & n1499 ;
  assign n1501 = n1462 & ~n1499 ;
  assign n1502 = n1500 | n1501 ;
  assign n1503 = n1461 | n1502 ;
  assign n1504 = n1461 & n1502 ;
  assign n1505 = n1503 & ~n1504 ;
  assign n1506 = ~n1460 & n1505 ;
  assign n1507 = n1460 & ~n1505 ;
  assign n1508 = n1506 | n1507 ;
  assign n1509 = n1459 | n1508 ;
  assign n1510 = n1459 & n1508 ;
  assign n1511 = n1509 & ~n1510 ;
  assign n1512 = ~n1458 & n1511 ;
  assign n1513 = n1458 & ~n1511 ;
  assign n1514 = n1512 | n1513 ;
  assign n1515 = n1457 | n1514 ;
  assign n1516 = n1457 & n1514 ;
  assign n1517 = n1515 & ~n1516 ;
  assign n1518 = ~n1456 & n1517 ;
  assign n1519 = n1456 & ~n1517 ;
  assign n1520 = n1518 | n1519 ;
  assign n1521 = n1455 | n1520 ;
  assign n1522 = n1455 & n1520 ;
  assign n1523 = n1521 & ~n1522 ;
  assign n1524 = ~n1454 & n1523 ;
  assign n1525 = n1454 & ~n1523 ;
  assign n1526 = n1524 | n1525 ;
  assign n1527 = n1453 | n1526 ;
  assign n1528 = n1453 & n1526 ;
  assign n1529 = n1527 & ~n1528 ;
  assign n1530 = ~n1452 & n1529 ;
  assign n1531 = n1452 & ~n1529 ;
  assign n1532 = n1530 | n1531 ;
  assign n1533 = n1527 & ~n1530 ;
  assign n1534 = n1521 & ~n1524 ;
  assign n1535 = N120 & N528 ;
  assign n1536 = n1515 & ~n1518 ;
  assign n1537 = N137 & N511 ;
  assign n1538 = n1509 & ~n1512 ;
  assign n1539 = N154 & N494 ;
  assign n1540 = n1503 & ~n1506 ;
  assign n1541 = N171 & N477 ;
  assign n1542 = n1497 & ~n1500 ;
  assign n1543 = N188 & N460 ;
  assign n1544 = n1491 & ~n1494 ;
  assign n1545 = N205 & N443 ;
  assign n1546 = n1485 & ~n1488 ;
  assign n1547 = N222 & N426 ;
  assign n1548 = n1479 & ~n1482 ;
  assign n1549 = N239 & N409 ;
  assign n1550 = N256 & N392 ;
  assign n1551 = n1473 & ~n1476 ;
  assign n1552 = n1550 | n1551 ;
  assign n1553 = n1550 & n1551 ;
  assign n1554 = n1552 & ~n1553 ;
  assign n1555 = ~n1549 & n1554 ;
  assign n1556 = n1549 & ~n1554 ;
  assign n1557 = n1555 | n1556 ;
  assign n1558 = n1548 | n1557 ;
  assign n1559 = n1548 & n1557 ;
  assign n1560 = n1558 & ~n1559 ;
  assign n1561 = ~n1547 & n1560 ;
  assign n1562 = n1547 & ~n1560 ;
  assign n1563 = n1561 | n1562 ;
  assign n1564 = n1546 | n1563 ;
  assign n1565 = n1546 & n1563 ;
  assign n1566 = n1564 & ~n1565 ;
  assign n1567 = ~n1545 & n1566 ;
  assign n1568 = n1545 & ~n1566 ;
  assign n1569 = n1567 | n1568 ;
  assign n1570 = n1544 | n1569 ;
  assign n1571 = n1544 & n1569 ;
  assign n1572 = n1570 & ~n1571 ;
  assign n1573 = ~n1543 & n1572 ;
  assign n1574 = n1543 & ~n1572 ;
  assign n1575 = n1573 | n1574 ;
  assign n1576 = n1542 | n1575 ;
  assign n1577 = n1542 & n1575 ;
  assign n1578 = n1576 & ~n1577 ;
  assign n1579 = ~n1541 & n1578 ;
  assign n1580 = n1541 & ~n1578 ;
  assign n1581 = n1579 | n1580 ;
  assign n1582 = n1540 | n1581 ;
  assign n1583 = n1540 & n1581 ;
  assign n1584 = n1582 & ~n1583 ;
  assign n1585 = ~n1539 & n1584 ;
  assign n1586 = n1539 & ~n1584 ;
  assign n1587 = n1585 | n1586 ;
  assign n1588 = n1538 | n1587 ;
  assign n1589 = n1538 & n1587 ;
  assign n1590 = n1588 & ~n1589 ;
  assign n1591 = ~n1537 & n1590 ;
  assign n1592 = n1537 & ~n1590 ;
  assign n1593 = n1591 | n1592 ;
  assign n1594 = n1536 | n1593 ;
  assign n1595 = n1536 & n1593 ;
  assign n1596 = n1594 & ~n1595 ;
  assign n1597 = ~n1535 & n1596 ;
  assign n1598 = n1535 & ~n1596 ;
  assign n1599 = n1597 | n1598 ;
  assign n1600 = n1534 | n1599 ;
  assign n1601 = n1534 & n1599 ;
  assign n1602 = n1600 & ~n1601 ;
  assign n1603 = ~n1533 & n1602 ;
  assign n1604 = n1533 & ~n1602 ;
  assign n1605 = n1603 | n1604 ;
  assign n1606 = n1600 & ~n1603 ;
  assign n1607 = n1594 & ~n1597 ;
  assign n1608 = N137 & N528 ;
  assign n1609 = n1588 & ~n1591 ;
  assign n1610 = N154 & N511 ;
  assign n1611 = n1582 & ~n1585 ;
  assign n1612 = N171 & N494 ;
  assign n1613 = n1576 & ~n1579 ;
  assign n1614 = N188 & N477 ;
  assign n1615 = n1570 & ~n1573 ;
  assign n1616 = N205 & N460 ;
  assign n1617 = n1564 & ~n1567 ;
  assign n1618 = N222 & N443 ;
  assign n1619 = n1558 & ~n1561 ;
  assign n1620 = N239 & N426 ;
  assign n1621 = N256 & N409 ;
  assign n1622 = n1552 & ~n1555 ;
  assign n1623 = n1621 | n1622 ;
  assign n1624 = n1621 & n1622 ;
  assign n1625 = n1623 & ~n1624 ;
  assign n1626 = ~n1620 & n1625 ;
  assign n1627 = n1620 & ~n1625 ;
  assign n1628 = n1626 | n1627 ;
  assign n1629 = n1619 | n1628 ;
  assign n1630 = n1619 & n1628 ;
  assign n1631 = n1629 & ~n1630 ;
  assign n1632 = ~n1618 & n1631 ;
  assign n1633 = n1618 & ~n1631 ;
  assign n1634 = n1632 | n1633 ;
  assign n1635 = n1617 | n1634 ;
  assign n1636 = n1617 & n1634 ;
  assign n1637 = n1635 & ~n1636 ;
  assign n1638 = ~n1616 & n1637 ;
  assign n1639 = n1616 & ~n1637 ;
  assign n1640 = n1638 | n1639 ;
  assign n1641 = n1615 | n1640 ;
  assign n1642 = n1615 & n1640 ;
  assign n1643 = n1641 & ~n1642 ;
  assign n1644 = ~n1614 & n1643 ;
  assign n1645 = n1614 & ~n1643 ;
  assign n1646 = n1644 | n1645 ;
  assign n1647 = n1613 | n1646 ;
  assign n1648 = n1613 & n1646 ;
  assign n1649 = n1647 & ~n1648 ;
  assign n1650 = ~n1612 & n1649 ;
  assign n1651 = n1612 & ~n1649 ;
  assign n1652 = n1650 | n1651 ;
  assign n1653 = n1611 | n1652 ;
  assign n1654 = n1611 & n1652 ;
  assign n1655 = n1653 & ~n1654 ;
  assign n1656 = ~n1610 & n1655 ;
  assign n1657 = n1610 & ~n1655 ;
  assign n1658 = n1656 | n1657 ;
  assign n1659 = n1609 | n1658 ;
  assign n1660 = n1609 & n1658 ;
  assign n1661 = n1659 & ~n1660 ;
  assign n1662 = ~n1608 & n1661 ;
  assign n1663 = n1608 & ~n1661 ;
  assign n1664 = n1662 | n1663 ;
  assign n1665 = n1607 | n1664 ;
  assign n1666 = n1607 & n1664 ;
  assign n1667 = n1665 & ~n1666 ;
  assign n1668 = ~n1606 & n1667 ;
  assign n1669 = n1606 & ~n1667 ;
  assign n1670 = n1668 | n1669 ;
  assign n1671 = n1665 & ~n1668 ;
  assign n1672 = n1659 & ~n1662 ;
  assign n1673 = N154 & N528 ;
  assign n1674 = n1653 & ~n1656 ;
  assign n1675 = N171 & N511 ;
  assign n1676 = n1647 & ~n1650 ;
  assign n1677 = N188 & N494 ;
  assign n1678 = n1641 & ~n1644 ;
  assign n1679 = N205 & N477 ;
  assign n1680 = n1635 & ~n1638 ;
  assign n1681 = N222 & N460 ;
  assign n1682 = n1629 & ~n1632 ;
  assign n1683 = N239 & N443 ;
  assign n1684 = N256 & N426 ;
  assign n1685 = n1623 & ~n1626 ;
  assign n1686 = n1684 | n1685 ;
  assign n1687 = n1684 & n1685 ;
  assign n1688 = n1686 & ~n1687 ;
  assign n1689 = ~n1683 & n1688 ;
  assign n1690 = n1683 & ~n1688 ;
  assign n1691 = n1689 | n1690 ;
  assign n1692 = n1682 | n1691 ;
  assign n1693 = n1682 & n1691 ;
  assign n1694 = n1692 & ~n1693 ;
  assign n1695 = ~n1681 & n1694 ;
  assign n1696 = n1681 & ~n1694 ;
  assign n1697 = n1695 | n1696 ;
  assign n1698 = n1680 | n1697 ;
  assign n1699 = n1680 & n1697 ;
  assign n1700 = n1698 & ~n1699 ;
  assign n1701 = ~n1679 & n1700 ;
  assign n1702 = n1679 & ~n1700 ;
  assign n1703 = n1701 | n1702 ;
  assign n1704 = n1678 | n1703 ;
  assign n1705 = n1678 & n1703 ;
  assign n1706 = n1704 & ~n1705 ;
  assign n1707 = ~n1677 & n1706 ;
  assign n1708 = n1677 & ~n1706 ;
  assign n1709 = n1707 | n1708 ;
  assign n1710 = n1676 | n1709 ;
  assign n1711 = n1676 & n1709 ;
  assign n1712 = n1710 & ~n1711 ;
  assign n1713 = ~n1675 & n1712 ;
  assign n1714 = n1675 & ~n1712 ;
  assign n1715 = n1713 | n1714 ;
  assign n1716 = n1674 | n1715 ;
  assign n1717 = n1674 & n1715 ;
  assign n1718 = n1716 & ~n1717 ;
  assign n1719 = ~n1673 & n1718 ;
  assign n1720 = n1673 & ~n1718 ;
  assign n1721 = n1719 | n1720 ;
  assign n1722 = n1672 | n1721 ;
  assign n1723 = n1672 & n1721 ;
  assign n1724 = n1722 & ~n1723 ;
  assign n1725 = ~n1671 & n1724 ;
  assign n1726 = n1671 & ~n1724 ;
  assign n1727 = n1725 | n1726 ;
  assign n1728 = n1722 & ~n1725 ;
  assign n1729 = n1716 & ~n1719 ;
  assign n1730 = N171 & N528 ;
  assign n1731 = n1710 & ~n1713 ;
  assign n1732 = N188 & N511 ;
  assign n1733 = n1704 & ~n1707 ;
  assign n1734 = N205 & N494 ;
  assign n1735 = n1698 & ~n1701 ;
  assign n1736 = N222 & N477 ;
  assign n1737 = n1692 & ~n1695 ;
  assign n1738 = N239 & N460 ;
  assign n1739 = N256 & N443 ;
  assign n1740 = n1686 & ~n1689 ;
  assign n1741 = n1739 | n1740 ;
  assign n1742 = n1739 & n1740 ;
  assign n1743 = n1741 & ~n1742 ;
  assign n1744 = ~n1738 & n1743 ;
  assign n1745 = n1738 & ~n1743 ;
  assign n1746 = n1744 | n1745 ;
  assign n1747 = n1737 | n1746 ;
  assign n1748 = n1737 & n1746 ;
  assign n1749 = n1747 & ~n1748 ;
  assign n1750 = ~n1736 & n1749 ;
  assign n1751 = n1736 & ~n1749 ;
  assign n1752 = n1750 | n1751 ;
  assign n1753 = n1735 | n1752 ;
  assign n1754 = n1735 & n1752 ;
  assign n1755 = n1753 & ~n1754 ;
  assign n1756 = ~n1734 & n1755 ;
  assign n1757 = n1734 & ~n1755 ;
  assign n1758 = n1756 | n1757 ;
  assign n1759 = n1733 | n1758 ;
  assign n1760 = n1733 & n1758 ;
  assign n1761 = n1759 & ~n1760 ;
  assign n1762 = ~n1732 & n1761 ;
  assign n1763 = n1732 & ~n1761 ;
  assign n1764 = n1762 | n1763 ;
  assign n1765 = n1731 | n1764 ;
  assign n1766 = n1731 & n1764 ;
  assign n1767 = n1765 & ~n1766 ;
  assign n1768 = ~n1730 & n1767 ;
  assign n1769 = n1730 & ~n1767 ;
  assign n1770 = n1768 | n1769 ;
  assign n1771 = n1729 | n1770 ;
  assign n1772 = n1729 & n1770 ;
  assign n1773 = n1771 & ~n1772 ;
  assign n1774 = ~n1728 & n1773 ;
  assign n1775 = n1728 & ~n1773 ;
  assign n1776 = n1774 | n1775 ;
  assign n1777 = n1771 & ~n1774 ;
  assign n1778 = n1765 & ~n1768 ;
  assign n1779 = N188 & N528 ;
  assign n1780 = n1759 & ~n1762 ;
  assign n1781 = N205 & N511 ;
  assign n1782 = n1753 & ~n1756 ;
  assign n1783 = N222 & N494 ;
  assign n1784 = n1747 & ~n1750 ;
  assign n1785 = N239 & N477 ;
  assign n1786 = N256 & N460 ;
  assign n1787 = n1741 & ~n1744 ;
  assign n1788 = n1786 | n1787 ;
  assign n1789 = n1786 & n1787 ;
  assign n1790 = n1788 & ~n1789 ;
  assign n1791 = ~n1785 & n1790 ;
  assign n1792 = n1785 & ~n1790 ;
  assign n1793 = n1791 | n1792 ;
  assign n1794 = n1784 | n1793 ;
  assign n1795 = n1784 & n1793 ;
  assign n1796 = n1794 & ~n1795 ;
  assign n1797 = ~n1783 & n1796 ;
  assign n1798 = n1783 & ~n1796 ;
  assign n1799 = n1797 | n1798 ;
  assign n1800 = n1782 | n1799 ;
  assign n1801 = n1782 & n1799 ;
  assign n1802 = n1800 & ~n1801 ;
  assign n1803 = ~n1781 & n1802 ;
  assign n1804 = n1781 & ~n1802 ;
  assign n1805 = n1803 | n1804 ;
  assign n1806 = n1780 | n1805 ;
  assign n1807 = n1780 & n1805 ;
  assign n1808 = n1806 & ~n1807 ;
  assign n1809 = ~n1779 & n1808 ;
  assign n1810 = n1779 & ~n1808 ;
  assign n1811 = n1809 | n1810 ;
  assign n1812 = n1778 | n1811 ;
  assign n1813 = n1778 & n1811 ;
  assign n1814 = n1812 & ~n1813 ;
  assign n1815 = ~n1777 & n1814 ;
  assign n1816 = n1777 & ~n1814 ;
  assign n1817 = n1815 | n1816 ;
  assign n1818 = n1812 & ~n1815 ;
  assign n1819 = n1806 & ~n1809 ;
  assign n1820 = N205 & N528 ;
  assign n1821 = n1800 & ~n1803 ;
  assign n1822 = N222 & N511 ;
  assign n1823 = n1794 & ~n1797 ;
  assign n1824 = N239 & N494 ;
  assign n1825 = N256 & N477 ;
  assign n1826 = n1788 & ~n1791 ;
  assign n1827 = n1825 | n1826 ;
  assign n1828 = n1825 & n1826 ;
  assign n1829 = n1827 & ~n1828 ;
  assign n1830 = ~n1824 & n1829 ;
  assign n1831 = n1824 & ~n1829 ;
  assign n1832 = n1830 | n1831 ;
  assign n1833 = n1823 | n1832 ;
  assign n1834 = n1823 & n1832 ;
  assign n1835 = n1833 & ~n1834 ;
  assign n1836 = ~n1822 & n1835 ;
  assign n1837 = n1822 & ~n1835 ;
  assign n1838 = n1836 | n1837 ;
  assign n1839 = n1821 | n1838 ;
  assign n1840 = n1821 & n1838 ;
  assign n1841 = n1839 & ~n1840 ;
  assign n1842 = ~n1820 & n1841 ;
  assign n1843 = n1820 & ~n1841 ;
  assign n1844 = n1842 | n1843 ;
  assign n1845 = n1819 | n1844 ;
  assign n1846 = n1819 & n1844 ;
  assign n1847 = n1845 & ~n1846 ;
  assign n1848 = ~n1818 & n1847 ;
  assign n1849 = n1818 & ~n1847 ;
  assign n1850 = n1848 | n1849 ;
  assign n1851 = n1845 & ~n1848 ;
  assign n1852 = n1839 & ~n1842 ;
  assign n1853 = N222 & N528 ;
  assign n1854 = n1833 & ~n1836 ;
  assign n1855 = N239 & N511 ;
  assign n1856 = N256 & N494 ;
  assign n1857 = n1827 & ~n1830 ;
  assign n1858 = n1856 | n1857 ;
  assign n1859 = n1856 & n1857 ;
  assign n1860 = n1858 & ~n1859 ;
  assign n1861 = ~n1855 & n1860 ;
  assign n1862 = n1855 & ~n1860 ;
  assign n1863 = n1861 | n1862 ;
  assign n1864 = n1854 | n1863 ;
  assign n1865 = n1854 & n1863 ;
  assign n1866 = n1864 & ~n1865 ;
  assign n1867 = ~n1853 & n1866 ;
  assign n1868 = n1853 & ~n1866 ;
  assign n1869 = n1867 | n1868 ;
  assign n1870 = n1852 | n1869 ;
  assign n1871 = n1852 & n1869 ;
  assign n1872 = n1870 & ~n1871 ;
  assign n1873 = ~n1851 & n1872 ;
  assign n1874 = n1851 & ~n1872 ;
  assign n1875 = n1873 | n1874 ;
  assign n1876 = n1870 & ~n1873 ;
  assign n1877 = n1864 & ~n1867 ;
  assign n1878 = N239 & N528 ;
  assign n1879 = N256 & N511 ;
  assign n1880 = n1858 & ~n1861 ;
  assign n1881 = n1879 | n1880 ;
  assign n1882 = n1879 & n1880 ;
  assign n1883 = n1881 & ~n1882 ;
  assign n1884 = ~n1878 & n1883 ;
  assign n1885 = n1878 & ~n1883 ;
  assign n1886 = n1884 | n1885 ;
  assign n1887 = n1877 | n1886 ;
  assign n1888 = n1877 & n1886 ;
  assign n1889 = n1887 & ~n1888 ;
  assign n1890 = ~n1876 & n1889 ;
  assign n1891 = n1876 & ~n1889 ;
  assign n1892 = n1890 | n1891 ;
  assign n1893 = N256 & N528 ;
  assign n1894 = n1881 & ~n1884 ;
  assign n1895 = n1893 | n1894 ;
  assign n1896 = n1887 & ~n1890 ;
  assign n1897 = n1893 & n1894 ;
  assign n1898 = n1895 & ~n1897 ;
  assign n1899 = ~n1896 & n1898 ;
  assign n1900 = n1895 & ~n1899 ;
  assign n1901 = n1896 & ~n1898 ;
  assign n1902 = n1899 | n1901 ;
  assign N1581 = n39 ;
  assign N1901 = n51 ;
  assign N2223 = n71 ;
  assign N2548 = n99 ;
  assign N2877 = n135 ;
  assign N3211 = n179 ;
  assign N3552 = n231 ;
  assign N3895 = n291 ;
  assign N4241 = n359 ;
  assign N4591 = n435 ;
  assign N4946 = n519 ;
  assign N5308 = n611 ;
  assign N545 = n34 ;
  assign N5672 = n711 ;
  assign N5971 = n819 ;
  assign N6123 = n934 ;
  assign N6150 = n1048 ;
  assign N6160 = n1160 ;
  assign N6170 = n1265 ;
  assign N6180 = n1362 ;
  assign N6190 = n1451 ;
  assign N6200 = n1532 ;
  assign N6210 = n1605 ;
  assign N6220 = n1670 ;
  assign N6230 = n1727 ;
  assign N6240 = n1776 ;
  assign N6250 = n1817 ;
  assign N6260 = n1850 ;
  assign N6270 = n1875 ;
  assign N6280 = n1892 ;
  assign N6287 = n1900 ;
  assign N6288 = n1902 ;
endmodule
