module top( x0 , x1 , x2 , x3 , x4 , x5 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 );
  input x0 , x1 , x2 , x3 , x4 , x5 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 ;
  wire n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 ;
  assign n7 = ( x1 & x2 ) | ( x1 & x3 ) | ( x2 & x3 ) ;
  assign n8 = x4 & ~n7 ;
  assign n9 = ( x1 & x4 ) | ( x1 & ~n8 ) | ( x4 & ~n8 ) ;
  assign n10 = x0 & n9 ;
  assign n11 = x1 & ~x2 ;
  assign n12 = x3 & ~x4 ;
  assign n13 = ( x2 & ~x3 ) | ( x2 & n12 ) | ( ~x3 & n12 ) ;
  assign n14 = ( ~x1 & x2 ) | ( ~x1 & n13 ) | ( x2 & n13 ) ;
  assign n15 = ( n11 & ~n13 ) | ( n11 & n14 ) | ( ~n13 & n14 ) ;
  assign n16 = x0 & ~n15 ;
  assign n17 = ( x0 & x3 ) | ( x0 & x4 ) | ( x3 & x4 ) ;
  assign n18 = ( x0 & x3 ) | ( x0 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n19 = n17 & ~n18 ;
  assign n20 = x2 & ~x4 ;
  assign n21 = x3 & n20 ;
  assign n22 = x1 | x3 ;
  assign n23 = ( x0 & ~x2 ) | ( x0 & n22 ) | ( ~x2 & n22 ) ;
  assign n24 = ( x0 & x3 ) | ( x0 & ~n22 ) | ( x3 & ~n22 ) ;
  assign n25 = ( x1 & ~n23 ) | ( x1 & n24 ) | ( ~n23 & n24 ) ;
  assign n26 = ( x0 & ~x1 ) | ( x0 & n25 ) | ( ~x1 & n25 ) ;
  assign n27 = n21 & ~n26 ;
  assign n28 = ( n21 & n25 ) | ( n21 & ~n27 ) | ( n25 & ~n27 ) ;
  assign n29 = ( x1 & ~x2 ) | ( x1 & n28 ) | ( ~x2 & n28 ) ;
  assign n30 = n19 & ~n29 ;
  assign n31 = ( n19 & n28 ) | ( n19 & ~n30 ) | ( n28 & ~n30 ) ;
  assign n34 = ( x1 & ~x3 ) | ( x1 & x5 ) | ( ~x3 & x5 ) ;
  assign n35 = ( x2 & ~x5 ) | ( x2 & n34 ) | ( ~x5 & n34 ) ;
  assign n36 = ( x1 & x2 ) | ( x1 & ~n34 ) | ( x2 & ~n34 ) ;
  assign n37 = n35 & ~n36 ;
  assign n38 = x0 & ~n37 ;
  assign n32 = ~x2 & x3 ;
  assign n33 = ~x5 & n32 ;
  assign n39 = x1 & n33 ;
  assign n40 = x0 | n39 ;
  assign n41 = ~n38 & n40 ;
  assign n57 = ~x4 & n41 ;
  assign n42 = ( x0 & ~x2 ) | ( x0 & x3 ) | ( ~x2 & x3 ) ;
  assign n43 = ( ~x0 & x1 ) | ( ~x0 & n42 ) | ( x1 & n42 ) ;
  assign n44 = ( ~x2 & x3 ) | ( ~x2 & n43 ) | ( x3 & n43 ) ;
  assign n45 = ~n42 & n44 ;
  assign n46 = ( ~n43 & n44 ) | ( ~n43 & n45 ) | ( n44 & n45 ) ;
  assign n48 = ( x1 & ~x2 ) | ( x1 & x3 ) | ( ~x2 & x3 ) ;
  assign n49 = x1 & x4 ;
  assign n50 = ( x3 & ~n48 ) | ( x3 & n49 ) | ( ~n48 & n49 ) ;
  assign n51 = ( ~x4 & n48 ) | ( ~x4 & n50 ) | ( n48 & n50 ) ;
  assign n52 = ( ~x3 & n50 ) | ( ~x3 & n51 ) | ( n50 & n51 ) ;
  assign n53 = x0 & ~n52 ;
  assign n47 = ~x4 & n32 ;
  assign n54 = x1 & n47 ;
  assign n55 = x0 | n54 ;
  assign n56 = ~n53 & n55 ;
  assign n58 = n46 | n56 ;
  assign n59 = ( n41 & ~n57 ) | ( n41 & n58 ) | ( ~n57 & n58 ) ;
  assign n62 = ( x1 & x2 ) | ( x1 & ~x5 ) | ( x2 & ~x5 ) ;
  assign n63 = n7 | n62 ;
  assign n64 = x5 & n63 ;
  assign n65 = ( ~n7 & n63 ) | ( ~n7 & n64 ) | ( n63 & n64 ) ;
  assign n66 = x4 & ~n65 ;
  assign n60 = ~x3 & x5 ;
  assign n61 = ( x1 & x5 ) | ( x1 & n60 ) | ( x5 & n60 ) ;
  assign n67 = x2 & n61 ;
  assign n68 = x4 | n67 ;
  assign n69 = ~n66 & n68 ;
  assign n86 = ~x0 & n69 ;
  assign n72 = x4 & ~x5 ;
  assign n70 = ~x0 & x1 ;
  assign n71 = ~x2 & n70 ;
  assign n73 = x3 & n71 ;
  assign n74 = n72 & n73 ;
  assign n77 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n78 = x2 | n77 ;
  assign n79 = ( x0 & ~x3 ) | ( x0 & n77 ) | ( ~x3 & n77 ) ;
  assign n80 = x2 & n79 ;
  assign n81 = n78 & ~n80 ;
  assign n82 = x4 & ~n81 ;
  assign n75 = x1 | x2 ;
  assign n76 = ( ~x1 & n11 ) | ( ~x1 & n75 ) | ( n11 & n75 ) ;
  assign n83 = x3 & n76 ;
  assign n84 = x4 | n83 ;
  assign n85 = ~n82 & n84 ;
  assign n87 = n74 | n85 ;
  assign n88 = ( n69 & ~n86 ) | ( n69 & n87 ) | ( ~n86 & n87 ) ;
  assign n89 = x2 | x3 ;
  assign n90 = ( x0 & ~x2 ) | ( x0 & n89 ) | ( ~x2 & n89 ) ;
  assign n91 = ( x0 & ~x1 ) | ( x0 & n89 ) | ( ~x1 & n89 ) ;
  assign n92 = ( n11 & ~n90 ) | ( n11 & n91 ) | ( ~n90 & n91 ) ;
  assign n126 = ~x4 & n92 ;
  assign n93 = x2 & ~x3 ;
  assign n94 = ( x0 & ~x4 ) | ( x0 & n93 ) | ( ~x4 & n93 ) ;
  assign n95 = ~x0 & n94 ;
  assign n96 = ( x0 & ~x3 ) | ( x0 & x5 ) | ( ~x3 & x5 ) ;
  assign n97 = ( ~x1 & x5 ) | ( ~x1 & n96 ) | ( x5 & n96 ) ;
  assign n98 = x5 & ~n97 ;
  assign n99 = n97 | n98 ;
  assign n100 = ( ~x5 & n98 ) | ( ~x5 & n99 ) | ( n98 & n99 ) ;
  assign n123 = ~x2 & n100 ;
  assign n101 = ~x2 & x5 ;
  assign n102 = ( x0 & x1 ) | ( x0 & n101 ) | ( x1 & n101 ) ;
  assign n103 = ~x1 & n102 ;
  assign n111 = ( x2 & x5 ) | ( x2 & n18 ) | ( x5 & n18 ) ;
  assign n112 = ( x0 & x3 ) | ( x0 & n111 ) | ( x3 & n111 ) ;
  assign n113 = n18 & ~n112 ;
  assign n114 = ( n111 & ~n112 ) | ( n111 & n113 ) | ( ~n112 & n113 ) ;
  assign n115 = x4 & ~n114 ;
  assign n107 = x2 | x5 ;
  assign n108 = x3 | x5 ;
  assign n109 = x2 & ~n108 ;
  assign n110 = ( ~x2 & n107 ) | ( ~x2 & n109 ) | ( n107 & n109 ) ;
  assign n116 = x0 & n110 ;
  assign n117 = x4 | n116 ;
  assign n118 = ~n115 & n117 ;
  assign n119 = x1 & ~n118 ;
  assign n104 = ( x2 & x4 ) | ( x2 & x5 ) | ( x4 & x5 ) ;
  assign n105 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n106 = n104 & ~n105 ;
  assign n120 = x0 & n106 ;
  assign n121 = x1 | n120 ;
  assign n122 = ~n119 & n121 ;
  assign n124 = n103 | n122 ;
  assign n125 = ( n100 & ~n123 ) | ( n100 & n124 ) | ( ~n123 & n124 ) ;
  assign n127 = n95 | n125 ;
  assign n128 = ( n92 & ~n126 ) | ( n92 & n127 ) | ( ~n126 & n127 ) ;
  assign n130 = ( x2 & x3 ) | ( x2 & x4 ) | ( x3 & x4 ) ;
  assign n131 = x1 & ~n130 ;
  assign n132 = ~x1 & n130 ;
  assign n133 = n131 | n132 ;
  assign n134 = x5 & ~n133 ;
  assign n129 = ( ~x2 & n89 ) | ( ~x2 & n93 ) | ( n89 & n93 ) ;
  assign n135 = x4 & n129 ;
  assign n136 = x5 | n135 ;
  assign n137 = ~n134 & n136 ;
  assign n138 = ( x2 & x3 ) | ( x2 & x5 ) | ( x3 & x5 ) ;
  assign n139 = x3 & x4 ;
  assign n140 = ( x3 & x5 ) | ( x3 & n139 ) | ( x5 & n139 ) ;
  assign n141 = ( n32 & n138 ) | ( n32 & ~n140 ) | ( n138 & ~n140 ) ;
  assign n142 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n143 = ~x4 & n142 ;
  assign n144 = ( ~x3 & n142 ) | ( ~x3 & n143 ) | ( n142 & n143 ) ;
  assign y0 = n10 ;
  assign y1 = n16 ;
  assign y2 = n31 ;
  assign y3 = n59 ;
  assign y4 = n88 ;
  assign y5 = n128 ;
  assign y6 = n137 ;
  assign y7 = n141 ;
  assign y8 = n144 ;
  assign y9 = n72 ;
  assign y10 = 1'b0 ;
  assign y11 = x5 ;
endmodule
