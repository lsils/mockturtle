module top( b_4_ , a_6_ , a_7_ , a_1_ , a_0_ , a_2_ , c , b_7_ , a_5_ , b_3_ , b_2_ , b_1_ , b_6_ , a_3_ , b_5_ , a_4_ , b_0_ , cout , s_6_ , s_3_ , s_4_ , s_5_ , s_0_ , s_2_ , s_7_ , s_1_ );
  input b_4_ , a_6_ , a_7_ , a_1_ , a_0_ , a_2_ , c , b_7_ , a_5_ , b_3_ , b_2_ , b_1_ , b_6_ , a_3_ , b_5_ , a_4_ , b_0_ ;
  output cout , s_6_ , s_3_ , s_4_ , s_5_ , s_0_ , s_2_ , s_7_ , s_1_ ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 ;
  assign n18 = a_7_ & b_7_ ;
  assign n19 = a_7_ | b_7_ ;
  assign n20 = ~n18 & n19 ;
  assign n21 = a_6_ & b_6_ ;
  assign n22 = a_6_ | b_6_ ;
  assign n23 = ~n21 & n22 ;
  assign n24 = a_5_ & b_5_ ;
  assign n25 = b_4_ & a_4_ ;
  assign n26 = b_3_ & a_3_ ;
  assign n27 = b_3_ | a_3_ ;
  assign n28 = ~n26 & n27 ;
  assign n29 = a_2_ & b_2_ ;
  assign n30 = a_2_ | b_2_ ;
  assign n31 = ~n29 & n30 ;
  assign n32 = a_1_ & b_1_ ;
  assign n33 = a_1_ | b_1_ ;
  assign n34 = a_0_ & b_0_ ;
  assign n35 = n33 & n34 ;
  assign n36 = n32 | n35 ;
  assign n37 = n31 & n36 ;
  assign n38 = n29 | n37 ;
  assign n39 = n28 & n38 ;
  assign n40 = n26 | n39 ;
  assign n41 = b_4_ | a_4_ ;
  assign n42 = ~n25 & n41 ;
  assign n43 = n40 & n42 ;
  assign n44 = n25 | n43 ;
  assign n45 = a_5_ | b_5_ ;
  assign n46 = ~n24 & n45 ;
  assign n47 = n44 & n46 ;
  assign n48 = n24 | n47 ;
  assign n49 = n23 & n48 ;
  assign n50 = n21 | n49 ;
  assign n51 = n20 & n50 ;
  assign n52 = n18 | n51 ;
  assign n53 = n20 | n50 ;
  assign n54 = ~n51 & n53 ;
  assign n55 = n23 | n48 ;
  assign n56 = ~n49 & n55 ;
  assign n57 = n40 | n42 ;
  assign n58 = ~n43 & n57 ;
  assign n59 = n28 | n38 ;
  assign n60 = ~n39 & n59 ;
  assign n61 = n31 | n36 ;
  assign n62 = ~n37 & n61 ;
  assign n63 = ~n32 & n33 ;
  assign n64 = a_0_ | b_0_ ;
  assign n65 = ~n34 & n64 ;
  assign n66 = c & n65 ;
  assign n67 = n63 & n66 ;
  assign n68 = n62 & n67 ;
  assign n69 = n60 & n68 ;
  assign n70 = n58 & n69 ;
  assign n71 = n44 | n46 ;
  assign n72 = ~n47 & n71 ;
  assign n73 = n70 & n72 ;
  assign n74 = n56 & n73 ;
  assign n75 = n54 & n74 ;
  assign n76 = n52 | n75 ;
  assign n77 = n56 | n73 ;
  assign n78 = ~n74 & n77 ;
  assign n79 = n60 | n68 ;
  assign n80 = ~n69 & n79 ;
  assign n81 = n58 | n69 ;
  assign n82 = ~n70 & n81 ;
  assign n83 = n70 | n72 ;
  assign n84 = ~n73 & n83 ;
  assign n85 = c | n65 ;
  assign n86 = ~n66 & n85 ;
  assign n87 = n62 | n67 ;
  assign n88 = ~n68 & n87 ;
  assign n89 = n54 | n74 ;
  assign n90 = ~n75 & n89 ;
  assign n91 = n34 | n66 ;
  assign n92 = n63 | n91 ;
  assign n93 = n63 & n91 ;
  assign n94 = n92 & ~n93 ;
  assign cout = n76 ;
  assign s_6_ = n78 ;
  assign s_3_ = n80 ;
  assign s_4_ = n82 ;
  assign s_5_ = n84 ;
  assign s_0_ = n86 ;
  assign s_2_ = n88 ;
  assign s_7_ = n90 ;
  assign s_1_ = n94 ;
endmodule
