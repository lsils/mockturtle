module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 ;
  wire n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 ;
  assign n136 = x72 & ~x75 ;
  assign n137 = ~x72 & x92 ;
  assign n138 = x91 & n137 ;
  assign n139 = x83 & n138 ;
  assign n140 = x2 | x3 ;
  assign n141 = x39 & ~n140 ;
  assign n142 = ( n139 & ~n140 ) | ( n139 & n141 ) | ( ~n140 & n141 ) ;
  assign n143 = x1 & ~x73 ;
  assign n144 = ( x73 & n142 ) | ( x73 & ~n143 ) | ( n142 & ~n143 ) ;
  assign n145 = ( x28 & ~x37 ) | ( x28 & x79 ) | ( ~x37 & x79 ) ;
  assign n146 = ( x79 & x80 ) | ( x79 & ~n145 ) | ( x80 & ~n145 ) ;
  assign n147 = ( ~x28 & x80 ) | ( ~x28 & n145 ) | ( x80 & n145 ) ;
  assign n148 = n146 & ~n147 ;
  assign n149 = ( x73 & ~x75 ) | ( x73 & n148 ) | ( ~x75 & n148 ) ;
  assign n150 = ~x34 & x86 ;
  assign n151 = x35 & ~x86 ;
  assign n152 = ( x86 & ~n150 ) | ( x86 & n151 ) | ( ~n150 & n151 ) ;
  assign n153 = x87 & x88 ;
  assign n154 = x87 & ~n153 ;
  assign n155 = n152 & n154 ;
  assign n156 = ~x32 & x86 ;
  assign n157 = x33 & ~x86 ;
  assign n158 = ( x86 & ~n156 ) | ( x86 & n157 ) | ( ~n156 & n157 ) ;
  assign n159 = ( ~n153 & n154 ) | ( ~n153 & n158 ) | ( n154 & n158 ) ;
  assign n160 = ( x88 & n155 ) | ( x88 & n159 ) | ( n155 & n159 ) ;
  assign n161 = x83 & x92 ;
  assign n162 = ( x83 & x91 ) | ( x83 & n161 ) | ( x91 & n161 ) ;
  assign n163 = x84 | x85 ;
  assign n164 = ( x75 & ~n162 ) | ( x75 & n163 ) | ( ~n162 & n163 ) ;
  assign n165 = ( ~n136 & n162 ) | ( ~n136 & n164 ) | ( n162 & n164 ) ;
  assign n166 = x90 | n165 ;
  assign n167 = ( x89 & n160 ) | ( x89 & n166 ) | ( n160 & n166 ) ;
  assign n168 = n160 & ~n167 ;
  assign n169 = x74 & x91 ;
  assign n170 = x28 & ~x91 ;
  assign n171 = ( x91 & ~n169 ) | ( x91 & n170 ) | ( ~n169 & n170 ) ;
  assign n172 = x92 & ~n171 ;
  assign n173 = ~x27 & x91 ;
  assign n174 = x92 | n173 ;
  assign n175 = ~n172 & n174 ;
  assign n176 = x83 & n175 ;
  assign n177 = x109 & ~n162 ;
  assign n178 = n176 | n177 ;
  assign n179 = ( n163 & n176 ) | ( n163 & n178 ) | ( n176 & n178 ) ;
  assign n180 = ( ~x72 & n168 ) | ( ~x72 & n179 ) | ( n168 & n179 ) ;
  assign n181 = x75 | n180 ;
  assign n182 = ( ~x75 & n168 ) | ( ~x75 & n181 ) | ( n168 & n181 ) ;
  assign n183 = ~x73 & n182 ;
  assign n184 = ( n148 & ~n149 ) | ( n148 & n183 ) | ( ~n149 & n183 ) ;
  assign n185 = ( x38 & x81 ) | ( x38 & ~x82 ) | ( x81 & ~x82 ) ;
  assign n186 = ~x38 & x77 ;
  assign n187 = ( x81 & ~n185 ) | ( x81 & n186 ) | ( ~n185 & n186 ) ;
  assign n188 = x16 & ~x73 ;
  assign n189 = ( x7 & x73 ) | ( x7 & ~n188 ) | ( x73 & ~n188 ) ;
  assign n190 = x40 & ~n189 ;
  assign n191 = x7 & ~x16 ;
  assign n192 = ~x73 & n191 ;
  assign n193 = n190 | n192 ;
  assign n194 = ( x8 & n190 ) | ( x8 & n193 ) | ( n190 & n193 ) ;
  assign n195 = x41 & ~n189 ;
  assign n196 = n192 | n195 ;
  assign n197 = ( x9 & n195 ) | ( x9 & n196 ) | ( n195 & n196 ) ;
  assign n198 = x42 & ~n189 ;
  assign n199 = n192 | n198 ;
  assign n200 = ( x10 & n198 ) | ( x10 & n199 ) | ( n198 & n199 ) ;
  assign n201 = x43 & ~n189 ;
  assign n202 = n192 | n201 ;
  assign n203 = ( x11 & n201 ) | ( x11 & n202 ) | ( n201 & n202 ) ;
  assign n204 = x44 & ~n189 ;
  assign n205 = n192 | n204 ;
  assign n206 = ( x12 & n204 ) | ( x12 & n205 ) | ( n204 & n205 ) ;
  assign n207 = x45 & ~n189 ;
  assign n208 = n192 | n207 ;
  assign n209 = ( x13 & n207 ) | ( x13 & n208 ) | ( n207 & n208 ) ;
  assign n210 = x46 & ~n189 ;
  assign n211 = n192 | n210 ;
  assign n212 = ( x14 & n210 ) | ( x14 & n211 ) | ( n210 & n211 ) ;
  assign n213 = x47 & ~n189 ;
  assign n214 = n192 | n213 ;
  assign n215 = ( x15 & n213 ) | ( x15 & n214 ) | ( n213 & n214 ) ;
  assign n216 = x16 | x73 ;
  assign n217 = ( x7 & x73 ) | ( x7 & n216 ) | ( x73 & n216 ) ;
  assign n218 = x48 & ~n217 ;
  assign n219 = x7 & ~x73 ;
  assign n220 = x16 & n219 ;
  assign n221 = n218 | n220 ;
  assign n222 = ( x8 & n218 ) | ( x8 & n221 ) | ( n218 & n221 ) ;
  assign n223 = x49 & ~n217 ;
  assign n224 = n220 | n223 ;
  assign n225 = ( x9 & n223 ) | ( x9 & n224 ) | ( n223 & n224 ) ;
  assign n226 = x50 & ~n217 ;
  assign n227 = n220 | n226 ;
  assign n228 = ( x10 & n226 ) | ( x10 & n227 ) | ( n226 & n227 ) ;
  assign n229 = x51 & ~n217 ;
  assign n230 = n220 | n229 ;
  assign n231 = ( x11 & n229 ) | ( x11 & n230 ) | ( n229 & n230 ) ;
  assign n232 = x52 & ~n217 ;
  assign n233 = n220 | n232 ;
  assign n234 = ( x12 & n232 ) | ( x12 & n233 ) | ( n232 & n233 ) ;
  assign n235 = x53 & ~n217 ;
  assign n236 = n220 | n235 ;
  assign n237 = ( x13 & n235 ) | ( x13 & n236 ) | ( n235 & n236 ) ;
  assign n238 = x54 & ~n217 ;
  assign n239 = n220 | n238 ;
  assign n240 = ( x14 & n238 ) | ( x14 & n239 ) | ( n238 & n239 ) ;
  assign n241 = x55 & ~n217 ;
  assign n242 = n220 | n241 ;
  assign n243 = ( x15 & n241 ) | ( x15 & n242 ) | ( n241 & n242 ) ;
  assign n244 = x26 & ~x73 ;
  assign n245 = ( x17 & x73 ) | ( x17 & ~n244 ) | ( x73 & ~n244 ) ;
  assign n246 = x56 & ~n245 ;
  assign n247 = x17 & ~x26 ;
  assign n248 = ~x73 & n247 ;
  assign n249 = n246 | n248 ;
  assign n250 = ( x18 & n246 ) | ( x18 & n249 ) | ( n246 & n249 ) ;
  assign n251 = x57 & ~n245 ;
  assign n252 = n248 | n251 ;
  assign n253 = ( x19 & n251 ) | ( x19 & n252 ) | ( n251 & n252 ) ;
  assign n254 = x58 & ~n245 ;
  assign n255 = n248 | n254 ;
  assign n256 = ( x20 & n254 ) | ( x20 & n255 ) | ( n254 & n255 ) ;
  assign n257 = x59 & ~n245 ;
  assign n258 = n248 | n257 ;
  assign n259 = ( x21 & n257 ) | ( x21 & n258 ) | ( n257 & n258 ) ;
  assign n260 = x60 & ~n245 ;
  assign n261 = n248 | n260 ;
  assign n262 = ( x22 & n260 ) | ( x22 & n261 ) | ( n260 & n261 ) ;
  assign n263 = x61 & ~n245 ;
  assign n264 = n248 | n263 ;
  assign n265 = ( x23 & n263 ) | ( x23 & n264 ) | ( n263 & n264 ) ;
  assign n266 = x62 & ~n245 ;
  assign n267 = n248 | n266 ;
  assign n268 = ( x24 & n266 ) | ( x24 & n267 ) | ( n266 & n267 ) ;
  assign n269 = x63 & ~n245 ;
  assign n270 = n248 | n269 ;
  assign n271 = ( x25 & n269 ) | ( x25 & n270 ) | ( n269 & n270 ) ;
  assign n272 = x26 | x73 ;
  assign n273 = ( x17 & x73 ) | ( x17 & n272 ) | ( x73 & n272 ) ;
  assign n274 = x64 & ~n273 ;
  assign n275 = x17 & ~x73 ;
  assign n276 = x26 & n275 ;
  assign n277 = n274 | n276 ;
  assign n278 = ( x18 & n274 ) | ( x18 & n277 ) | ( n274 & n277 ) ;
  assign n279 = x65 & ~n273 ;
  assign n280 = n276 | n279 ;
  assign n281 = ( x19 & n279 ) | ( x19 & n280 ) | ( n279 & n280 ) ;
  assign n282 = x66 & ~n273 ;
  assign n283 = n276 | n282 ;
  assign n284 = ( x20 & n282 ) | ( x20 & n283 ) | ( n282 & n283 ) ;
  assign n285 = x67 & ~n273 ;
  assign n286 = n276 | n285 ;
  assign n287 = ( x21 & n285 ) | ( x21 & n286 ) | ( n285 & n286 ) ;
  assign n288 = x68 & ~n273 ;
  assign n289 = n276 | n288 ;
  assign n290 = ( x22 & n288 ) | ( x22 & n289 ) | ( n288 & n289 ) ;
  assign n291 = x69 & ~n273 ;
  assign n292 = n276 | n291 ;
  assign n293 = ( x23 & n291 ) | ( x23 & n292 ) | ( n291 & n292 ) ;
  assign n294 = x70 & ~n273 ;
  assign n295 = n276 | n294 ;
  assign n296 = ( x24 & n294 ) | ( x24 & n295 ) | ( n294 & n295 ) ;
  assign n297 = x71 & ~n273 ;
  assign n298 = n276 | n297 ;
  assign n299 = ( x25 & n297 ) | ( x25 & n298 ) | ( n297 & n298 ) ;
  assign n300 = ~x1 & x72 ;
  assign n301 = ~n140 & n300 ;
  assign n302 = x73 | n301 ;
  assign n303 = x38 | n139 ;
  assign n304 = ~x109 & n163 ;
  assign n305 = ~x90 & n160 ;
  assign n306 = ~x89 & n305 ;
  assign n307 = n163 | n306 ;
  assign n308 = ~n304 & n307 ;
  assign n309 = ( x74 & n162 ) | ( x74 & ~n308 ) | ( n162 & ~n308 ) ;
  assign n310 = x72 & x74 ;
  assign n311 = ( ~n162 & n309 ) | ( ~n162 & n310 ) | ( n309 & n310 ) ;
  assign n312 = x74 | n162 ;
  assign n313 = ( x72 & n308 ) | ( x72 & n312 ) | ( n308 & n312 ) ;
  assign n314 = n308 & ~n313 ;
  assign n315 = x27 & x91 ;
  assign n316 = x92 | n315 ;
  assign n317 = ( ~x28 & n315 ) | ( ~x28 & n316 ) | ( n315 & n316 ) ;
  assign n318 = x74 & ~n317 ;
  assign n319 = ( x28 & n173 ) | ( x28 & n174 ) | ( n173 & n174 ) ;
  assign n320 = ~x72 & n319 ;
  assign n321 = x74 | n320 ;
  assign n322 = ~n318 & n321 ;
  assign n323 = ( x83 & n139 ) | ( x83 & n322 ) | ( n139 & n322 ) ;
  assign n324 = ( ~x73 & n314 ) | ( ~x73 & n323 ) | ( n314 & n323 ) ;
  assign n325 = ~n311 & n324 ;
  assign n326 = ( ~x73 & n311 ) | ( ~x73 & n325 ) | ( n311 & n325 ) ;
  assign n327 = ~x35 & x133 ;
  assign n328 = ( x34 & ~x132 ) | ( x34 & n327 ) | ( ~x132 & n327 ) ;
  assign n329 = x35 & ~x133 ;
  assign n330 = ( ~x34 & x132 ) | ( ~x34 & n329 ) | ( x132 & n329 ) ;
  assign n331 = n328 | n330 ;
  assign n332 = x126 & x128 ;
  assign n333 = ( ~x125 & x127 ) | ( ~x125 & n332 ) | ( x127 & n332 ) ;
  assign n334 = x125 & n333 ;
  assign n335 = x134 & n334 ;
  assign n336 = ( x129 & n331 ) | ( x129 & n335 ) | ( n331 & n335 ) ;
  assign n337 = ~n331 & n336 ;
  assign n338 = ( ~x33 & x131 ) | ( ~x33 & n337 ) | ( x131 & n337 ) ;
  assign n339 = ~x131 & n338 ;
  assign n340 = ( x33 & n338 ) | ( x33 & n339 ) | ( n338 & n339 ) ;
  assign n341 = ( x32 & x130 ) | ( x32 & n340 ) | ( x130 & n340 ) ;
  assign n342 = ~x130 & n341 ;
  assign n343 = ( ~x32 & n341 ) | ( ~x32 & n342 ) | ( n341 & n342 ) ;
  assign n344 = ~x35 & x78 ;
  assign n345 = ( x34 & x36 ) | ( x34 & n344 ) | ( x36 & n344 ) ;
  assign n346 = ~x34 & n345 ;
  assign n347 = x75 & ~x80 ;
  assign n348 = ( x75 & ~x79 ) | ( x75 & n347 ) | ( ~x79 & n347 ) ;
  assign n349 = ( x32 & x33 ) | ( x32 & ~n348 ) | ( x33 & ~n348 ) ;
  assign n350 = n346 & n349 ;
  assign n351 = ( n346 & n348 ) | ( n346 & ~n350 ) | ( n348 & ~n350 ) ;
  assign n352 = ~x73 & n351 ;
  assign n353 = ( ~x73 & n343 ) | ( ~x73 & n352 ) | ( n343 & n352 ) ;
  assign n354 = x36 | x38 ;
  assign n355 = x130 & ~x131 ;
  assign n356 = ~x132 & n355 ;
  assign n357 = x127 & x129 ;
  assign n358 = ( ~x126 & x128 ) | ( ~x126 & n357 ) | ( x128 & n357 ) ;
  assign n359 = x126 & n358 ;
  assign n360 = ~x133 & n359 ;
  assign n361 = n356 & n360 ;
  assign n362 = ( x125 & n354 ) | ( x125 & n361 ) | ( n354 & n361 ) ;
  assign n363 = ~x76 & n362 ;
  assign n364 = ( x76 & n354 ) | ( x76 & ~n362 ) | ( n354 & ~n362 ) ;
  assign n365 = ( ~n354 & n363 ) | ( ~n354 & n364 ) | ( n363 & n364 ) ;
  assign n366 = ( x76 & n354 ) | ( x76 & n361 ) | ( n354 & n361 ) ;
  assign n367 = x125 & ~n366 ;
  assign n368 = ( x125 & n354 ) | ( x125 & ~n367 ) | ( n354 & ~n367 ) ;
  assign n369 = x77 & n368 ;
  assign n370 = x125 & n361 ;
  assign n371 = ~n354 & n370 ;
  assign n372 = x76 & n371 ;
  assign n373 = x77 | n372 ;
  assign n374 = ~n369 & n373 ;
  assign n375 = ~x36 & x78 ;
  assign n376 = x0 & ~x38 ;
  assign n377 = ( x36 & n375 ) | ( x36 & n376 ) | ( n375 & n376 ) ;
  assign n378 = ~x82 & n377 ;
  assign n379 = ( ~x81 & n377 ) | ( ~x81 & n378 ) | ( n377 & n378 ) ;
  assign n380 = x36 & ~x38 ;
  assign n381 = x33 | x35 ;
  assign n382 = x34 | n381 ;
  assign n383 = x78 & ~n382 ;
  assign n384 = ( x32 & n380 ) | ( x32 & n383 ) | ( n380 & n383 ) ;
  assign n385 = ~x32 & n384 ;
  assign n386 = ( x75 & ~n343 ) | ( x75 & n385 ) | ( ~n343 & n385 ) ;
  assign n387 = x38 & ~n385 ;
  assign n388 = ( n343 & n386 ) | ( n343 & ~n387 ) | ( n386 & ~n387 ) ;
  assign n389 = x79 | n388 ;
  assign n390 = x35 | x133 ;
  assign n391 = x125 & x132 ;
  assign n392 = ( x35 & ~n390 ) | ( x35 & n391 ) | ( ~n390 & n391 ) ;
  assign n393 = x34 | n392 ;
  assign n394 = ~x34 & x132 ;
  assign n395 = x133 | n394 ;
  assign n396 = ( ~x35 & n394 ) | ( ~x35 & n395 ) | ( n394 & n395 ) ;
  assign n397 = x125 & ~n396 ;
  assign n398 = x130 & n359 ;
  assign n399 = ( x32 & n359 ) | ( x32 & n398 ) | ( n359 & n398 ) ;
  assign n400 = x131 & x134 ;
  assign n401 = ( ~x33 & n399 ) | ( ~x33 & n400 ) | ( n399 & n400 ) ;
  assign n402 = n397 & ~n401 ;
  assign n403 = ( x33 & ~n397 ) | ( x33 & n402 ) | ( ~n397 & n402 ) ;
  assign n404 = x34 | x132 ;
  assign n405 = x125 & x133 ;
  assign n406 = ( x34 & ~n404 ) | ( x34 & n405 ) | ( ~n404 & n405 ) ;
  assign n407 = ~x36 & n396 ;
  assign n408 = x35 | n407 ;
  assign n409 = ( ~n406 & n407 ) | ( ~n406 & n408 ) | ( n407 & n408 ) ;
  assign n410 = n403 | n409 ;
  assign n411 = ( ~n392 & n393 ) | ( ~n392 & n410 ) | ( n393 & n410 ) ;
  assign n412 = x78 & ~n397 ;
  assign n413 = ~x130 & n359 ;
  assign n414 = ~x131 & x134 ;
  assign n415 = ( x33 & x134 ) | ( x33 & n414 ) | ( x134 & n414 ) ;
  assign n416 = ( ~x32 & n413 ) | ( ~x32 & n415 ) | ( n413 & n415 ) ;
  assign n417 = n397 & ~n416 ;
  assign n418 = ( x32 & ~n397 ) | ( x32 & n417 ) | ( ~n397 & n417 ) ;
  assign n419 = n346 | n415 ;
  assign n420 = ( n346 & n399 ) | ( n346 & n419 ) | ( n399 & n419 ) ;
  assign n421 = ~n418 & n420 ;
  assign n422 = ( n397 & n412 ) | ( n397 & n421 ) | ( n412 & n421 ) ;
  assign n423 = x125 | n354 ;
  assign n424 = ( n411 & n422 ) | ( n411 & n423 ) | ( n422 & n423 ) ;
  assign n425 = x38 & n423 ;
  assign n426 = ( ~n411 & n424 ) | ( ~n411 & n425 ) | ( n424 & n425 ) ;
  assign n427 = x75 | n426 ;
  assign n428 = x79 & n427 ;
  assign n429 = n389 & ~n428 ;
  assign n430 = ( x38 & n427 ) | ( x38 & n428 ) | ( n427 & n428 ) ;
  assign n431 = x80 & n430 ;
  assign n432 = x79 & n388 ;
  assign n433 = x80 | n432 ;
  assign n434 = ~n431 & n433 ;
  assign n435 = ~x38 & x82 ;
  assign n436 = ( ~x84 & x89 ) | ( ~x84 & x90 ) | ( x89 & x90 ) ;
  assign n437 = x89 & n436 ;
  assign n438 = x89 | x90 ;
  assign n439 = ( x31 & n437 ) | ( x31 & ~n438 ) | ( n437 & ~n438 ) ;
  assign n440 = n437 | n439 ;
  assign n441 = ~x87 & x88 ;
  assign n442 = x86 & n441 ;
  assign n443 = ~n440 & n442 ;
  assign n444 = ( x72 & ~x73 ) | ( x72 & n443 ) | ( ~x73 & n443 ) ;
  assign n445 = ~x73 & x83 ;
  assign n446 = ( ~x72 & n444 ) | ( ~x72 & n445 ) | ( n444 & n445 ) ;
  assign n447 = x30 & x31 ;
  assign n448 = ( x29 & x31 ) | ( x29 & n447 ) | ( x31 & n447 ) ;
  assign n449 = x89 | n448 ;
  assign n450 = ~x72 & n442 ;
  assign n451 = ( x90 & n449 ) | ( x90 & ~n450 ) | ( n449 & ~n450 ) ;
  assign n452 = n449 & ~n451 ;
  assign n453 = ( ~x73 & x84 ) | ( ~x73 & n452 ) | ( x84 & n452 ) ;
  assign n454 = x72 | x90 ;
  assign n455 = x89 | n454 ;
  assign n456 = n442 & n448 ;
  assign n457 = ( x84 & ~n455 ) | ( x84 & n456 ) | ( ~n455 & n456 ) ;
  assign n458 = ~x84 & n457 ;
  assign n459 = ~x73 & n458 ;
  assign n460 = ( ~n452 & n453 ) | ( ~n452 & n459 ) | ( n453 & n459 ) ;
  assign n461 = ( x29 & x30 ) | ( x29 & ~x90 ) | ( x30 & ~x90 ) ;
  assign n462 = x31 & n461 ;
  assign n463 = ( x31 & x90 ) | ( x31 & ~n462 ) | ( x90 & ~n462 ) ;
  assign n464 = ( x89 & ~n450 ) | ( x89 & n463 ) | ( ~n450 & n463 ) ;
  assign n465 = n463 & ~n464 ;
  assign n466 = ( x73 & x85 ) | ( x73 & n465 ) | ( x85 & n465 ) ;
  assign n467 = n465 & ~n466 ;
  assign n468 = ( x85 & ~n466 ) | ( x85 & n467 ) | ( ~n466 & n467 ) ;
  assign n469 = ( x73 & x86 ) | ( x73 & ~n301 ) | ( x86 & ~n301 ) ;
  assign n470 = n301 | n469 ;
  assign n471 = ( ~x86 & n469 ) | ( ~x86 & n470 ) | ( n469 & n470 ) ;
  assign n472 = ~x87 & n469 ;
  assign n473 = ( x73 & x87 ) | ( x73 & ~n469 ) | ( x87 & ~n469 ) ;
  assign n474 = ( ~x73 & n472 ) | ( ~x73 & n473 ) | ( n472 & n473 ) ;
  assign n475 = x87 & ~n469 ;
  assign n476 = ( x73 & x87 ) | ( x73 & ~n475 ) | ( x87 & ~n475 ) ;
  assign n477 = x88 & n476 ;
  assign n478 = x87 & ~n302 ;
  assign n479 = x86 & n478 ;
  assign n480 = ~x88 & n479 ;
  assign n481 = ( x88 & ~n477 ) | ( x88 & n480 ) | ( ~n477 & n480 ) ;
  assign n482 = x86 & x88 ;
  assign n483 = ( x87 & n301 ) | ( x87 & n482 ) | ( n301 & n482 ) ;
  assign n484 = ~n301 & n483 ;
  assign n485 = x73 | n484 ;
  assign n486 = x89 & n485 ;
  assign n487 = x88 & n479 ;
  assign n488 = x89 | n487 ;
  assign n489 = ~n486 & n488 ;
  assign n490 = ~x89 & n484 ;
  assign n491 = ~x73 & x90 ;
  assign n492 = ( ~n484 & n490 ) | ( ~n484 & n491 ) | ( n490 & n491 ) ;
  assign n493 = x88 & x89 ;
  assign n494 = ( ~x90 & n492 ) | ( ~x90 & n493 ) | ( n492 & n493 ) ;
  assign n495 = n479 & ~n494 ;
  assign n496 = ( n479 & n492 ) | ( n479 & ~n495 ) | ( n492 & ~n495 ) ;
  assign n497 = ~x72 & x83 ;
  assign n498 = ( ~x72 & n443 ) | ( ~x72 & n497 ) | ( n443 & n497 ) ;
  assign n499 = ( x73 & x91 ) | ( x73 & n498 ) | ( x91 & n498 ) ;
  assign n500 = n498 & ~n499 ;
  assign n501 = ( x91 & ~n499 ) | ( x91 & n500 ) | ( ~n499 & n500 ) ;
  assign n502 = ~x92 & n499 ;
  assign n503 = ( x73 & x92 ) | ( x73 & ~n499 ) | ( x92 & ~n499 ) ;
  assign n504 = ( ~x73 & n502 ) | ( ~x73 & n503 ) | ( n502 & n503 ) ;
  assign n505 = x4 & ~x6 ;
  assign n506 = ~x73 & n505 ;
  assign n507 = x94 & n506 ;
  assign n508 = x6 & ~x73 ;
  assign n509 = ( x4 & x73 ) | ( x4 & ~n508 ) | ( x73 & ~n508 ) ;
  assign n510 = ~n507 & n509 ;
  assign n511 = ( x93 & n507 ) | ( x93 & ~n510 ) | ( n507 & ~n510 ) ;
  assign n512 = x95 & n506 ;
  assign n513 = n509 & ~n512 ;
  assign n514 = ( x94 & n512 ) | ( x94 & ~n513 ) | ( n512 & ~n513 ) ;
  assign n515 = x96 & n506 ;
  assign n516 = n509 & ~n515 ;
  assign n517 = ( x95 & n515 ) | ( x95 & ~n516 ) | ( n515 & ~n516 ) ;
  assign n518 = x97 & n506 ;
  assign n519 = n509 & ~n518 ;
  assign n520 = ( x96 & n518 ) | ( x96 & ~n519 ) | ( n518 & ~n519 ) ;
  assign n521 = x98 & n506 ;
  assign n522 = n509 & ~n521 ;
  assign n523 = ( x97 & n521 ) | ( x97 & ~n522 ) | ( n521 & ~n522 ) ;
  assign n524 = x99 & n506 ;
  assign n525 = n509 & ~n524 ;
  assign n526 = ( x98 & n524 ) | ( x98 & ~n525 ) | ( n524 & ~n525 ) ;
  assign n527 = x100 & n506 ;
  assign n528 = n509 & ~n527 ;
  assign n529 = ( x99 & n527 ) | ( x99 & ~n528 ) | ( n527 & ~n528 ) ;
  assign n530 = x5 & n506 ;
  assign n531 = x100 | n530 ;
  assign n532 = ( ~n509 & n530 ) | ( ~n509 & n531 ) | ( n530 & n531 ) ;
  assign n533 = x4 & ~x73 ;
  assign n534 = x6 & n533 ;
  assign n535 = x102 & n534 ;
  assign n536 = x6 | x73 ;
  assign n537 = ( x4 & x73 ) | ( x4 & n536 ) | ( x73 & n536 ) ;
  assign n538 = ~n535 & n537 ;
  assign n539 = ( x101 & n535 ) | ( x101 & ~n538 ) | ( n535 & ~n538 ) ;
  assign n540 = x103 & n534 ;
  assign n541 = n537 & ~n540 ;
  assign n542 = ( x102 & n540 ) | ( x102 & ~n541 ) | ( n540 & ~n541 ) ;
  assign n543 = x104 & n534 ;
  assign n544 = n537 & ~n543 ;
  assign n545 = ( x103 & n543 ) | ( x103 & ~n544 ) | ( n543 & ~n544 ) ;
  assign n546 = x105 & n534 ;
  assign n547 = n537 & ~n546 ;
  assign n548 = ( x104 & n546 ) | ( x104 & ~n547 ) | ( n546 & ~n547 ) ;
  assign n549 = x106 & n534 ;
  assign n550 = n537 & ~n549 ;
  assign n551 = ( x105 & n549 ) | ( x105 & ~n550 ) | ( n549 & ~n550 ) ;
  assign n552 = x107 & n534 ;
  assign n553 = n537 & ~n552 ;
  assign n554 = ( x106 & n552 ) | ( x106 & ~n553 ) | ( n552 & ~n553 ) ;
  assign n555 = x108 & n534 ;
  assign n556 = n537 & ~n555 ;
  assign n557 = ( x107 & n555 ) | ( x107 & ~n556 ) | ( n555 & ~n556 ) ;
  assign n558 = x5 & n534 ;
  assign n559 = x108 | n558 ;
  assign n560 = ( ~n537 & n558 ) | ( ~n537 & n559 ) | ( n558 & n559 ) ;
  assign n561 = x2 & ~x3 ;
  assign n562 = ( ~x40 & x73 ) | ( ~x40 & n561 ) | ( x73 & n561 ) ;
  assign n563 = x3 & ~x56 ;
  assign n564 = ~x72 & n163 ;
  assign n565 = ~x1 & n564 ;
  assign n566 = ( x1 & n163 ) | ( x1 & ~n300 ) | ( n163 & ~n300 ) ;
  assign n567 = x109 & ~n566 ;
  assign n568 = x1 | n567 ;
  assign n569 = ( x93 & n567 ) | ( x93 & n568 ) | ( n567 & n568 ) ;
  assign n570 = x110 | n569 ;
  assign n571 = ( n565 & n569 ) | ( n565 & n570 ) | ( n569 & n570 ) ;
  assign n572 = ~x2 & n571 ;
  assign n573 = x3 | n572 ;
  assign n574 = ~n563 & n573 ;
  assign n575 = ~x73 & n574 ;
  assign n576 = ( n561 & ~n562 ) | ( n561 & n575 ) | ( ~n562 & n575 ) ;
  assign n577 = x1 & ~x2 ;
  assign n578 = ~x94 & n577 ;
  assign n579 = ~x2 & x111 ;
  assign n580 = n565 & n579 ;
  assign n581 = x2 & ~x41 ;
  assign n582 = x110 & ~n566 ;
  assign n583 = x2 | n582 ;
  assign n584 = ~n581 & n583 ;
  assign n585 = n580 | n584 ;
  assign n586 = ( n577 & ~n578 ) | ( n577 & n585 ) | ( ~n578 & n585 ) ;
  assign n587 = ( x3 & ~x73 ) | ( x3 & n586 ) | ( ~x73 & n586 ) ;
  assign n588 = ( x3 & ~x57 ) | ( x3 & x73 ) | ( ~x57 & x73 ) ;
  assign n589 = n587 & ~n588 ;
  assign n590 = ~x95 & n577 ;
  assign n591 = ~x2 & x112 ;
  assign n592 = n565 & n591 ;
  assign n593 = x2 & ~x42 ;
  assign n594 = x111 & ~n566 ;
  assign n595 = x2 | n594 ;
  assign n596 = ~n593 & n595 ;
  assign n597 = n592 | n596 ;
  assign n598 = ( n577 & ~n590 ) | ( n577 & n597 ) | ( ~n590 & n597 ) ;
  assign n599 = ( x3 & ~x73 ) | ( x3 & n598 ) | ( ~x73 & n598 ) ;
  assign n600 = ( x3 & ~x58 ) | ( x3 & x73 ) | ( ~x58 & x73 ) ;
  assign n601 = n599 & ~n600 ;
  assign n602 = x3 & ~x73 ;
  assign n603 = ~x59 & n602 ;
  assign n604 = x2 & ~x73 ;
  assign n605 = ( x3 & x43 ) | ( x3 & n604 ) | ( x43 & n604 ) ;
  assign n606 = ~x3 & n605 ;
  assign n607 = x2 | x73 ;
  assign n608 = x3 | n607 ;
  assign n609 = ( ~x113 & n565 ) | ( ~x113 & n608 ) | ( n565 & n608 ) ;
  assign n610 = x112 & ~n566 ;
  assign n611 = x1 | n610 ;
  assign n612 = ( x96 & n610 ) | ( x96 & n611 ) | ( n610 & n611 ) ;
  assign n613 = ~n608 & n612 ;
  assign n614 = ( n565 & ~n609 ) | ( n565 & n613 ) | ( ~n609 & n613 ) ;
  assign n615 = n606 | n614 ;
  assign n616 = ( n602 & ~n603 ) | ( n602 & n615 ) | ( ~n603 & n615 ) ;
  assign n617 = ~x60 & n602 ;
  assign n618 = ( x3 & x44 ) | ( x3 & n604 ) | ( x44 & n604 ) ;
  assign n619 = ~x3 & n618 ;
  assign n620 = ( ~x114 & n565 ) | ( ~x114 & n608 ) | ( n565 & n608 ) ;
  assign n621 = x113 & ~n566 ;
  assign n622 = x1 | n621 ;
  assign n623 = ( x97 & n621 ) | ( x97 & n622 ) | ( n621 & n622 ) ;
  assign n624 = ~n608 & n623 ;
  assign n625 = ( n565 & ~n620 ) | ( n565 & n624 ) | ( ~n620 & n624 ) ;
  assign n626 = n619 | n625 ;
  assign n627 = ( n602 & ~n617 ) | ( n602 & n626 ) | ( ~n617 & n626 ) ;
  assign n628 = ~x61 & n602 ;
  assign n629 = ( x3 & x45 ) | ( x3 & n604 ) | ( x45 & n604 ) ;
  assign n630 = ~x3 & n629 ;
  assign n631 = ( ~x115 & n565 ) | ( ~x115 & n608 ) | ( n565 & n608 ) ;
  assign n632 = x114 & ~n566 ;
  assign n633 = x1 | n632 ;
  assign n634 = ( x98 & n632 ) | ( x98 & n633 ) | ( n632 & n633 ) ;
  assign n635 = ~n608 & n634 ;
  assign n636 = ( n565 & ~n631 ) | ( n565 & n635 ) | ( ~n631 & n635 ) ;
  assign n637 = n630 | n636 ;
  assign n638 = ( n602 & ~n628 ) | ( n602 & n637 ) | ( ~n628 & n637 ) ;
  assign n639 = ~x62 & n602 ;
  assign n640 = ( x3 & x46 ) | ( x3 & n604 ) | ( x46 & n604 ) ;
  assign n641 = ~x3 & n640 ;
  assign n642 = ( ~x116 & n565 ) | ( ~x116 & n608 ) | ( n565 & n608 ) ;
  assign n643 = x115 & ~n566 ;
  assign n644 = x1 | n643 ;
  assign n645 = ( x99 & n643 ) | ( x99 & n644 ) | ( n643 & n644 ) ;
  assign n646 = ~n608 & n645 ;
  assign n647 = ( n565 & ~n642 ) | ( n565 & n646 ) | ( ~n642 & n646 ) ;
  assign n648 = n641 | n647 ;
  assign n649 = ( n602 & ~n639 ) | ( n602 & n648 ) | ( ~n639 & n648 ) ;
  assign n650 = ( ~x47 & x73 ) | ( ~x47 & n561 ) | ( x73 & n561 ) ;
  assign n651 = x3 & ~x63 ;
  assign n652 = x116 & ~n566 ;
  assign n653 = x1 | n652 ;
  assign n654 = ( x100 & n652 ) | ( x100 & n653 ) | ( n652 & n653 ) ;
  assign n655 = x117 | n654 ;
  assign n656 = ( n565 & n654 ) | ( n565 & n655 ) | ( n654 & n655 ) ;
  assign n657 = ~x2 & n656 ;
  assign n658 = x3 | n657 ;
  assign n659 = ~n651 & n658 ;
  assign n660 = ~x73 & n659 ;
  assign n661 = ( n561 & ~n650 ) | ( n561 & n660 ) | ( ~n650 & n660 ) ;
  assign n662 = ~x64 & n602 ;
  assign n663 = ( x3 & x48 ) | ( x3 & n604 ) | ( x48 & n604 ) ;
  assign n664 = ~x3 & n663 ;
  assign n665 = ( ~x118 & n565 ) | ( ~x118 & n608 ) | ( n565 & n608 ) ;
  assign n666 = x117 & ~n566 ;
  assign n667 = x1 | n666 ;
  assign n668 = ( x101 & n666 ) | ( x101 & n667 ) | ( n666 & n667 ) ;
  assign n669 = ~n608 & n668 ;
  assign n670 = ( n565 & ~n665 ) | ( n565 & n669 ) | ( ~n665 & n669 ) ;
  assign n671 = n664 | n670 ;
  assign n672 = ( n602 & ~n662 ) | ( n602 & n671 ) | ( ~n662 & n671 ) ;
  assign n673 = ~x102 & n577 ;
  assign n674 = ~x2 & x119 ;
  assign n675 = n565 & n674 ;
  assign n676 = x2 & ~x49 ;
  assign n677 = x118 & ~n566 ;
  assign n678 = x2 | n677 ;
  assign n679 = ~n676 & n678 ;
  assign n680 = n675 | n679 ;
  assign n681 = ( n577 & ~n673 ) | ( n577 & n680 ) | ( ~n673 & n680 ) ;
  assign n682 = ( x3 & ~x73 ) | ( x3 & n681 ) | ( ~x73 & n681 ) ;
  assign n683 = ( x3 & ~x65 ) | ( x3 & x73 ) | ( ~x65 & x73 ) ;
  assign n684 = n682 & ~n683 ;
  assign n685 = ( x3 & ~x66 ) | ( x3 & x73 ) | ( ~x66 & x73 ) ;
  assign n686 = x119 & ~n566 ;
  assign n687 = x1 | n686 ;
  assign n688 = ( x103 & n686 ) | ( x103 & n687 ) | ( n686 & n687 ) ;
  assign n689 = x120 | n688 ;
  assign n690 = ( n565 & n688 ) | ( n565 & n689 ) | ( n688 & n689 ) ;
  assign n691 = ( x2 & ~x3 ) | ( x2 & n690 ) | ( ~x3 & n690 ) ;
  assign n692 = ( x2 & x3 ) | ( x2 & ~x50 ) | ( x3 & ~x50 ) ;
  assign n693 = n691 & ~n692 ;
  assign n694 = ~x73 & n693 ;
  assign n695 = ( x3 & ~n685 ) | ( x3 & n694 ) | ( ~n685 & n694 ) ;
  assign n696 = ( x3 & ~x67 ) | ( x3 & x73 ) | ( ~x67 & x73 ) ;
  assign n697 = x120 & ~n566 ;
  assign n698 = x1 | n697 ;
  assign n699 = ( x104 & n697 ) | ( x104 & n698 ) | ( n697 & n698 ) ;
  assign n700 = x121 | n699 ;
  assign n701 = ( n565 & n699 ) | ( n565 & n700 ) | ( n699 & n700 ) ;
  assign n702 = ( x2 & ~x3 ) | ( x2 & n701 ) | ( ~x3 & n701 ) ;
  assign n703 = ( x2 & x3 ) | ( x2 & ~x51 ) | ( x3 & ~x51 ) ;
  assign n704 = n702 & ~n703 ;
  assign n705 = ~x73 & n704 ;
  assign n706 = ( x3 & ~n696 ) | ( x3 & n705 ) | ( ~n696 & n705 ) ;
  assign n707 = ( x3 & ~x68 ) | ( x3 & x73 ) | ( ~x68 & x73 ) ;
  assign n708 = x121 & ~n566 ;
  assign n709 = x1 | n708 ;
  assign n710 = ( x105 & n708 ) | ( x105 & n709 ) | ( n708 & n709 ) ;
  assign n711 = x122 | n710 ;
  assign n712 = ( n565 & n710 ) | ( n565 & n711 ) | ( n710 & n711 ) ;
  assign n713 = ( x2 & ~x3 ) | ( x2 & n712 ) | ( ~x3 & n712 ) ;
  assign n714 = ( x2 & x3 ) | ( x2 & ~x52 ) | ( x3 & ~x52 ) ;
  assign n715 = n713 & ~n714 ;
  assign n716 = ~x73 & n715 ;
  assign n717 = ( x3 & ~n707 ) | ( x3 & n716 ) | ( ~n707 & n716 ) ;
  assign n718 = ~x69 & n602 ;
  assign n719 = ( x3 & x53 ) | ( x3 & n604 ) | ( x53 & n604 ) ;
  assign n720 = ~x3 & n719 ;
  assign n721 = ( ~x123 & n565 ) | ( ~x123 & n608 ) | ( n565 & n608 ) ;
  assign n722 = x122 & ~n566 ;
  assign n723 = x1 | n722 ;
  assign n724 = ( x106 & n722 ) | ( x106 & n723 ) | ( n722 & n723 ) ;
  assign n725 = ~n608 & n724 ;
  assign n726 = ( n565 & ~n721 ) | ( n565 & n725 ) | ( ~n721 & n725 ) ;
  assign n727 = n720 | n726 ;
  assign n728 = ( n602 & ~n718 ) | ( n602 & n727 ) | ( ~n718 & n727 ) ;
  assign n729 = ~x70 & n602 ;
  assign n730 = ( x3 & x54 ) | ( x3 & n604 ) | ( x54 & n604 ) ;
  assign n731 = ~x3 & n730 ;
  assign n732 = ( ~x124 & n565 ) | ( ~x124 & n608 ) | ( n565 & n608 ) ;
  assign n733 = x123 & ~n566 ;
  assign n734 = x1 | n733 ;
  assign n735 = ( x107 & n733 ) | ( x107 & n734 ) | ( n733 & n734 ) ;
  assign n736 = ~n608 & n735 ;
  assign n737 = ( n565 & ~n732 ) | ( n565 & n736 ) | ( ~n732 & n736 ) ;
  assign n738 = n731 | n737 ;
  assign n739 = ( n602 & ~n729 ) | ( n602 & n738 ) | ( ~n729 & n738 ) ;
  assign n740 = x2 & ~x55 ;
  assign n741 = x124 & ~n566 ;
  assign n742 = x2 | n741 ;
  assign n743 = ~n740 & n742 ;
  assign n744 = x108 | n743 ;
  assign n745 = ( n577 & n743 ) | ( n577 & n744 ) | ( n743 & n744 ) ;
  assign n746 = ( x3 & ~x73 ) | ( x3 & n745 ) | ( ~x73 & n745 ) ;
  assign n747 = ( x3 & ~x71 ) | ( x3 & x73 ) | ( ~x71 & x73 ) ;
  assign n748 = n746 & ~n747 ;
  assign n749 = ( x125 & x126 ) | ( x125 & ~n354 ) | ( x126 & ~n354 ) ;
  assign n750 = ~x126 & n749 ;
  assign n751 = ( ~x125 & n749 ) | ( ~x125 & n750 ) | ( n749 & n750 ) ;
  assign n752 = ( x125 & x126 ) | ( x125 & n354 ) | ( x126 & n354 ) ;
  assign n753 = ~x127 & n752 ;
  assign n754 = ( x127 & n354 ) | ( x127 & ~n752 ) | ( n354 & ~n752 ) ;
  assign n755 = ( ~n354 & n753 ) | ( ~n354 & n754 ) | ( n753 & n754 ) ;
  assign n756 = x127 & ~n752 ;
  assign n757 = ( x127 & n354 ) | ( x127 & ~n756 ) | ( n354 & ~n756 ) ;
  assign n758 = x128 & n757 ;
  assign n759 = x125 & x127 ;
  assign n760 = ( x126 & n354 ) | ( x126 & n759 ) | ( n354 & n759 ) ;
  assign n761 = ~n354 & n760 ;
  assign n762 = ~x128 & n761 ;
  assign n763 = ( x128 & ~n758 ) | ( x128 & n762 ) | ( ~n758 & n762 ) ;
  assign n764 = x127 & x128 ;
  assign n765 = ( x125 & n354 ) | ( x125 & n764 ) | ( n354 & n764 ) ;
  assign n766 = x126 & ~n765 ;
  assign n767 = ( x126 & n354 ) | ( x126 & ~n766 ) | ( n354 & ~n766 ) ;
  assign n768 = x129 & n767 ;
  assign n769 = n334 & ~n354 ;
  assign n770 = x129 | n769 ;
  assign n771 = ~n768 & n770 ;
  assign n772 = ( x125 & n354 ) | ( x125 & n359 ) | ( n354 & n359 ) ;
  assign n773 = ~x130 & n772 ;
  assign n774 = ( x130 & n354 ) | ( x130 & ~n772 ) | ( n354 & ~n772 ) ;
  assign n775 = ( ~n354 & n773 ) | ( ~n354 & n774 ) | ( n773 & n774 ) ;
  assign n776 = ( x125 & n354 ) | ( x125 & n413 ) | ( n354 & n413 ) ;
  assign n777 = ~x131 & n776 ;
  assign n778 = ( x131 & n354 ) | ( x131 & ~n776 ) | ( n354 & ~n776 ) ;
  assign n779 = ( ~n354 & n777 ) | ( ~n354 & n778 ) | ( n777 & n778 ) ;
  assign n780 = x131 & ~n776 ;
  assign n781 = ( x131 & n354 ) | ( x131 & ~n780 ) | ( n354 & ~n780 ) ;
  assign n782 = x132 & n781 ;
  assign n783 = x131 & n413 ;
  assign n784 = x125 & n783 ;
  assign n785 = ~n354 & n784 ;
  assign n786 = x132 | n785 ;
  assign n787 = ~n782 & n786 ;
  assign n788 = x131 & x132 ;
  assign n789 = ( n354 & n413 ) | ( n354 & n788 ) | ( n413 & n788 ) ;
  assign n790 = x125 & ~n789 ;
  assign n791 = ( x125 & n354 ) | ( x125 & ~n790 ) | ( n354 & ~n790 ) ;
  assign n792 = x133 & n791 ;
  assign n793 = x132 & n784 ;
  assign n794 = ~n354 & n793 ;
  assign n795 = x133 | n794 ;
  assign n796 = ~n792 & n795 ;
  assign n797 = x81 & ~x82 ;
  assign n798 = ( ~x36 & x38 ) | ( ~x36 & x78 ) | ( x38 & x78 ) ;
  assign n799 = ~x38 & x134 ;
  assign n800 = ( x78 & ~n798 ) | ( x78 & n799 ) | ( ~n798 & n799 ) ;
  assign n801 = x0 & n800 ;
  assign n802 = ( ~x81 & n797 ) | ( ~x81 & n801 ) | ( n797 & n801 ) ;
  assign y0 = ~n136 ;
  assign y1 = n144 ;
  assign y2 = n184 ;
  assign y3 = n187 ;
  assign y4 = n194 ;
  assign y5 = n197 ;
  assign y6 = n200 ;
  assign y7 = n203 ;
  assign y8 = n206 ;
  assign y9 = n209 ;
  assign y10 = n212 ;
  assign y11 = n215 ;
  assign y12 = n222 ;
  assign y13 = n225 ;
  assign y14 = n228 ;
  assign y15 = n231 ;
  assign y16 = n234 ;
  assign y17 = n237 ;
  assign y18 = n240 ;
  assign y19 = n243 ;
  assign y20 = n250 ;
  assign y21 = n253 ;
  assign y22 = n256 ;
  assign y23 = n259 ;
  assign y24 = n262 ;
  assign y25 = n265 ;
  assign y26 = n268 ;
  assign y27 = n271 ;
  assign y28 = n278 ;
  assign y29 = n281 ;
  assign y30 = n284 ;
  assign y31 = n287 ;
  assign y32 = n290 ;
  assign y33 = n293 ;
  assign y34 = n296 ;
  assign y35 = n299 ;
  assign y36 = n302 ;
  assign y37 = n303 ;
  assign y38 = n326 ;
  assign y39 = n353 ;
  assign y40 = n365 ;
  assign y41 = n374 ;
  assign y42 = n379 ;
  assign y43 = n429 ;
  assign y44 = n434 ;
  assign y45 = n435 ;
  assign y46 = n380 ;
  assign y47 = n446 ;
  assign y48 = n460 ;
  assign y49 = n468 ;
  assign y50 = ~n471 ;
  assign y51 = n474 ;
  assign y52 = n481 ;
  assign y53 = n489 ;
  assign y54 = n496 ;
  assign y55 = n501 ;
  assign y56 = n504 ;
  assign y57 = n511 ;
  assign y58 = n514 ;
  assign y59 = n517 ;
  assign y60 = n520 ;
  assign y61 = n523 ;
  assign y62 = n526 ;
  assign y63 = n529 ;
  assign y64 = n532 ;
  assign y65 = n539 ;
  assign y66 = n542 ;
  assign y67 = n545 ;
  assign y68 = n548 ;
  assign y69 = n551 ;
  assign y70 = n554 ;
  assign y71 = n557 ;
  assign y72 = n560 ;
  assign y73 = n576 ;
  assign y74 = n589 ;
  assign y75 = n601 ;
  assign y76 = n616 ;
  assign y77 = n627 ;
  assign y78 = n638 ;
  assign y79 = n649 ;
  assign y80 = n661 ;
  assign y81 = n672 ;
  assign y82 = n684 ;
  assign y83 = n695 ;
  assign y84 = n706 ;
  assign y85 = n717 ;
  assign y86 = n728 ;
  assign y87 = n739 ;
  assign y88 = n748 ;
  assign y89 = ~n423 ;
  assign y90 = n751 ;
  assign y91 = n755 ;
  assign y92 = n763 ;
  assign y93 = n771 ;
  assign y94 = n775 ;
  assign y95 = n779 ;
  assign y96 = n787 ;
  assign y97 = n796 ;
  assign y98 = n802 ;
endmodule
