module top( N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 , N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 );
  input N1 , N101 , N106 , N111 , N116 , N121 , N126 , N13 , N130 , N135 , N138 , N143 , N146 , N149 , N152 , N153 , N156 , N159 , N165 , N17 , N171 , N177 , N183 , N189 , N195 , N201 , N207 , N210 , N219 , N228 , N237 , N246 , N255 , N259 , N26 , N260 , N261 , N267 , N268 , N29 , N36 , N42 , N51 , N55 , N59 , N68 , N72 , N73 , N74 , N75 , N8 , N80 , N85 , N86 , N87 , N88 , N89 , N90 , N91 , N96 ;
  output N388 , N389 , N390 , N391 , N418 , N419 , N420 , N421 , N422 , N423 , N446 , N447 , N448 , N449 , N450 , N767 , N768 , N850 , N863 , N864 , N865 , N866 , N874 , N878 , N879 , N880 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 ;
  assign n61 = N29 & N75 ;
  assign n62 = N42 & n61 ;
  assign n63 = N29 & N36 ;
  assign n64 = N80 & n63 ;
  assign n65 = N42 & n63 ;
  assign n66 = N85 & N86 ;
  assign n67 = N1 & N8 ;
  assign n68 = N13 & N17 ;
  assign n69 = n67 & n68 ;
  assign n70 = N1 & N26 ;
  assign n71 = n68 & n70 ;
  assign n72 = ~n65 & n71 ;
  assign n73 = N59 & N75 ;
  assign n74 = N80 & n73 ;
  assign n75 = N36 & N59 ;
  assign n76 = N80 & n75 ;
  assign n77 = N42 & n75 ;
  assign n78 = N87 | N88 ;
  assign n79 = N90 & n78 ;
  assign n80 = n65 & n71 ;
  assign n81 = N51 & n70 ;
  assign n82 = N13 & N55 ;
  assign n83 = n67 & n82 ;
  assign n84 = N29 & N68 ;
  assign n85 = n83 & n84 ;
  assign n86 = N59 & N68 ;
  assign n87 = N74 & n86 ;
  assign n88 = n83 & n87 ;
  assign n89 = N89 & n78 ;
  assign n90 = N130 | N96 ;
  assign n91 = N130 & N96 ;
  assign n92 = n90 & ~n91 ;
  assign n93 = N91 & n92 ;
  assign n94 = N91 | n92 ;
  assign n95 = ~n93 & n94 ;
  assign n96 = N121 | N135 ;
  assign n97 = N121 & N135 ;
  assign n98 = n96 & ~n97 ;
  assign n99 = N126 & ~n98 ;
  assign n100 = ~N126 & n98 ;
  assign n101 = n99 | n100 ;
  assign n102 = N101 & ~N106 ;
  assign n103 = ~N101 & N106 ;
  assign n104 = n102 | n103 ;
  assign n105 = N111 | N116 ;
  assign n106 = N111 & N116 ;
  assign n107 = n105 & ~n106 ;
  assign n108 = n104 | n107 ;
  assign n109 = n104 & n107 ;
  assign n110 = n108 & ~n109 ;
  assign n111 = n101 | n110 ;
  assign n112 = n101 & n110 ;
  assign n113 = n111 & ~n112 ;
  assign n114 = ~n95 & n113 ;
  assign n115 = n95 & ~n113 ;
  assign n116 = n114 | n115 ;
  assign n117 = N159 | N177 ;
  assign n118 = N159 & N177 ;
  assign n119 = n117 & ~n118 ;
  assign n120 = N130 & ~n119 ;
  assign n121 = ~N130 & n119 ;
  assign n122 = n120 | n121 ;
  assign n123 = N189 | N195 ;
  assign n124 = N189 & N195 ;
  assign n125 = n123 & ~n124 ;
  assign n126 = N207 & ~n125 ;
  assign n127 = ~N207 & n125 ;
  assign n128 = n126 | n127 ;
  assign n129 = ~N165 & N201 ;
  assign n130 = N165 & ~N201 ;
  assign n131 = n129 | n130 ;
  assign n132 = N171 & ~N183 ;
  assign n133 = ~N171 & N183 ;
  assign n134 = n132 | n133 ;
  assign n135 = n131 & ~n134 ;
  assign n136 = ~n131 & n134 ;
  assign n137 = n135 | n136 ;
  assign n138 = ~n128 & n137 ;
  assign n139 = n128 & ~n137 ;
  assign n140 = n138 | n139 ;
  assign n141 = n122 & ~n140 ;
  assign n142 = ~n122 & n140 ;
  assign n143 = n141 | n142 ;
  assign n144 = N156 & N59 ;
  assign n145 = n81 & ~n144 ;
  assign n146 = N17 & n145 ;
  assign n147 = N1 & ~n146 ;
  assign n148 = N153 & ~n147 ;
  assign n149 = N80 & n61 ;
  assign n150 = n81 & n149 ;
  assign n151 = N55 & n150 ;
  assign n152 = ~N268 & n151 ;
  assign n153 = N17 & ~N42 ;
  assign n154 = ~N17 & N42 ;
  assign n155 = n153 | n154 ;
  assign n156 = n81 & n144 ;
  assign n157 = n155 & n156 ;
  assign n158 = N42 & n73 ;
  assign n159 = N17 & N51 ;
  assign n160 = n67 & n159 ;
  assign n161 = ~n158 & n160 ;
  assign n162 = n157 | n161 ;
  assign n163 = N126 & n162 ;
  assign n164 = n152 | n163 ;
  assign n165 = n148 | n164 ;
  assign n166 = N201 | n165 ;
  assign n167 = N201 & n165 ;
  assign n168 = n166 & ~n167 ;
  assign n169 = N261 & n168 ;
  assign n170 = N261 | n168 ;
  assign n171 = N219 & n170 ;
  assign n172 = ~n169 & n171 ;
  assign n173 = N228 & n168 ;
  assign n174 = N237 & n167 ;
  assign n175 = N246 & n165 ;
  assign n176 = N42 & N72 ;
  assign n177 = N73 & n176 ;
  assign n178 = n86 & n177 ;
  assign n179 = n83 & n178 ;
  assign n180 = N201 & n179 ;
  assign n181 = N255 & N267 ;
  assign n182 = N121 & N210 ;
  assign n183 = n181 | n182 ;
  assign n184 = n180 | n183 ;
  assign n185 = n175 | n184 ;
  assign n186 = n174 | n185 ;
  assign n187 = n173 | n186 ;
  assign n188 = n172 | n187 ;
  assign n189 = N146 & ~n147 ;
  assign n190 = N116 & n162 ;
  assign n191 = n152 | n190 ;
  assign n192 = n189 | n191 ;
  assign n193 = N189 & n192 ;
  assign n194 = N189 | n192 ;
  assign n195 = N149 & ~n147 ;
  assign n196 = N121 & n162 ;
  assign n197 = n152 | n196 ;
  assign n198 = n195 | n197 ;
  assign n199 = N195 & n198 ;
  assign n200 = N195 | n198 ;
  assign n201 = N261 | n167 ;
  assign n202 = n166 & n201 ;
  assign n203 = n200 & n202 ;
  assign n204 = n199 | n203 ;
  assign n205 = n194 & n204 ;
  assign n206 = n193 | n205 ;
  assign n207 = N111 & n162 ;
  assign n208 = N143 & ~n147 ;
  assign n209 = n207 | n208 ;
  assign n210 = n152 | n209 ;
  assign n211 = N183 & n210 ;
  assign n212 = N183 | n210 ;
  assign n213 = ~n211 & n212 ;
  assign n214 = n206 | n213 ;
  assign n215 = n206 & n213 ;
  assign n216 = n214 & ~n215 ;
  assign n217 = N219 & n216 ;
  assign n218 = N228 & n213 ;
  assign n219 = N237 & n211 ;
  assign n220 = N246 & n210 ;
  assign n221 = N183 & n179 ;
  assign n222 = N106 & N210 ;
  assign n223 = n221 | n222 ;
  assign n224 = n220 | n223 ;
  assign n225 = n219 | n224 ;
  assign n226 = n218 | n225 ;
  assign n227 = n217 | n226 ;
  assign n228 = ~n193 & n194 ;
  assign n229 = n204 | n228 ;
  assign n230 = n204 & n228 ;
  assign n231 = n229 & ~n230 ;
  assign n232 = N219 & n231 ;
  assign n233 = N228 & n228 ;
  assign n234 = N237 & n193 ;
  assign n235 = N246 & n192 ;
  assign n236 = N189 & n179 ;
  assign n237 = N111 & N210 ;
  assign n238 = N255 & N259 ;
  assign n239 = n237 | n238 ;
  assign n240 = n236 | n239 ;
  assign n241 = n235 | n240 ;
  assign n242 = n234 | n241 ;
  assign n243 = n233 | n242 ;
  assign n244 = n232 | n243 ;
  assign n245 = ~n199 & n200 ;
  assign n246 = n202 | n245 ;
  assign n247 = n202 & n245 ;
  assign n248 = n246 & ~n247 ;
  assign n249 = N219 & n248 ;
  assign n250 = N228 & n245 ;
  assign n251 = N237 & n199 ;
  assign n252 = N246 & n198 ;
  assign n253 = N195 & n179 ;
  assign n254 = N255 & N260 ;
  assign n255 = N116 & N210 ;
  assign n256 = n254 | n255 ;
  assign n257 = n253 | n256 ;
  assign n258 = n252 | n257 ;
  assign n259 = n251 | n258 ;
  assign n260 = n250 | n259 ;
  assign n261 = n249 | n260 ;
  assign n262 = N91 & n162 ;
  assign n263 = N55 & n145 ;
  assign n264 = N143 & n263 ;
  assign n265 = N17 & ~N268 ;
  assign n266 = n150 & n265 ;
  assign n267 = N138 & N8 ;
  assign n268 = n266 | n267 ;
  assign n269 = n264 | n268 ;
  assign n270 = n262 | n269 ;
  assign n271 = N159 & n270 ;
  assign n272 = N159 | n270 ;
  assign n273 = N96 & n162 ;
  assign n274 = N146 & n263 ;
  assign n275 = N138 & N51 ;
  assign n276 = n266 | n275 ;
  assign n277 = n274 | n276 ;
  assign n278 = n273 | n277 ;
  assign n279 = N165 & n278 ;
  assign n280 = N165 | n278 ;
  assign n281 = N101 & n162 ;
  assign n282 = N149 & n263 ;
  assign n283 = N138 & N17 ;
  assign n284 = n266 | n283 ;
  assign n285 = n282 | n284 ;
  assign n286 = n281 | n285 ;
  assign n287 = N171 & n286 ;
  assign n288 = N171 | n286 ;
  assign n289 = N106 & n162 ;
  assign n290 = N153 & n263 ;
  assign n291 = N138 & N152 ;
  assign n292 = n266 | n291 ;
  assign n293 = n290 | n292 ;
  assign n294 = n289 | n293 ;
  assign n295 = N177 & n294 ;
  assign n296 = N177 | n294 ;
  assign n297 = n206 & n212 ;
  assign n298 = n211 | n297 ;
  assign n299 = n296 & n298 ;
  assign n300 = n295 | n299 ;
  assign n301 = n288 & n300 ;
  assign n302 = n287 | n301 ;
  assign n303 = n280 & n302 ;
  assign n304 = n279 | n303 ;
  assign n305 = n272 & n304 ;
  assign n306 = n271 | n305 ;
  assign n307 = ~n295 & n296 ;
  assign n308 = N219 & ~n298 ;
  assign n309 = N228 | n308 ;
  assign n310 = n307 & n309 ;
  assign n311 = N219 & ~n307 ;
  assign n312 = n298 & n311 ;
  assign n313 = N237 & n295 ;
  assign n314 = N246 & n294 ;
  assign n315 = N177 & n179 ;
  assign n316 = N101 & N210 ;
  assign n317 = n315 | n316 ;
  assign n318 = n314 | n317 ;
  assign n319 = n313 | n318 ;
  assign n320 = n312 | n319 ;
  assign n321 = n310 | n320 ;
  assign n322 = ~n271 & n272 ;
  assign n323 = n304 | n322 ;
  assign n324 = n304 & n322 ;
  assign n325 = N219 & ~n324 ;
  assign n326 = n323 & n325 ;
  assign n327 = N228 & n322 ;
  assign n328 = N237 & n271 ;
  assign n329 = N246 & n270 ;
  assign n330 = N159 & n179 ;
  assign n331 = N210 & N268 ;
  assign n332 = n330 | n331 ;
  assign n333 = n329 | n332 ;
  assign n334 = n328 | n333 ;
  assign n335 = n327 | n334 ;
  assign n336 = n326 | n335 ;
  assign n337 = ~n279 & n280 ;
  assign n338 = n302 & n337 ;
  assign n339 = n302 | n337 ;
  assign n340 = N219 & n339 ;
  assign n341 = ~n338 & n340 ;
  assign n342 = N228 & n337 ;
  assign n343 = N237 & n279 ;
  assign n344 = N246 & n278 ;
  assign n345 = N210 & N91 ;
  assign n346 = N165 & n179 ;
  assign n347 = n345 | n346 ;
  assign n348 = n344 | n347 ;
  assign n349 = n343 | n348 ;
  assign n350 = n342 | n349 ;
  assign n351 = n341 | n350 ;
  assign n352 = ~n287 & n288 ;
  assign n353 = n300 & n352 ;
  assign n354 = n300 | n352 ;
  assign n355 = N219 & n354 ;
  assign n356 = ~n353 & n355 ;
  assign n357 = N228 & n352 ;
  assign n358 = N237 & n287 ;
  assign n359 = N246 & n286 ;
  assign n360 = N210 & N96 ;
  assign n361 = N171 & n179 ;
  assign n362 = n360 | n361 ;
  assign n363 = n359 | n362 ;
  assign n364 = n358 | n363 ;
  assign n365 = n357 | n364 ;
  assign n366 = n356 | n365 ;
  assign N388 = n62 ;
  assign N389 = n64 ;
  assign N390 = n65 ;
  assign N391 = n66 ;
  assign N418 = n69 ;
  assign N419 = ~n72 ;
  assign N420 = ~n74 ;
  assign N421 = ~n76 ;
  assign N422 = ~n77 ;
  assign N423 = n79 ;
  assign N446 = ~n80 ;
  assign N447 = n81 ;
  assign N448 = n85 ;
  assign N449 = n88 ;
  assign N450 = n89 ;
  assign N767 = n116 ;
  assign N768 = n143 ;
  assign N850 = n188 ;
  assign N863 = n227 ;
  assign N864 = n244 ;
  assign N865 = n261 ;
  assign N866 = n306 ;
  assign N874 = n321 ;
  assign N878 = n336 ;
  assign N879 = n351 ;
  assign N880 = n366 ;
endmodule
