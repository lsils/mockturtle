module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 ;
  assign n42 = x18 | x19 ;
  assign n43 = x17 | n42 ;
  assign n44 = x16 | n43 ;
  assign n45 = ( x17 & x18 ) | ( x17 & ~x19 ) | ( x18 & ~x19 ) ;
  assign n46 = ( x15 & x19 ) | ( x15 & n45 ) | ( x19 & n45 ) ;
  assign n47 = ( x17 & x19 ) | ( x17 & ~n46 ) | ( x19 & ~n46 ) ;
  assign n48 = n45 | n47 ;
  assign n49 = ( x15 & ~n46 ) | ( x15 & n48 ) | ( ~n46 & n48 ) ;
  assign n50 = ~x16 & n49 ;
  assign n51 = ~x17 & x19 ;
  assign n52 = ( ~x17 & x18 ) | ( ~x17 & n51 ) | ( x18 & n51 ) ;
  assign n53 = x15 & n52 ;
  assign n54 = x16 & ~n53 ;
  assign n55 = n50 | n54 ;
  assign n56 = x13 & n55 ;
  assign n57 = ( n43 & ~n44 ) | ( n43 & n56 ) | ( ~n44 & n56 ) ;
  assign n58 = x12 & x40 ;
  assign n59 = ( x14 & n57 ) | ( x14 & n58 ) | ( n57 & n58 ) ;
  assign n60 = ~n57 & n59 ;
  assign n61 = ~x4 & n60 ;
  assign n62 = ( x3 & ~x5 ) | ( x3 & n61 ) | ( ~x5 & n61 ) ;
  assign n63 = ~x3 & n62 ;
  assign n64 = ( x15 & x17 ) | ( x15 & x19 ) | ( x17 & x19 ) ;
  assign n65 = ( x15 & x18 ) | ( x15 & ~n64 ) | ( x18 & ~n64 ) ;
  assign n66 = x18 & x19 ;
  assign n67 = ( x15 & n64 ) | ( x15 & n66 ) | ( n64 & n66 ) ;
  assign n68 = ( x19 & n65 ) | ( x19 & ~n67 ) | ( n65 & ~n67 ) ;
  assign n69 = ( ~x16 & x40 ) | ( ~x16 & n68 ) | ( x40 & n68 ) ;
  assign n70 = ~x18 & x19 ;
  assign n71 = x16 & x17 ;
  assign n72 = ( x18 & n70 ) | ( x18 & n71 ) | ( n70 & n71 ) ;
  assign n73 = ~x15 & n72 ;
  assign n74 = x40 & n73 ;
  assign n75 = ( ~n68 & n69 ) | ( ~n68 & n74 ) | ( n69 & n74 ) ;
  assign n76 = x15 | x16 ;
  assign n77 = x17 & ~n42 ;
  assign n78 = x5 & n77 ;
  assign n79 = ~n76 & n78 ;
  assign n80 = x5 & ~n79 ;
  assign n81 = ( n75 & n79 ) | ( n75 & ~n80 ) | ( n79 & ~n80 ) ;
  assign n82 = ( x3 & x13 ) | ( x3 & n81 ) | ( x13 & n81 ) ;
  assign n83 = x5 | x15 ;
  assign n84 = ~x16 & x17 ;
  assign n85 = ~n42 & n84 ;
  assign n86 = x3 & n85 ;
  assign n87 = ~n83 & n86 ;
  assign n88 = ~x13 & n87 ;
  assign n89 = ( n81 & ~n82 ) | ( n81 & n88 ) | ( ~n82 & n88 ) ;
  assign n90 = ~x4 & x12 ;
  assign n91 = ( x2 & n89 ) | ( x2 & n90 ) | ( n89 & n90 ) ;
  assign n92 = ~x2 & n91 ;
  assign n93 = ( x1 & ~x14 ) | ( x1 & n92 ) | ( ~x14 & n92 ) ;
  assign n94 = x15 & ~x16 ;
  assign n95 = x17 | x18 ;
  assign n96 = x17 & n66 ;
  assign n97 = ( ~x15 & n94 ) | ( ~x15 & n96 ) | ( n94 & n96 ) ;
  assign n98 = n95 & ~n97 ;
  assign n99 = ( x16 & n94 ) | ( x16 & ~n98 ) | ( n94 & ~n98 ) ;
  assign n100 = ~x12 & n99 ;
  assign n101 = ~x28 & x31 ;
  assign n102 = x24 & x25 ;
  assign n103 = x28 & ~n102 ;
  assign n104 = n101 | n103 ;
  assign n105 = ~x15 & n104 ;
  assign n106 = x12 & ~n105 ;
  assign n107 = n100 | n106 ;
  assign n108 = x40 & n107 ;
  assign n109 = x15 & ~n95 ;
  assign n110 = ~x15 & x16 ;
  assign n111 = n109 | n110 ;
  assign n112 = ( n96 & n109 ) | ( n96 & n111 ) | ( n109 & n111 ) ;
  assign n113 = ~x12 & n112 ;
  assign n114 = x4 & ~x5 ;
  assign n115 = ( x5 & ~n113 ) | ( x5 & n114 ) | ( ~n113 & n114 ) ;
  assign n116 = ( x5 & ~n108 ) | ( x5 & n114 ) | ( ~n108 & n114 ) ;
  assign n117 = ( n108 & ~n115 ) | ( n108 & n116 ) | ( ~n115 & n116 ) ;
  assign n118 = x2 & ~x3 ;
  assign n119 = ( x3 & ~n113 ) | ( x3 & n118 ) | ( ~n113 & n118 ) ;
  assign n120 = ( x3 & ~n117 ) | ( x3 & n118 ) | ( ~n117 & n118 ) ;
  assign n121 = ( n117 & ~n119 ) | ( n117 & n120 ) | ( ~n119 & n120 ) ;
  assign n122 = ( x1 & ~x13 ) | ( x1 & n121 ) | ( ~x13 & n121 ) ;
  assign n123 = x2 | x3 ;
  assign n124 = ~x4 & x15 ;
  assign n125 = ~n123 & n124 ;
  assign n126 = x16 & ~x17 ;
  assign n127 = n70 & n126 ;
  assign n128 = n125 & ~n127 ;
  assign n129 = x4 | x5 ;
  assign n130 = n94 & ~n129 ;
  assign n131 = ( n43 & ~n123 ) | ( n43 & n130 ) | ( ~n123 & n130 ) ;
  assign n132 = ~n43 & n131 ;
  assign n133 = x16 & ~x19 ;
  assign n134 = x16 | x19 ;
  assign n135 = ( ~x16 & n133 ) | ( ~x16 & n134 ) | ( n133 & n134 ) ;
  assign n136 = x15 & ~x17 ;
  assign n137 = ( x18 & n135 ) | ( x18 & ~n136 ) | ( n135 & ~n136 ) ;
  assign n138 = n135 & ~n137 ;
  assign n139 = n110 | n138 ;
  assign n140 = ( n96 & n138 ) | ( n96 & n139 ) | ( n138 & n139 ) ;
  assign n141 = n132 | n140 ;
  assign n142 = ( n125 & ~n128 ) | ( n125 & n141 ) | ( ~n128 & n141 ) ;
  assign n143 = x1 & n142 ;
  assign n144 = ~x12 & n143 ;
  assign n145 = x13 & n144 ;
  assign n146 = ( n121 & ~n122 ) | ( n121 & n145 ) | ( ~n122 & n145 ) ;
  assign n147 = ~x14 & n146 ;
  assign n148 = ( ~x1 & n93 ) | ( ~x1 & n147 ) | ( n93 & n147 ) ;
  assign n149 = ( x1 & x2 ) | ( x1 & ~n148 ) | ( x2 & ~n148 ) ;
  assign n150 = n63 & n149 ;
  assign n151 = ( n63 & n148 ) | ( n63 & ~n150 ) | ( n148 & ~n150 ) ;
  assign n152 = ( x0 & ~x36 ) | ( x0 & n151 ) | ( ~x36 & n151 ) ;
  assign n153 = x12 & ~x13 ;
  assign n154 = ~x5 & n153 ;
  assign n155 = x3 | x4 ;
  assign n156 = ~n76 & n77 ;
  assign n157 = ~n155 & n156 ;
  assign n158 = n154 & n157 ;
  assign n159 = x16 | x17 ;
  assign n160 = n70 & ~n159 ;
  assign n161 = ( x15 & ~x18 ) | ( x15 & x19 ) | ( ~x18 & x19 ) ;
  assign n162 = ( ~x17 & x19 ) | ( ~x17 & n161 ) | ( x19 & n161 ) ;
  assign n163 = x19 & ~n162 ;
  assign n164 = n162 | n163 ;
  assign n165 = ( ~x19 & n163 ) | ( ~x19 & n164 ) | ( n163 & n164 ) ;
  assign n166 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n167 = n165 & ~n166 ;
  assign n168 = x16 & n167 ;
  assign n169 = ~x5 & x15 ;
  assign n170 = ~n155 & n169 ;
  assign n171 = n168 | n170 ;
  assign n172 = ( n160 & n168 ) | ( n160 & n171 ) | ( n168 & n171 ) ;
  assign n173 = ( ~x12 & n158 ) | ( ~x12 & n172 ) | ( n158 & n172 ) ;
  assign n174 = x13 & ~n173 ;
  assign n175 = ( x13 & n158 ) | ( x13 & ~n174 ) | ( n158 & ~n174 ) ;
  assign n176 = x1 | x14 ;
  assign n177 = ( x2 & n175 ) | ( x2 & n176 ) | ( n175 & n176 ) ;
  assign n178 = n175 & ~n177 ;
  assign n179 = ( x0 & x36 ) | ( x0 & ~n178 ) | ( x36 & ~n178 ) ;
  assign n180 = n152 & ~n179 ;
  assign n181 = ~x10 & n180 ;
  assign n182 = ( x9 & ~x11 ) | ( x9 & n181 ) | ( ~x11 & n181 ) ;
  assign n183 = ~x9 & n182 ;
  assign n184 = ~x8 & n183 ;
  assign n185 = x15 | x17 ;
  assign n186 = ~x15 & n70 ;
  assign n187 = x17 & n186 ;
  assign n188 = ( ~x17 & n185 ) | ( ~x17 & n187 ) | ( n185 & n187 ) ;
  assign n189 = ( ~x14 & x16 ) | ( ~x14 & n188 ) | ( x16 & n188 ) ;
  assign n190 = ~x13 & x14 ;
  assign n191 = ( n188 & ~n189 ) | ( n188 & n190 ) | ( ~n189 & n190 ) ;
  assign n192 = x13 & ~x15 ;
  assign n193 = ( x14 & ~x28 ) | ( x14 & n192 ) | ( ~x28 & n192 ) ;
  assign n194 = ~x14 & n193 ;
  assign n195 = ~n191 & n194 ;
  assign n196 = ~x36 & x40 ;
  assign n197 = ( n191 & n195 ) | ( n191 & n196 ) | ( n195 & n196 ) ;
  assign n198 = ~x11 & x12 ;
  assign n199 = ( x10 & n197 ) | ( x10 & n198 ) | ( n197 & n198 ) ;
  assign n200 = ~x10 & n199 ;
  assign n201 = ~x8 & n200 ;
  assign n202 = ( x5 & ~x9 ) | ( x5 & n201 ) | ( ~x9 & n201 ) ;
  assign n203 = ~x5 & n202 ;
  assign n204 = ~x3 & n203 ;
  assign n205 = ( x2 & ~x4 ) | ( x2 & n204 ) | ( ~x4 & n204 ) ;
  assign n206 = ~x2 & n205 ;
  assign n207 = ~x0 & n206 ;
  assign n208 = ~x1 & n207 ;
  assign n209 = x15 & ~n159 ;
  assign n210 = ( ~x13 & x14 ) | ( ~x13 & n209 ) | ( x14 & n209 ) ;
  assign n211 = x14 & n210 ;
  assign n212 = ( x15 & x24 ) | ( x15 & x25 ) | ( x24 & x25 ) ;
  assign n213 = x28 & ~n212 ;
  assign n214 = ( x15 & x28 ) | ( x15 & ~n213 ) | ( x28 & ~n213 ) ;
  assign n215 = x13 & ~x14 ;
  assign n216 = ( n211 & ~n214 ) | ( n211 & n215 ) | ( ~n214 & n215 ) ;
  assign n217 = n211 | n216 ;
  assign n218 = ( x12 & n196 ) | ( x12 & ~n217 ) | ( n196 & ~n217 ) ;
  assign n219 = n217 & n218 ;
  assign n220 = ~x10 & n219 ;
  assign n221 = ( x9 & ~x11 ) | ( x9 & n220 ) | ( ~x11 & n220 ) ;
  assign n222 = ~x9 & n221 ;
  assign n223 = ~x5 & n222 ;
  assign n224 = ( x4 & ~x8 ) | ( x4 & n223 ) | ( ~x8 & n223 ) ;
  assign n225 = ~x4 & n224 ;
  assign n226 = ~x2 & n225 ;
  assign n227 = ( x1 & ~x3 ) | ( x1 & n226 ) | ( ~x3 & n226 ) ;
  assign n228 = ~x1 & n227 ;
  assign n229 = ~x0 & n228 ;
  assign n230 = ( x4 & ~n114 ) | ( x4 & n123 ) | ( ~n114 & n123 ) ;
  assign n231 = ~x14 & x16 ;
  assign n232 = ( x18 & n230 ) | ( x18 & ~n231 ) | ( n230 & ~n231 ) ;
  assign n233 = n230 & ~n232 ;
  assign n234 = ~x2 & x12 ;
  assign n235 = ~x3 & n234 ;
  assign n236 = x3 & ~x14 ;
  assign n237 = ( x2 & ~x14 ) | ( x2 & n236 ) | ( ~x14 & n236 ) ;
  assign n238 = x12 | n237 ;
  assign n239 = x14 & x40 ;
  assign n240 = ~n123 & n239 ;
  assign n241 = x12 & ~n240 ;
  assign n242 = n238 & ~n241 ;
  assign n243 = ~x18 & n242 ;
  assign n244 = x18 & x40 ;
  assign n245 = x14 & n244 ;
  assign n246 = n243 | n245 ;
  assign n247 = ( n235 & n243 ) | ( n235 & n246 ) | ( n243 & n246 ) ;
  assign n248 = x5 | n247 ;
  assign n249 = x14 | x18 ;
  assign n250 = ~x2 & x3 ;
  assign n251 = ( x2 & ~n249 ) | ( x2 & n250 ) | ( ~n249 & n250 ) ;
  assign n252 = ~x12 & n251 ;
  assign n253 = x5 & ~n252 ;
  assign n254 = n248 & ~n253 ;
  assign n255 = ( x4 & ~x16 ) | ( x4 & n254 ) | ( ~x16 & n254 ) ;
  assign n256 = ( x3 & x5 ) | ( x3 & ~x18 ) | ( x5 & ~x18 ) ;
  assign n257 = ~x2 & n256 ;
  assign n258 = ( x2 & ~x18 ) | ( x2 & n257 ) | ( ~x18 & n257 ) ;
  assign n259 = ~x12 & n258 ;
  assign n260 = ~x14 & n259 ;
  assign n261 = ( x4 & x16 ) | ( x4 & ~n260 ) | ( x16 & ~n260 ) ;
  assign n262 = n255 & ~n261 ;
  assign n263 = x12 & ~n262 ;
  assign n264 = ( n233 & n262 ) | ( n233 & ~n263 ) | ( n262 & ~n263 ) ;
  assign n265 = x1 | n264 ;
  assign n266 = x5 & x16 ;
  assign n267 = ( x5 & n249 ) | ( x5 & ~n266 ) | ( n249 & ~n266 ) ;
  assign n268 = x4 | n267 ;
  assign n269 = ( ~x3 & x12 ) | ( ~x3 & n268 ) | ( x12 & n268 ) ;
  assign n270 = x3 | n269 ;
  assign n271 = x2 | n270 ;
  assign n272 = x1 & n271 ;
  assign n273 = n265 & ~n272 ;
  assign n274 = ~x15 & n273 ;
  assign n275 = x3 | n129 ;
  assign n276 = x14 | x15 ;
  assign n277 = ~x18 & x40 ;
  assign n278 = x16 & n277 ;
  assign n279 = ( x12 & ~n276 ) | ( x12 & n278 ) | ( ~n276 & n278 ) ;
  assign n280 = ~x12 & n279 ;
  assign n281 = ~x2 & n280 ;
  assign n282 = ( x1 & ~n275 ) | ( x1 & n281 ) | ( ~n275 & n281 ) ;
  assign n283 = ~x1 & n282 ;
  assign n284 = x2 | x4 ;
  assign n285 = x3 | n284 ;
  assign n286 = x1 & ~n285 ;
  assign n287 = ~x4 & x40 ;
  assign n288 = ~x5 & n287 ;
  assign n289 = ~n123 & n288 ;
  assign n290 = x1 | n289 ;
  assign n291 = ~n286 & n290 ;
  assign n292 = ( x18 & ~n135 ) | ( x18 & n291 ) | ( ~n135 & n291 ) ;
  assign n293 = ( x4 & x5 ) | ( x4 & ~n135 ) | ( x5 & ~n135 ) ;
  assign n294 = ( x1 & x4 ) | ( x1 & x5 ) | ( x4 & x5 ) ;
  assign n295 = n293 & ~n294 ;
  assign n296 = ~x16 & x19 ;
  assign n297 = x1 & x5 ;
  assign n298 = ( x4 & n296 ) | ( x4 & n297 ) | ( n296 & n297 ) ;
  assign n299 = ~x4 & n298 ;
  assign n300 = ~n295 & n299 ;
  assign n301 = ( ~n123 & n295 ) | ( ~n123 & n300 ) | ( n295 & n300 ) ;
  assign n302 = ~x18 & n301 ;
  assign n303 = ( n291 & ~n292 ) | ( n291 & n302 ) | ( ~n292 & n302 ) ;
  assign n304 = ~x14 & x15 ;
  assign n305 = ( x12 & n303 ) | ( x12 & n304 ) | ( n303 & n304 ) ;
  assign n306 = ~x12 & n305 ;
  assign n307 = n283 | n306 ;
  assign n308 = ( n273 & ~n274 ) | ( n273 & n307 ) | ( ~n274 & n307 ) ;
  assign n309 = ~x17 & n308 ;
  assign n310 = x2 | x5 ;
  assign n311 = ( ~x1 & x3 ) | ( ~x1 & n310 ) | ( x3 & n310 ) ;
  assign n312 = x1 | n311 ;
  assign n313 = x17 & x19 ;
  assign n314 = ( x18 & ~n312 ) | ( x18 & n313 ) | ( ~n312 & n313 ) ;
  assign n315 = n312 & n314 ;
  assign n316 = ( x12 & n110 ) | ( x12 & n315 ) | ( n110 & n315 ) ;
  assign n317 = ~x12 & n316 ;
  assign n318 = x4 & n317 ;
  assign n319 = ( x2 & x3 ) | ( x2 & x19 ) | ( x3 & x19 ) ;
  assign n320 = ~x1 & n319 ;
  assign n321 = ( x1 & x19 ) | ( x1 & n320 ) | ( x19 & n320 ) ;
  assign n322 = x16 & x18 ;
  assign n323 = ( x17 & ~n321 ) | ( x17 & n322 ) | ( ~n321 & n322 ) ;
  assign n324 = n321 & n323 ;
  assign n325 = x5 & ~x15 ;
  assign n326 = ( x12 & n324 ) | ( x12 & n325 ) | ( n324 & n325 ) ;
  assign n327 = ~x12 & n326 ;
  assign n328 = ( x2 & x3 ) | ( x2 & x16 ) | ( x3 & x16 ) ;
  assign n329 = ~x40 & n328 ;
  assign n330 = ( x16 & x40 ) | ( x16 & n329 ) | ( x40 & n329 ) ;
  assign n331 = x15 | n330 ;
  assign n332 = ~x16 & x40 ;
  assign n333 = ~n123 & n332 ;
  assign n334 = x15 & ~n333 ;
  assign n335 = n331 & ~n334 ;
  assign n336 = ( x18 & n313 ) | ( x18 & ~n335 ) | ( n313 & ~n335 ) ;
  assign n337 = n335 & n336 ;
  assign n338 = ~x12 & n337 ;
  assign n339 = x15 & ~x29 ;
  assign n340 = x25 & x28 ;
  assign n341 = x27 & n340 ;
  assign n342 = x24 & n341 ;
  assign n343 = x15 | n342 ;
  assign n344 = ~n339 & n343 ;
  assign n345 = ~x3 & x40 ;
  assign n346 = ( x12 & ~n344 ) | ( x12 & n345 ) | ( ~n344 & n345 ) ;
  assign n347 = n344 & n346 ;
  assign n348 = n338 | n347 ;
  assign n349 = ( ~x2 & n338 ) | ( ~x2 & n348 ) | ( n338 & n348 ) ;
  assign n350 = ( x1 & ~x5 ) | ( x1 & n349 ) | ( ~x5 & n349 ) ;
  assign n351 = ( x12 & n96 ) | ( x12 & n110 ) | ( n96 & n110 ) ;
  assign n352 = ~x12 & n351 ;
  assign n353 = ( x1 & x5 ) | ( x1 & ~n352 ) | ( x5 & ~n352 ) ;
  assign n354 = n350 & ~n353 ;
  assign n355 = n327 | n354 ;
  assign n356 = ~x4 & n355 ;
  assign n357 = n318 | n356 ;
  assign n358 = n309 | n357 ;
  assign n359 = ( ~x14 & n309 ) | ( ~x14 & n358 ) | ( n309 & n358 ) ;
  assign n360 = x0 | n359 ;
  assign n361 = x2 | x14 ;
  assign n362 = ( x12 & n172 ) | ( x12 & n361 ) | ( n172 & n361 ) ;
  assign n363 = n172 & ~n362 ;
  assign n364 = ~x1 & n363 ;
  assign n365 = x0 & ~n364 ;
  assign n366 = n360 & ~n365 ;
  assign n367 = x13 & n366 ;
  assign n368 = ( x15 & x16 ) | ( x15 & ~x18 ) | ( x16 & ~x18 ) ;
  assign n369 = ~x16 & x18 ;
  assign n370 = ( x15 & x40 ) | ( x15 & ~n369 ) | ( x40 & ~n369 ) ;
  assign n371 = ~n368 & n370 ;
  assign n372 = x3 | n371 ;
  assign n373 = x16 | x18 ;
  assign n374 = x15 | n373 ;
  assign n375 = x3 & n374 ;
  assign n376 = n372 & ~n375 ;
  assign n377 = x0 | n376 ;
  assign n378 = x3 | n374 ;
  assign n379 = x0 & n378 ;
  assign n380 = n377 & ~n379 ;
  assign n381 = x17 & n380 ;
  assign n382 = ~x19 & n381 ;
  assign n383 = x12 & ~x14 ;
  assign n384 = ( x13 & n382 ) | ( x13 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ~x13 & n384 ;
  assign n386 = ~x4 & n385 ;
  assign n387 = ( x2 & ~x5 ) | ( x2 & n386 ) | ( ~x5 & n386 ) ;
  assign n388 = ~x2 & n387 ;
  assign n389 = n367 | n388 ;
  assign n390 = ( ~x1 & n367 ) | ( ~x1 & n389 ) | ( n367 & n389 ) ;
  assign n391 = x10 | x36 ;
  assign n392 = ( x11 & n390 ) | ( x11 & n391 ) | ( n390 & n391 ) ;
  assign n393 = n390 & ~n392 ;
  assign n394 = ~x8 & n393 ;
  assign n395 = ~x9 & n394 ;
  assign n396 = ~x17 & x40 ;
  assign n397 = x14 & n396 ;
  assign n398 = ( x15 & x16 ) | ( x15 & n397 ) | ( x16 & n397 ) ;
  assign n399 = ~x16 & n398 ;
  assign n400 = x13 & n399 ;
  assign n401 = ( x5 & x12 ) | ( x5 & n400 ) | ( x12 & n400 ) ;
  assign n402 = ~x5 & n401 ;
  assign n403 = ~x3 & n402 ;
  assign n404 = ( x2 & ~x4 ) | ( x2 & n403 ) | ( ~x4 & n403 ) ;
  assign n405 = ~x2 & n404 ;
  assign n406 = x1 | x12 ;
  assign n407 = ( x2 & n172 ) | ( x2 & n406 ) | ( n172 & n406 ) ;
  assign n408 = n172 & ~n407 ;
  assign n409 = x0 & n408 ;
  assign n410 = x15 & x29 ;
  assign n411 = ( x24 & x27 ) | ( x24 & n340 ) | ( x27 & n340 ) ;
  assign n412 = ~x27 & n411 ;
  assign n413 = ~x15 & n412 ;
  assign n414 = ( x15 & ~n410 ) | ( x15 & n413 ) | ( ~n410 & n413 ) ;
  assign n415 = ( x12 & ~x40 ) | ( x12 & n414 ) | ( ~x40 & n414 ) ;
  assign n416 = ~x17 & x18 ;
  assign n417 = ( x15 & x16 ) | ( x15 & n416 ) | ( x16 & n416 ) ;
  assign n418 = x17 & ~x18 ;
  assign n419 = ( x15 & x16 ) | ( x15 & ~n418 ) | ( x16 & ~n418 ) ;
  assign n420 = ~n417 & n419 ;
  assign n421 = x16 & ~n43 ;
  assign n422 = x19 | n421 ;
  assign n423 = ( n420 & n421 ) | ( n420 & n422 ) | ( n421 & n422 ) ;
  assign n424 = ( x12 & x40 ) | ( x12 & n423 ) | ( x40 & n423 ) ;
  assign n425 = ~n415 & n424 ;
  assign n426 = ( x3 & n118 ) | ( x3 & ~n425 ) | ( n118 & ~n425 ) ;
  assign n427 = ( ~n119 & n425 ) | ( ~n119 & n426 ) | ( n425 & n426 ) ;
  assign n428 = x5 | n427 ;
  assign n429 = ( x2 & x16 ) | ( x2 & x19 ) | ( x16 & x19 ) ;
  assign n430 = ( x18 & n134 ) | ( x18 & ~n429 ) | ( n134 & ~n429 ) ;
  assign n431 = x17 | n430 ;
  assign n432 = x15 & ~n431 ;
  assign n433 = ( n96 & n110 ) | ( n96 & n432 ) | ( n110 & n432 ) ;
  assign n434 = x2 & ~n433 ;
  assign n435 = ( x2 & n432 ) | ( x2 & ~n434 ) | ( n432 & ~n434 ) ;
  assign n436 = ( ~x2 & n140 ) | ( ~x2 & n435 ) | ( n140 & n435 ) ;
  assign n437 = x3 & ~n436 ;
  assign n438 = ( x3 & n435 ) | ( x3 & ~n437 ) | ( n435 & ~n437 ) ;
  assign n439 = ~x12 & n438 ;
  assign n440 = x5 & ~n439 ;
  assign n441 = n428 & ~n440 ;
  assign n442 = ( ~x1 & x4 ) | ( ~x1 & n441 ) | ( x4 & n441 ) ;
  assign n443 = ~x2 & x5 ;
  assign n444 = ( x3 & n140 ) | ( x3 & ~n443 ) | ( n140 & ~n443 ) ;
  assign n445 = n140 & ~n444 ;
  assign n446 = ~x12 & n445 ;
  assign n447 = ( ~x12 & n438 ) | ( ~x12 & n446 ) | ( n438 & n446 ) ;
  assign n448 = ( x1 & x4 ) | ( x1 & ~n447 ) | ( x4 & ~n447 ) ;
  assign n449 = n442 & ~n448 ;
  assign n450 = n144 | n449 ;
  assign n451 = ~x0 & n450 ;
  assign n452 = n409 | n451 ;
  assign n453 = ( ~x13 & x14 ) | ( ~x13 & n452 ) | ( x14 & n452 ) ;
  assign n454 = ~x13 & n382 ;
  assign n455 = ( x5 & x12 ) | ( x5 & n454 ) | ( x12 & n454 ) ;
  assign n456 = ~x5 & n455 ;
  assign n457 = ~x2 & n456 ;
  assign n458 = ( x1 & ~x4 ) | ( x1 & n457 ) | ( ~x4 & n457 ) ;
  assign n459 = ~x1 & n458 ;
  assign n460 = ~x14 & n459 ;
  assign n461 = ( n452 & ~n453 ) | ( n452 & n460 ) | ( ~n453 & n460 ) ;
  assign n462 = ( x0 & x1 ) | ( x0 & ~n461 ) | ( x1 & ~n461 ) ;
  assign n463 = n405 & n462 ;
  assign n464 = ( n405 & n461 ) | ( n405 & ~n463 ) | ( n461 & ~n463 ) ;
  assign n465 = ( x11 & n391 ) | ( x11 & n464 ) | ( n391 & n464 ) ;
  assign n466 = n464 & ~n465 ;
  assign n467 = ~x8 & n466 ;
  assign n468 = ~x9 & n467 ;
  assign n469 = x5 & x15 ;
  assign n470 = x16 & ~x40 ;
  assign n471 = ( x5 & x16 ) | ( x5 & ~n470 ) | ( x16 & ~n470 ) ;
  assign n472 = ( x5 & x15 ) | ( x5 & n471 ) | ( x15 & n471 ) ;
  assign n473 = ( n469 & n471 ) | ( n469 & ~n472 ) | ( n471 & ~n472 ) ;
  assign n474 = x17 | x19 ;
  assign n475 = ( x18 & n473 ) | ( x18 & n474 ) | ( n473 & n474 ) ;
  assign n476 = n473 & ~n475 ;
  assign n477 = x17 & x18 ;
  assign n478 = n109 | n477 ;
  assign n479 = ( n109 & n110 ) | ( n109 & n478 ) | ( n110 & n478 ) ;
  assign n480 = ( ~x5 & x19 ) | ( ~x5 & n479 ) | ( x19 & n479 ) ;
  assign n481 = ( x40 & ~n94 ) | ( x40 & n477 ) | ( ~n94 & n477 ) ;
  assign n482 = ~n95 & n110 ;
  assign n483 = x40 & n482 ;
  assign n484 = ( n94 & n481 ) | ( n94 & n483 ) | ( n481 & n483 ) ;
  assign n485 = ( x5 & x19 ) | ( x5 & n484 ) | ( x19 & n484 ) ;
  assign n486 = n480 & n485 ;
  assign n487 = ~x5 & x40 ;
  assign n488 = ( x12 & n414 ) | ( x12 & n487 ) | ( n414 & n487 ) ;
  assign n489 = ~n414 & n488 ;
  assign n490 = ( ~n476 & n486 ) | ( ~n476 & n489 ) | ( n486 & n489 ) ;
  assign n491 = x12 & ~n489 ;
  assign n492 = ( n476 & n490 ) | ( n476 & ~n491 ) | ( n490 & ~n491 ) ;
  assign n493 = x3 & ~x4 ;
  assign n494 = ( x4 & ~n113 ) | ( x4 & n493 ) | ( ~n113 & n493 ) ;
  assign n495 = ( x4 & ~n492 ) | ( x4 & n493 ) | ( ~n492 & n493 ) ;
  assign n496 = ( n492 & ~n494 ) | ( n492 & n495 ) | ( ~n494 & n495 ) ;
  assign n497 = ( ~x1 & x2 ) | ( ~x1 & n496 ) | ( x2 & n496 ) ;
  assign n498 = ( x1 & x2 ) | ( x1 & ~n113 ) | ( x2 & ~n113 ) ;
  assign n499 = n497 & ~n498 ;
  assign n500 = ~x5 & n165 ;
  assign n501 = ( ~x4 & n165 ) | ( ~x4 & n500 ) | ( n165 & n500 ) ;
  assign n502 = ( x4 & n160 ) | ( x4 & n169 ) | ( n160 & n169 ) ;
  assign n503 = ~x4 & n502 ;
  assign n504 = x16 | n503 ;
  assign n505 = ( n501 & n503 ) | ( n501 & n504 ) | ( n503 & n504 ) ;
  assign n506 = x2 | x12 ;
  assign n507 = ( x3 & n505 ) | ( x3 & n506 ) | ( n505 & n506 ) ;
  assign n508 = n505 & ~n507 ;
  assign n509 = ~x1 & n508 ;
  assign n510 = x0 & n509 ;
  assign n511 = ( ~n144 & n499 ) | ( ~n144 & n510 ) | ( n499 & n510 ) ;
  assign n512 = x0 & ~n510 ;
  assign n513 = ( n144 & n511 ) | ( n144 & ~n512 ) | ( n511 & ~n512 ) ;
  assign n514 = ~x14 & n513 ;
  assign n515 = ~x5 & x12 ;
  assign n516 = ( x4 & n399 ) | ( x4 & n515 ) | ( n399 & n515 ) ;
  assign n517 = ~x4 & n516 ;
  assign n518 = ~x2 & n517 ;
  assign n519 = ( x1 & ~x3 ) | ( x1 & n518 ) | ( ~x3 & n518 ) ;
  assign n520 = ~x1 & n519 ;
  assign n521 = n514 | n520 ;
  assign n522 = ( ~x0 & n514 ) | ( ~x0 & n521 ) | ( n514 & n521 ) ;
  assign n523 = x13 & n522 ;
  assign n524 = ( x15 & x16 ) | ( x15 & x18 ) | ( x16 & x18 ) ;
  assign n525 = ( x15 & x16 ) | ( x15 & ~x40 ) | ( x16 & ~x40 ) ;
  assign n526 = n524 & ~n525 ;
  assign n527 = x5 | n526 ;
  assign n528 = x5 & n374 ;
  assign n529 = n527 & ~n528 ;
  assign n530 = ~x14 & x17 ;
  assign n531 = ( x19 & n529 ) | ( x19 & ~n530 ) | ( n529 & ~n530 ) ;
  assign n532 = n529 & ~n531 ;
  assign n533 = ~x13 & n532 ;
  assign n534 = ( x4 & x12 ) | ( x4 & n533 ) | ( x12 & n533 ) ;
  assign n535 = ~x4 & n534 ;
  assign n536 = ~x2 & n535 ;
  assign n537 = ( x1 & ~x3 ) | ( x1 & n536 ) | ( ~x3 & n536 ) ;
  assign n538 = ~x1 & n537 ;
  assign n539 = n523 | n538 ;
  assign n540 = ( ~x0 & n523 ) | ( ~x0 & n539 ) | ( n523 & n539 ) ;
  assign n541 = ( x11 & n391 ) | ( x11 & n540 ) | ( n391 & n540 ) ;
  assign n542 = n540 & ~n541 ;
  assign n543 = ~x8 & n542 ;
  assign n544 = ~x9 & n543 ;
  assign n545 = ( ~x17 & n42 ) | ( ~x17 & n110 ) | ( n42 & n110 ) ;
  assign n546 = x15 & n369 ;
  assign n547 = ~x17 & n546 ;
  assign n548 = ( ~n42 & n545 ) | ( ~n42 & n547 ) | ( n545 & n547 ) ;
  assign n549 = ( ~x12 & x13 ) | ( ~x12 & n548 ) | ( x13 & n548 ) ;
  assign n550 = x13 & n549 ;
  assign n551 = ( x15 & n153 ) | ( x15 & n550 ) | ( n153 & n550 ) ;
  assign n552 = n550 | n551 ;
  assign n553 = ( x14 & n487 ) | ( x14 & ~n552 ) | ( n487 & ~n552 ) ;
  assign n554 = n552 & n553 ;
  assign n555 = ~x3 & n554 ;
  assign n556 = ( x2 & ~x4 ) | ( x2 & n555 ) | ( ~x4 & n555 ) ;
  assign n557 = ~x2 & n556 ;
  assign n558 = x12 & x13 ;
  assign n559 = x13 & ~n558 ;
  assign n560 = n109 & n559 ;
  assign n561 = x22 & x23 ;
  assign n562 = ~x20 & x21 ;
  assign n563 = ( ~x24 & n561 ) | ( ~x24 & n562 ) | ( n561 & n562 ) ;
  assign n564 = ~n561 & n563 ;
  assign n565 = x21 & ~n564 ;
  assign n566 = ( x20 & n564 ) | ( x20 & ~n565 ) | ( n564 & ~n565 ) ;
  assign n567 = x27 & n566 ;
  assign n568 = ~x19 & n567 ;
  assign n569 = x18 & n568 ;
  assign n570 = ~x15 & x17 ;
  assign n571 = n569 & n570 ;
  assign n572 = ( ~n558 & n559 ) | ( ~n558 & n571 ) | ( n559 & n571 ) ;
  assign n573 = ( x12 & n560 ) | ( x12 & n572 ) | ( n560 & n572 ) ;
  assign n574 = n109 | n570 ;
  assign n575 = ( n66 & n109 ) | ( n66 & n574 ) | ( n109 & n574 ) ;
  assign n576 = ~x12 & x16 ;
  assign n577 = ( x13 & ~n575 ) | ( x13 & n576 ) | ( ~n575 & n576 ) ;
  assign n578 = n575 & n577 ;
  assign n579 = x16 & ~n578 ;
  assign n580 = ( n573 & n578 ) | ( n573 & ~n579 ) | ( n578 & ~n579 ) ;
  assign n581 = x4 & n580 ;
  assign n582 = ( x15 & x17 ) | ( x15 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n583 = ~x17 & n582 ;
  assign n584 = ( ~x15 & x16 ) | ( ~x15 & n583 ) | ( x16 & n583 ) ;
  assign n585 = ( n582 & n583 ) | ( n582 & n584 ) | ( n583 & n584 ) ;
  assign n586 = n559 & n585 ;
  assign n587 = ( x22 & ~x23 ) | ( x22 & x24 ) | ( ~x23 & x24 ) ;
  assign n588 = x23 & n587 ;
  assign n589 = x24 & ~x26 ;
  assign n590 = ( x22 & ~n587 ) | ( x22 & n589 ) | ( ~n587 & n589 ) ;
  assign n591 = ( x24 & ~n588 ) | ( x24 & n590 ) | ( ~n588 & n590 ) ;
  assign n592 = ~x20 & x27 ;
  assign n593 = ( x21 & ~n591 ) | ( x21 & n592 ) | ( ~n591 & n592 ) ;
  assign n594 = n591 & n593 ;
  assign n595 = n566 | n594 ;
  assign n596 = x18 & n595 ;
  assign n597 = ( x15 & n84 ) | ( x15 & n596 ) | ( n84 & n596 ) ;
  assign n598 = ~x15 & n597 ;
  assign n599 = ( ~n558 & n559 ) | ( ~n558 & n598 ) | ( n559 & n598 ) ;
  assign n600 = ( x12 & n586 ) | ( x12 & n599 ) | ( n586 & n599 ) ;
  assign n601 = x5 | x40 ;
  assign n602 = ( x19 & n600 ) | ( x19 & ~n601 ) | ( n600 & ~n601 ) ;
  assign n603 = ~x12 & x19 ;
  assign n604 = ( x13 & ~n479 ) | ( x13 & n603 ) | ( ~n479 & n603 ) ;
  assign n605 = n479 & n604 ;
  assign n606 = n601 & n605 ;
  assign n607 = ( n600 & ~n602 ) | ( n600 & n606 ) | ( ~n602 & n606 ) ;
  assign n608 = x13 | x15 ;
  assign n609 = x12 & ~n608 ;
  assign n610 = ( x5 & ~n85 ) | ( x5 & n609 ) | ( ~n85 & n609 ) ;
  assign n611 = n85 & n610 ;
  assign n612 = ~x30 & x31 ;
  assign n613 = x32 & x33 ;
  assign n614 = x30 & ~n613 ;
  assign n615 = n612 | n614 ;
  assign n616 = x13 & ~n615 ;
  assign n617 = ( x15 & x16 ) | ( x15 & ~x19 ) | ( x16 & ~x19 ) ;
  assign n618 = x38 & x39 ;
  assign n619 = ( x15 & n617 ) | ( x15 & n618 ) | ( n617 & n618 ) ;
  assign n620 = n617 & n619 ;
  assign n621 = n76 & ~n620 ;
  assign n622 = x17 & n621 ;
  assign n623 = ~x18 & n622 ;
  assign n624 = x24 & ~x27 ;
  assign n625 = x22 | n624 ;
  assign n626 = ( x22 & x23 ) | ( x22 & ~n624 ) | ( x23 & ~n624 ) ;
  assign n627 = ( x23 & ~x24 ) | ( x23 & x26 ) | ( ~x24 & x26 ) ;
  assign n628 = x23 & ~x27 ;
  assign n629 = ( x24 & n627 ) | ( x24 & n628 ) | ( n627 & n628 ) ;
  assign n630 = x22 & n629 ;
  assign n631 = ( n625 & ~n626 ) | ( n625 & n630 ) | ( ~n626 & n630 ) ;
  assign n632 = x21 & n631 ;
  assign n633 = ~x20 & n632 ;
  assign n634 = x17 & n633 ;
  assign n635 = x15 & x16 ;
  assign n636 = ( x15 & n110 ) | ( x15 & ~n635 ) | ( n110 & ~n635 ) ;
  assign n637 = ( n634 & ~n635 ) | ( n634 & n636 ) | ( ~n635 & n636 ) ;
  assign n638 = ( ~x18 & x19 ) | ( ~x18 & n637 ) | ( x19 & n637 ) ;
  assign n639 = n51 & n94 ;
  assign n640 = x18 & n639 ;
  assign n641 = ( n637 & ~n638 ) | ( n637 & n640 ) | ( ~n638 & n640 ) ;
  assign n642 = n623 | n641 ;
  assign n643 = ~x13 & n642 ;
  assign n644 = n616 | n643 ;
  assign n645 = x12 & ~n644 ;
  assign n646 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n647 = ~n45 & n646 ;
  assign n648 = ( ~x15 & n482 ) | ( ~x15 & n647 ) | ( n482 & n647 ) ;
  assign n649 = ( x15 & n84 ) | ( x15 & n482 ) | ( n84 & n482 ) ;
  assign n650 = n648 | n649 ;
  assign n651 = x13 & n650 ;
  assign n652 = x12 | n651 ;
  assign n653 = ~n645 & n652 ;
  assign n654 = ( ~x5 & n611 ) | ( ~x5 & n653 ) | ( n611 & n653 ) ;
  assign n655 = x40 & ~n654 ;
  assign n656 = ( x40 & n611 ) | ( x40 & ~n655 ) | ( n611 & ~n655 ) ;
  assign n657 = n607 | n656 ;
  assign n658 = ~x4 & n657 ;
  assign n659 = n581 | n658 ;
  assign n660 = x13 & n112 ;
  assign n661 = ~x12 & n660 ;
  assign n662 = ( x3 & n118 ) | ( x3 & ~n661 ) | ( n118 & ~n661 ) ;
  assign n663 = ( x3 & n118 ) | ( x3 & ~n659 ) | ( n118 & ~n659 ) ;
  assign n664 = ( n659 & ~n662 ) | ( n659 & n663 ) | ( ~n662 & n663 ) ;
  assign n665 = ~x12 & x13 ;
  assign n666 = ( x1 & ~n142 ) | ( x1 & n665 ) | ( ~n142 & n665 ) ;
  assign n667 = n142 & n666 ;
  assign n668 = x1 & ~n667 ;
  assign n669 = ( n664 & n667 ) | ( n664 & ~n668 ) | ( n667 & ~n668 ) ;
  assign n670 = ( x0 & ~x14 ) | ( x0 & n669 ) | ( ~x14 & n669 ) ;
  assign n671 = n153 & n156 ;
  assign n672 = ~n129 & n671 ;
  assign n673 = ( ~x12 & n505 ) | ( ~x12 & n672 ) | ( n505 & n672 ) ;
  assign n674 = x13 & ~n673 ;
  assign n675 = ( x13 & n672 ) | ( x13 & ~n674 ) | ( n672 & ~n674 ) ;
  assign n676 = x1 | x3 ;
  assign n677 = ( x2 & n675 ) | ( x2 & n676 ) | ( n675 & n676 ) ;
  assign n678 = n675 & ~n677 ;
  assign n679 = ( x0 & x14 ) | ( x0 & ~n678 ) | ( x14 & ~n678 ) ;
  assign n680 = n670 & ~n679 ;
  assign n681 = ( x0 & x1 ) | ( x0 & ~n680 ) | ( x1 & ~n680 ) ;
  assign n682 = n557 & n681 ;
  assign n683 = ( n557 & n680 ) | ( n557 & ~n682 ) | ( n680 & ~n682 ) ;
  assign n684 = ( x11 & n391 ) | ( x11 & n683 ) | ( n391 & n683 ) ;
  assign n685 = n683 & ~n684 ;
  assign n686 = ~x8 & n685 ;
  assign n687 = ~x9 & n686 ;
  assign n688 = x19 | n618 ;
  assign n689 = x18 | n688 ;
  assign n690 = x17 & ~n689 ;
  assign n691 = ( x15 & x16 ) | ( x15 & n690 ) | ( x16 & n690 ) ;
  assign n692 = ~x15 & n691 ;
  assign n693 = x38 | x39 ;
  assign n694 = x37 | n693 ;
  assign n695 = x18 & ~n694 ;
  assign n696 = n665 & n695 ;
  assign n697 = n94 & n696 ;
  assign n698 = x15 & ~x18 ;
  assign n699 = x16 | n694 ;
  assign n700 = x15 & n699 ;
  assign n701 = ( n322 & n698 ) | ( n322 & ~n700 ) | ( n698 & ~n700 ) ;
  assign n702 = ( ~x13 & n697 ) | ( ~x13 & n701 ) | ( n697 & n701 ) ;
  assign n703 = x12 & ~n702 ;
  assign n704 = ( x12 & n697 ) | ( x12 & ~n703 ) | ( n697 & ~n703 ) ;
  assign n705 = ( x17 & x19 ) | ( x17 & n704 ) | ( x19 & n704 ) ;
  assign n706 = n94 & n665 ;
  assign n707 = ( n66 & n694 ) | ( n66 & n706 ) | ( n694 & n706 ) ;
  assign n708 = ~n694 & n707 ;
  assign n709 = ~x17 & n708 ;
  assign n710 = ( n704 & ~n705 ) | ( n704 & n709 ) | ( ~n705 & n709 ) ;
  assign n711 = ( x12 & ~x13 ) | ( x12 & n710 ) | ( ~x13 & n710 ) ;
  assign n712 = n692 & ~n711 ;
  assign n713 = ( n692 & n710 ) | ( n692 & ~n712 ) | ( n710 & ~n712 ) ;
  assign n714 = ~x14 & x40 ;
  assign n715 = ( x36 & n713 ) | ( x36 & ~n714 ) | ( n713 & ~n714 ) ;
  assign n716 = n713 & ~n715 ;
  assign n717 = ~x10 & n716 ;
  assign n718 = ( x9 & ~x11 ) | ( x9 & n717 ) | ( ~x11 & n717 ) ;
  assign n719 = ~x9 & n718 ;
  assign n720 = ~x4 & n719 ;
  assign n721 = ( x3 & ~x5 ) | ( x3 & n720 ) | ( ~x5 & n720 ) ;
  assign n722 = ~x3 & n721 ;
  assign n723 = ~x1 & n722 ;
  assign n724 = ( x0 & ~x2 ) | ( x0 & n723 ) | ( ~x2 & n723 ) ;
  assign n725 = ~x0 & n724 ;
  assign n726 = x9 & x11 ;
  assign n727 = ( x9 & ~x10 ) | ( x9 & n726 ) | ( ~x10 & n726 ) ;
  assign n728 = ~x8 & n727 ;
  assign n729 = ( ~x8 & n725 ) | ( ~x8 & n728 ) | ( n725 & n728 ) ;
  assign n730 = ~x14 & x30 ;
  assign n731 = ~x16 & n416 ;
  assign n732 = x15 & n731 ;
  assign n733 = x14 & ~n732 ;
  assign n734 = n730 | n733 ;
  assign n735 = ( x12 & x13 ) | ( x12 & n734 ) | ( x13 & n734 ) ;
  assign n736 = x18 | n618 ;
  assign n737 = x17 & ~n736 ;
  assign n738 = ( ~x17 & n95 ) | ( ~x17 & n737 ) | ( n95 & n737 ) ;
  assign n739 = ( x19 & ~n110 ) | ( x19 & n738 ) | ( ~n110 & n738 ) ;
  assign n740 = n738 & ~n739 ;
  assign n741 = ~x13 & n740 ;
  assign n742 = ~x14 & n741 ;
  assign n743 = x12 & n742 ;
  assign n744 = ( ~n734 & n735 ) | ( ~n734 & n743 ) | ( n735 & n743 ) ;
  assign n745 = x14 & ~x15 ;
  assign n746 = n744 | n745 ;
  assign n747 = ( n665 & n744 ) | ( n665 & n746 ) | ( n744 & n746 ) ;
  assign n748 = ~x11 & x40 ;
  assign n749 = ( x36 & n747 ) | ( x36 & ~n748 ) | ( n747 & ~n748 ) ;
  assign n750 = n747 & ~n749 ;
  assign n751 = ~x9 & n750 ;
  assign n752 = ( x8 & ~x10 ) | ( x8 & n751 ) | ( ~x10 & n751 ) ;
  assign n753 = ~x8 & n752 ;
  assign n754 = ~x4 & n753 ;
  assign n755 = ( x3 & ~x5 ) | ( x3 & n754 ) | ( ~x5 & n754 ) ;
  assign n756 = ~x3 & n755 ;
  assign n757 = ~x1 & n756 ;
  assign n758 = ( x0 & ~x2 ) | ( x0 & n757 ) | ( ~x2 & n757 ) ;
  assign n759 = ~x0 & n758 ;
  assign n760 = ( x14 & x30 ) | ( x14 & x32 ) | ( x30 & x32 ) ;
  assign n761 = x33 & ~n760 ;
  assign n762 = ( x14 & x33 ) | ( x14 & ~n761 ) | ( x33 & ~n761 ) ;
  assign n763 = x12 & ~n762 ;
  assign n764 = x12 | n231 ;
  assign n765 = ~n763 & n764 ;
  assign n766 = ~x15 & n765 ;
  assign n767 = ~x14 & n762 ;
  assign n768 = ( ~n731 & n762 ) | ( ~n731 & n767 ) | ( n762 & n767 ) ;
  assign n769 = x12 & ~n768 ;
  assign n770 = x15 & ~n769 ;
  assign n771 = n766 | n770 ;
  assign n772 = x13 | n743 ;
  assign n773 = ( n743 & ~n771 ) | ( n743 & n772 ) | ( ~n771 & n772 ) ;
  assign n774 = ( x36 & ~n748 ) | ( x36 & n773 ) | ( ~n748 & n773 ) ;
  assign n775 = n773 & ~n774 ;
  assign n776 = ~x9 & n775 ;
  assign n777 = ( x8 & ~x10 ) | ( x8 & n776 ) | ( ~x10 & n776 ) ;
  assign n778 = ~x8 & n777 ;
  assign n779 = ~x4 & n778 ;
  assign n780 = ( x3 & ~x5 ) | ( x3 & n779 ) | ( ~x5 & n779 ) ;
  assign n781 = ~x3 & n780 ;
  assign n782 = ~x1 & n781 ;
  assign n783 = ( x0 & ~x2 ) | ( x0 & n782 ) | ( ~x2 & n782 ) ;
  assign n784 = ~x0 & n783 ;
  assign n785 = ( x15 & n84 ) | ( x15 & n569 ) | ( n84 & n569 ) ;
  assign n786 = ~x15 & n785 ;
  assign n787 = ( x13 & n383 ) | ( x13 & n786 ) | ( n383 & n786 ) ;
  assign n788 = ~x13 & n787 ;
  assign n789 = ( x0 & ~x4 ) | ( x0 & n788 ) | ( ~x4 & n788 ) ;
  assign n790 = ( ~x12 & x14 ) | ( ~x12 & x18 ) | ( x14 & x18 ) ;
  assign n791 = x12 & ~n790 ;
  assign n792 = ( x14 & ~n695 ) | ( x14 & n790 ) | ( ~n695 & n790 ) ;
  assign n793 = ~x12 & n792 ;
  assign n794 = n791 | n793 ;
  assign n795 = ( x16 & x17 ) | ( x16 & ~n794 ) | ( x17 & ~n794 ) ;
  assign n796 = x12 | x14 ;
  assign n797 = x16 & ~x18 ;
  assign n798 = ~n796 & n797 ;
  assign n799 = ~x17 & n798 ;
  assign n800 = ( n794 & n795 ) | ( n794 & ~n799 ) | ( n795 & ~n799 ) ;
  assign n801 = x30 & x32 ;
  assign n802 = ( x33 & x35 ) | ( x33 & n801 ) | ( x35 & n801 ) ;
  assign n803 = ~x35 & n802 ;
  assign n804 = ( x14 & n800 ) | ( x14 & n803 ) | ( n800 & n803 ) ;
  assign n805 = x12 & n804 ;
  assign n806 = ( ~x12 & n800 ) | ( ~x12 & n805 ) | ( n800 & n805 ) ;
  assign n807 = x15 & n806 ;
  assign n808 = x12 & n803 ;
  assign n809 = x16 & n96 ;
  assign n810 = x12 | n809 ;
  assign n811 = ~n808 & n810 ;
  assign n812 = ~x14 & n811 ;
  assign n813 = x15 | n812 ;
  assign n814 = ~n807 & n813 ;
  assign n815 = ( x13 & x40 ) | ( x13 & ~n814 ) | ( x40 & ~n814 ) ;
  assign n816 = ( x16 & ~x17 ) | ( x16 & x19 ) | ( ~x17 & x19 ) ;
  assign n817 = x19 & ~n816 ;
  assign n818 = ( x17 & n694 ) | ( x17 & ~n817 ) | ( n694 & ~n817 ) ;
  assign n819 = ( n816 & ~n817 ) | ( n816 & n818 ) | ( ~n817 & n818 ) ;
  assign n820 = ( x15 & ~x18 ) | ( x15 & n819 ) | ( ~x18 & n819 ) ;
  assign n821 = x19 & n110 ;
  assign n822 = x17 & n821 ;
  assign n823 = ~x18 & n822 ;
  assign n824 = ( ~n819 & n820 ) | ( ~n819 & n823 ) | ( n820 & n823 ) ;
  assign n825 = ( x13 & n383 ) | ( x13 & n824 ) | ( n383 & n824 ) ;
  assign n826 = ~x13 & n825 ;
  assign n827 = x40 & n826 ;
  assign n828 = ( n814 & n815 ) | ( n814 & n827 ) | ( n815 & n827 ) ;
  assign n829 = ( ~x4 & x5 ) | ( ~x4 & n828 ) | ( x5 & n828 ) ;
  assign n830 = ( x19 & n665 ) | ( x19 & ~n797 ) | ( n665 & ~n797 ) ;
  assign n831 = x12 & ~x16 ;
  assign n832 = ( x13 & n596 ) | ( x13 & n831 ) | ( n596 & n831 ) ;
  assign n833 = ~x13 & n832 ;
  assign n834 = ~x19 & n833 ;
  assign n835 = ( n665 & ~n830 ) | ( n665 & n834 ) | ( ~n830 & n834 ) ;
  assign n836 = ( x14 & n570 ) | ( x14 & n835 ) | ( n570 & n835 ) ;
  assign n837 = ~x14 & n836 ;
  assign n838 = ( x4 & x5 ) | ( x4 & ~n837 ) | ( x5 & ~n837 ) ;
  assign n839 = n829 & ~n838 ;
  assign n840 = ~x0 & n839 ;
  assign n841 = ( n788 & ~n789 ) | ( n788 & n840 ) | ( ~n789 & n840 ) ;
  assign n842 = ~x4 & n154 ;
  assign n843 = x0 & n842 ;
  assign n844 = n77 & n843 ;
  assign n845 = ( x14 & ~n76 ) | ( x14 & n844 ) | ( ~n76 & n844 ) ;
  assign n846 = ~x14 & n845 ;
  assign n847 = ~n841 & n846 ;
  assign n848 = x11 | x36 ;
  assign n849 = ( n841 & n847 ) | ( n841 & ~n848 ) | ( n847 & ~n848 ) ;
  assign n850 = ~x9 & n849 ;
  assign n851 = ( x3 & ~x10 ) | ( x3 & n850 ) | ( ~x10 & n850 ) ;
  assign n852 = ~x3 & n851 ;
  assign n853 = ( x1 & x2 ) | ( x1 & ~n727 ) | ( x2 & ~n727 ) ;
  assign n854 = n852 & n853 ;
  assign n855 = ( n727 & n852 ) | ( n727 & ~n854 ) | ( n852 & ~n854 ) ;
  assign n856 = ~x8 & n855 ;
  assign n857 = ~x5 & n788 ;
  assign n858 = x4 & n857 ;
  assign n859 = ( n839 & n846 ) | ( n839 & ~n858 ) | ( n846 & ~n858 ) ;
  assign n860 = x0 & ~n846 ;
  assign n861 = ( n858 & n859 ) | ( n858 & ~n860 ) | ( n859 & ~n860 ) ;
  assign n862 = ( x11 & n391 ) | ( x11 & n861 ) | ( n391 & n861 ) ;
  assign n863 = n861 & ~n862 ;
  assign n864 = ~x8 & n863 ;
  assign n865 = ( x3 & ~x9 ) | ( x3 & n864 ) | ( ~x9 & n864 ) ;
  assign n866 = ~x3 & n865 ;
  assign n867 = ~x1 & n866 ;
  assign n868 = ~x2 & n867 ;
  assign n869 = ( x36 & n156 ) | ( x36 & ~n843 ) | ( n156 & ~n843 ) ;
  assign n870 = ~x19 & n595 ;
  assign n871 = x18 & n870 ;
  assign n872 = x17 & n871 ;
  assign n873 = ~x15 & n872 ;
  assign n874 = ( x13 & ~x16 ) | ( x13 & n873 ) | ( ~x16 & n873 ) ;
  assign n875 = ~x13 & n874 ;
  assign n876 = x5 & ~n875 ;
  assign n877 = x13 & ~n803 ;
  assign n878 = x18 & ~x19 ;
  assign n879 = ~x17 & n110 ;
  assign n880 = n878 & n879 ;
  assign n881 = n623 | n880 ;
  assign n882 = ~x13 & n881 ;
  assign n883 = n877 | n882 ;
  assign n884 = x40 & n883 ;
  assign n885 = x5 | n884 ;
  assign n886 = ~n876 & n885 ;
  assign n887 = x12 & ~n886 ;
  assign n888 = x40 & n575 ;
  assign n889 = x5 | n888 ;
  assign n890 = ~x15 & n77 ;
  assign n891 = x5 & ~n890 ;
  assign n892 = n889 & ~n891 ;
  assign n893 = x16 & n892 ;
  assign n894 = ( x16 & n136 ) | ( x16 & n277 ) | ( n136 & n277 ) ;
  assign n895 = ~x16 & n894 ;
  assign n896 = n893 | n895 ;
  assign n897 = ( ~x5 & n893 ) | ( ~x5 & n896 ) | ( n893 & n896 ) ;
  assign n898 = x13 & n897 ;
  assign n899 = x12 | n898 ;
  assign n900 = ~n887 & n899 ;
  assign n901 = ( ~x0 & x4 ) | ( ~x0 & n900 ) | ( x4 & n900 ) ;
  assign n902 = x5 & n786 ;
  assign n903 = ( x12 & x13 ) | ( x12 & n902 ) | ( x13 & n902 ) ;
  assign n904 = ~x13 & n903 ;
  assign n905 = ( x0 & x4 ) | ( x0 & ~n904 ) | ( x4 & ~n904 ) ;
  assign n906 = n901 & ~n905 ;
  assign n907 = ~x36 & n906 ;
  assign n908 = ( n156 & ~n869 ) | ( n156 & n907 ) | ( ~n869 & n907 ) ;
  assign n909 = ~x11 & n908 ;
  assign n910 = ( x10 & ~x14 ) | ( x10 & n909 ) | ( ~x14 & n909 ) ;
  assign n911 = ~x10 & n910 ;
  assign n912 = ~x3 & n911 ;
  assign n913 = ( x2 & ~x9 ) | ( x2 & n912 ) | ( ~x9 & n912 ) ;
  assign n914 = ~x2 & n913 ;
  assign n915 = ( x1 & ~x8 ) | ( x1 & n914 ) | ( ~x8 & n914 ) ;
  assign n916 = ( ~x1 & n728 ) | ( ~x1 & n915 ) | ( n728 & n915 ) ;
  assign n917 = x5 | n564 ;
  assign n918 = x20 & ~x21 ;
  assign n919 = x5 & ~n918 ;
  assign n920 = n917 & ~n919 ;
  assign n921 = ~x19 & x27 ;
  assign n922 = ( x18 & ~n920 ) | ( x18 & n921 ) | ( ~n920 & n921 ) ;
  assign n923 = n920 & n922 ;
  assign n924 = ( x15 & n84 ) | ( x15 & n923 ) | ( n84 & n923 ) ;
  assign n925 = ~x15 & n924 ;
  assign n926 = ( x13 & n383 ) | ( x13 & n925 ) | ( n383 & n925 ) ;
  assign n927 = ~x13 & n926 ;
  assign n928 = x2 & ~x4 ;
  assign n929 = ( x3 & n927 ) | ( x3 & n928 ) | ( n927 & n928 ) ;
  assign n930 = ~x3 & n929 ;
  assign n931 = ~x15 & x40 ;
  assign n932 = ( x5 & x16 ) | ( x5 & n931 ) | ( x16 & n931 ) ;
  assign n933 = ~x5 & n932 ;
  assign n934 = ~x4 & n933 ;
  assign n935 = x1 | n934 ;
  assign n936 = ( x4 & x5 ) | ( x4 & ~x16 ) | ( x5 & ~x16 ) ;
  assign n937 = ( x4 & ~x19 ) | ( x4 & n936 ) | ( ~x19 & n936 ) ;
  assign n938 = x4 & ~n937 ;
  assign n939 = n937 | n938 ;
  assign n940 = ( ~x4 & n938 ) | ( ~x4 & n939 ) | ( n938 & n939 ) ;
  assign n941 = x15 & n940 ;
  assign n942 = x1 & ~n941 ;
  assign n943 = n935 & ~n942 ;
  assign n944 = ( x17 & x18 ) | ( x17 & n943 ) | ( x18 & n943 ) ;
  assign n945 = ( x5 & n110 ) | ( x5 & n244 ) | ( n110 & n244 ) ;
  assign n946 = ~x5 & n945 ;
  assign n947 = ~x1 & n946 ;
  assign n948 = ~x4 & n947 ;
  assign n949 = ~x17 & n948 ;
  assign n950 = ( n943 & ~n944 ) | ( n943 & n949 ) | ( ~n944 & n949 ) ;
  assign n951 = ( x40 & n94 ) | ( x40 & ~n96 ) | ( n94 & ~n96 ) ;
  assign n952 = ( ~x18 & n42 ) | ( ~x18 & n878 ) | ( n42 & n878 ) ;
  assign n953 = x17 & n952 ;
  assign n954 = x16 & n953 ;
  assign n955 = ( x15 & n76 ) | ( x15 & ~n954 ) | ( n76 & ~n954 ) ;
  assign n956 = x40 & ~n955 ;
  assign n957 = ( n96 & n951 ) | ( n96 & n956 ) | ( n951 & n956 ) ;
  assign n958 = x5 | n957 ;
  assign n959 = n77 & n110 ;
  assign n960 = x5 & ~n959 ;
  assign n961 = n958 & ~n960 ;
  assign n962 = ( ~x1 & n950 ) | ( ~x1 & n961 ) | ( n950 & n961 ) ;
  assign n963 = x4 | n962 ;
  assign n964 = ( ~x4 & n950 ) | ( ~x4 & n963 ) | ( n950 & n963 ) ;
  assign n965 = ( x12 & ~x13 ) | ( x12 & n964 ) | ( ~x13 & n964 ) ;
  assign n966 = ( ~x15 & n58 ) | ( ~x15 & n94 ) | ( n58 & n94 ) ;
  assign n967 = ~x4 & n966 ;
  assign n968 = ( x1 & ~x5 ) | ( x1 & n967 ) | ( ~x5 & n967 ) ;
  assign n969 = ~x1 & n968 ;
  assign n970 = x13 & n969 ;
  assign n971 = ( n964 & ~n965 ) | ( n964 & n970 ) | ( ~n965 & n970 ) ;
  assign n972 = x20 & x21 ;
  assign n973 = ~x19 & n972 ;
  assign n974 = ( x4 & n570 ) | ( x4 & n973 ) | ( n570 & n973 ) ;
  assign n975 = ~x4 & n974 ;
  assign n976 = ( x4 & n51 ) | ( x4 & n975 ) | ( n51 & n975 ) ;
  assign n977 = x15 & ~n976 ;
  assign n978 = ( x15 & n975 ) | ( x15 & ~n977 ) | ( n975 & ~n977 ) ;
  assign n979 = x5 & ~n978 ;
  assign n980 = ( x15 & x19 ) | ( x15 & ~x40 ) | ( x19 & ~x40 ) ;
  assign n981 = ( x15 & ~x17 ) | ( x15 & x40 ) | ( ~x17 & x40 ) ;
  assign n982 = ~n980 & n981 ;
  assign n983 = ( x19 & ~n980 ) | ( x19 & n982 ) | ( ~n980 & n982 ) ;
  assign n984 = ~x4 & n983 ;
  assign n985 = x5 | n984 ;
  assign n986 = ~n979 & n985 ;
  assign n987 = x18 & n986 ;
  assign n988 = ~x38 & x39 ;
  assign n989 = x37 & n988 ;
  assign n990 = ( x15 & n64 ) | ( x15 & ~n989 ) | ( n64 & ~n989 ) ;
  assign n991 = n64 & n990 ;
  assign n992 = n185 & ~n991 ;
  assign n993 = ( ~x18 & n487 ) | ( ~x18 & n992 ) | ( n487 & n992 ) ;
  assign n994 = ~n992 & n993 ;
  assign n995 = n987 | n994 ;
  assign n996 = ( ~x4 & n987 ) | ( ~x4 & n995 ) | ( n987 & n995 ) ;
  assign n997 = ( x13 & x16 ) | ( x13 & n996 ) | ( x16 & n996 ) ;
  assign n998 = ~x19 & n618 ;
  assign n999 = x17 & n998 ;
  assign n1000 = ( ~x17 & n474 ) | ( ~x17 & n999 ) | ( n474 & n999 ) ;
  assign n1001 = x18 & n1000 ;
  assign n1002 = x16 & x40 ;
  assign n1003 = ( ~n1000 & n1001 ) | ( ~n1000 & n1002 ) | ( n1001 & n1002 ) ;
  assign n1004 = ~x5 & n1003 ;
  assign n1005 = ( x4 & ~x15 ) | ( x4 & n1004 ) | ( ~x15 & n1004 ) ;
  assign n1006 = ~x4 & n1005 ;
  assign n1007 = ~x13 & n1006 ;
  assign n1008 = ( n996 & ~n997 ) | ( n996 & n1007 ) | ( ~n997 & n1007 ) ;
  assign n1009 = ( ~x1 & n971 ) | ( ~x1 & n1008 ) | ( n971 & n1008 ) ;
  assign n1010 = x12 & ~n1009 ;
  assign n1011 = ( x12 & n971 ) | ( x12 & ~n1010 ) | ( n971 & ~n1010 ) ;
  assign n1012 = ~x14 & n1011 ;
  assign n1013 = ( ~x16 & x17 ) | ( ~x16 & n51 ) | ( x17 & n51 ) ;
  assign n1014 = ( x15 & ~x16 ) | ( x15 & n51 ) | ( ~x16 & n51 ) ;
  assign n1015 = ( n136 & n1013 ) | ( n136 & ~n1014 ) | ( n1013 & ~n1014 ) ;
  assign n1016 = x17 & n70 ;
  assign n1017 = ~n76 & n1016 ;
  assign n1018 = x18 | n1017 ;
  assign n1019 = ( n1015 & n1017 ) | ( n1015 & n1018 ) | ( n1017 & n1018 ) ;
  assign n1020 = ( x16 & x18 ) | ( x16 & x19 ) | ( x18 & x19 ) ;
  assign n1021 = x17 | n1020 ;
  assign n1022 = x13 & n1021 ;
  assign n1023 = ~n1019 & n1022 ;
  assign n1024 = ( x12 & ~x40 ) | ( x12 & n1023 ) | ( ~x40 & n1023 ) ;
  assign n1025 = ~x13 & x15 ;
  assign n1026 = ( x13 & n731 ) | ( x13 & ~n1025 ) | ( n731 & ~n1025 ) ;
  assign n1027 = ( x12 & x40 ) | ( x12 & n1026 ) | ( x40 & n1026 ) ;
  assign n1028 = ~n1024 & n1027 ;
  assign n1029 = ~x5 & x14 ;
  assign n1030 = ( x4 & n1028 ) | ( x4 & n1029 ) | ( n1028 & n1029 ) ;
  assign n1031 = ~x4 & n1030 ;
  assign n1032 = n1012 | n1031 ;
  assign n1033 = ( ~x1 & n1012 ) | ( ~x1 & n1032 ) | ( n1012 & n1032 ) ;
  assign n1034 = x3 | n1033 ;
  assign n1035 = ~x4 & x5 ;
  assign n1036 = x23 & ~x25 ;
  assign n1037 = ( ~x23 & n624 ) | ( ~x23 & n1036 ) | ( n624 & n1036 ) ;
  assign n1038 = x22 & n1037 ;
  assign n1039 = ~x4 & n1038 ;
  assign n1040 = ~x4 & x27 ;
  assign n1041 = x22 | x24 ;
  assign n1042 = x23 & ~x24 ;
  assign n1043 = x22 & n1042 ;
  assign n1044 = ( ~x22 & n1041 ) | ( ~x22 & n1043 ) | ( n1041 & n1043 ) ;
  assign n1045 = ( ~x4 & x27 ) | ( ~x4 & n1044 ) | ( x27 & n1044 ) ;
  assign n1046 = ( n1039 & ~n1040 ) | ( n1039 & n1045 ) | ( ~n1040 & n1045 ) ;
  assign n1047 = x5 | n1046 ;
  assign n1048 = x24 & x27 ;
  assign n1049 = x23 & x25 ;
  assign n1050 = ( x24 & x27 ) | ( x24 & ~n1049 ) | ( x27 & ~n1049 ) ;
  assign n1051 = ( n1042 & ~n1048 ) | ( n1042 & n1050 ) | ( ~n1048 & n1050 ) ;
  assign n1052 = x22 | x27 ;
  assign n1053 = x24 | n1052 ;
  assign n1054 = ~x22 & n1053 ;
  assign n1055 = ( n1051 & n1053 ) | ( n1051 & n1054 ) | ( n1053 & n1054 ) ;
  assign n1056 = x4 | n1055 ;
  assign n1057 = x5 & n1056 ;
  assign n1058 = n1047 & ~n1057 ;
  assign n1059 = x21 & n1058 ;
  assign n1060 = ~x20 & n1059 ;
  assign n1061 = ~x27 & n918 ;
  assign n1062 = n1060 | n1061 ;
  assign n1063 = ( n1035 & n1060 ) | ( n1035 & n1062 ) | ( n1060 & n1062 ) ;
  assign n1064 = x18 & ~n1063 ;
  assign n1065 = ~x18 & n129 ;
  assign n1066 = n1064 | n1065 ;
  assign n1067 = ( ~x19 & n84 ) | ( ~x19 & n1066 ) | ( n84 & n1066 ) ;
  assign n1068 = ~n1066 & n1067 ;
  assign n1069 = ~x14 & n1068 ;
  assign n1070 = ( x13 & ~x15 ) | ( x13 & n1069 ) | ( ~x15 & n1069 ) ;
  assign n1071 = ~x13 & n1070 ;
  assign n1072 = x12 & n1071 ;
  assign n1073 = ~x1 & n1072 ;
  assign n1074 = x3 & ~n1073 ;
  assign n1075 = n1034 & ~n1074 ;
  assign n1076 = ( x0 & ~x2 ) | ( x0 & n1075 ) | ( ~x2 & n1075 ) ;
  assign n1077 = ( x3 & x16 ) | ( x3 & ~n165 ) | ( x16 & ~n165 ) ;
  assign n1078 = ~x17 & n70 ;
  assign n1079 = ~x3 & x15 ;
  assign n1080 = n1078 & n1079 ;
  assign n1081 = x16 & n1080 ;
  assign n1082 = ( n165 & n1077 ) | ( n165 & n1081 ) | ( n1077 & n1081 ) ;
  assign n1083 = x3 | n43 ;
  assign n1084 = n94 & ~n1083 ;
  assign n1085 = ~n1082 & n1084 ;
  assign n1086 = ( n665 & n1082 ) | ( n665 & n1085 ) | ( n1082 & n1085 ) ;
  assign n1087 = ( x3 & n85 ) | ( x3 & n609 ) | ( n85 & n609 ) ;
  assign n1088 = ~x3 & n1087 ;
  assign n1089 = ~n1086 & n1088 ;
  assign n1090 = x5 | x14 ;
  assign n1091 = ( n1086 & n1089 ) | ( n1086 & ~n1090 ) | ( n1089 & ~n1090 ) ;
  assign n1092 = ~x1 & n1091 ;
  assign n1093 = ~x4 & n1092 ;
  assign n1094 = ( x0 & x2 ) | ( x0 & ~n1093 ) | ( x2 & ~n1093 ) ;
  assign n1095 = n1076 & ~n1094 ;
  assign n1096 = ( x0 & x1 ) | ( x0 & ~n1095 ) | ( x1 & ~n1095 ) ;
  assign n1097 = n930 & n1096 ;
  assign n1098 = ( n930 & n1095 ) | ( n930 & ~n1097 ) | ( n1095 & ~n1097 ) ;
  assign n1099 = ( x11 & n391 ) | ( x11 & n1098 ) | ( n391 & n1098 ) ;
  assign n1100 = n1098 & ~n1099 ;
  assign n1101 = ~x8 & n1100 ;
  assign n1102 = ~x9 & n1101 ;
  assign n1103 = ~x5 & x8 ;
  assign n1104 = ( x4 & ~x36 ) | ( x4 & n1103 ) | ( ~x36 & n1103 ) ;
  assign n1105 = ~x4 & n1104 ;
  assign n1106 = ~x2 & n1105 ;
  assign n1107 = ( x1 & ~x3 ) | ( x1 & n1106 ) | ( ~x3 & n1106 ) ;
  assign n1108 = ~x1 & n1107 ;
  assign n1109 = ~x0 & n1108 ;
  assign n1110 = x10 | n1109 ;
  assign n1111 = ( ~x8 & n1109 ) | ( ~x8 & n1110 ) | ( n1109 & n1110 ) ;
  assign n1112 = x9 & n1111 ;
  assign n1113 = ~x8 & x9 ;
  assign n1114 = ~x10 & n1113 ;
  assign n1115 = ~x13 & n304 ;
  assign n1116 = x16 & ~n95 ;
  assign n1117 = x13 & n745 ;
  assign n1118 = n1116 & n1117 ;
  assign n1119 = ~x16 & n477 ;
  assign n1120 = n1118 | n1119 ;
  assign n1121 = ( n1115 & n1118 ) | ( n1115 & n1120 ) | ( n1118 & n1120 ) ;
  assign n1122 = ( x5 & x19 ) | ( x5 & ~n1121 ) | ( x19 & ~n1121 ) ;
  assign n1123 = ~x38 & n84 ;
  assign n1124 = ( x18 & x37 ) | ( x18 & n1123 ) | ( x37 & n1123 ) ;
  assign n1125 = ~x18 & n1124 ;
  assign n1126 = x13 | n276 ;
  assign n1127 = ( x5 & n1125 ) | ( x5 & ~n1126 ) | ( n1125 & ~n1126 ) ;
  assign n1128 = ~x5 & n1127 ;
  assign n1129 = x19 & n1128 ;
  assign n1130 = ( n1121 & n1122 ) | ( n1121 & n1129 ) | ( n1122 & n1129 ) ;
  assign n1131 = x18 | n693 ;
  assign n1132 = x19 | n1131 ;
  assign n1133 = ( x16 & n136 ) | ( x16 & ~n1132 ) | ( n136 & ~n1132 ) ;
  assign n1134 = ~x16 & n1133 ;
  assign n1135 = ~x13 & n1134 ;
  assign n1136 = ( x5 & ~x14 ) | ( x5 & n1135 ) | ( ~x14 & n1135 ) ;
  assign n1137 = ~x5 & n1136 ;
  assign n1138 = ( x13 & x14 ) | ( x13 & ~x15 ) | ( x14 & ~x15 ) ;
  assign n1139 = x17 & ~n693 ;
  assign n1140 = x13 & ~x16 ;
  assign n1141 = ( n693 & n1139 ) | ( n693 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1142 = x18 & ~n1141 ;
  assign n1143 = x13 & ~n71 ;
  assign n1144 = x18 | n1143 ;
  assign n1145 = ~n1142 & n1144 ;
  assign n1146 = ( x14 & x15 ) | ( x14 & n1145 ) | ( x15 & n1145 ) ;
  assign n1147 = n1138 | n1146 ;
  assign n1148 = ~x5 & n1147 ;
  assign n1149 = ~x15 & n84 ;
  assign n1150 = x14 & n76 ;
  assign n1151 = ( x14 & n1149 ) | ( x14 & n1150 ) | ( n1149 & n1150 ) ;
  assign n1152 = ~x13 & n1151 ;
  assign n1153 = x5 & ~n1152 ;
  assign n1154 = n1148 | n1153 ;
  assign n1155 = ~x12 & n1154 ;
  assign n1156 = x14 & ~n190 ;
  assign n1157 = x17 & n1156 ;
  assign n1158 = ( x16 & ~n190 ) | ( x16 & n1156 ) | ( ~n190 & n1156 ) ;
  assign n1159 = ( ~x13 & n1157 ) | ( ~x13 & n1158 ) | ( n1157 & n1158 ) ;
  assign n1160 = x15 & ~n1159 ;
  assign n1161 = x13 & x14 ;
  assign n1162 = n71 & n1161 ;
  assign n1163 = x15 | n1162 ;
  assign n1164 = ~n1160 & n1163 ;
  assign n1165 = x16 & n416 ;
  assign n1166 = n1164 | n1165 ;
  assign n1167 = ( n1117 & n1164 ) | ( n1117 & n1166 ) | ( n1164 & n1166 ) ;
  assign n1168 = x5 & n1167 ;
  assign n1169 = x12 & ~n1168 ;
  assign n1170 = n1155 | n1169 ;
  assign n1171 = ( n1130 & ~n1137 ) | ( n1130 & n1170 ) | ( ~n1137 & n1170 ) ;
  assign n1172 = ~x12 & n1170 ;
  assign n1173 = ( ~n1130 & n1171 ) | ( ~n1130 & n1172 ) | ( n1171 & n1172 ) ;
  assign n1174 = ( ~x36 & n748 ) | ( ~x36 & n1173 ) | ( n748 & n1173 ) ;
  assign n1175 = ~n1173 & n1174 ;
  assign n1176 = ~x9 & n1175 ;
  assign n1177 = ( x4 & ~x10 ) | ( x4 & n1176 ) | ( ~x10 & n1176 ) ;
  assign n1178 = ~x4 & n1177 ;
  assign n1179 = ~x2 & n1178 ;
  assign n1180 = ( x1 & ~x3 ) | ( x1 & n1179 ) | ( ~x3 & n1179 ) ;
  assign n1181 = ~x1 & n1180 ;
  assign n1182 = ( x0 & ~x8 ) | ( x0 & n1181 ) | ( ~x8 & n1181 ) ;
  assign n1183 = x10 & n726 ;
  assign n1184 = ~x8 & n1183 ;
  assign n1185 = ( ~x0 & n1182 ) | ( ~x0 & n1184 ) | ( n1182 & n1184 ) ;
  assign n1186 = n1114 | n1185 ;
  assign n1187 = ( n1111 & ~n1112 ) | ( n1111 & n1186 ) | ( ~n1112 & n1186 ) ;
  assign n1188 = ( x8 & ~x9 ) | ( x8 & x10 ) | ( ~x9 & x10 ) ;
  assign n1189 = x10 & ~n1188 ;
  assign n1190 = ( n165 & n503 ) | ( n165 & n504 ) | ( n503 & n504 ) ;
  assign n1191 = ( x14 & ~n665 ) | ( x14 & n1190 ) | ( ~n665 & n1190 ) ;
  assign n1192 = n1190 & ~n1191 ;
  assign n1193 = ~x2 & n1192 ;
  assign n1194 = ( x1 & ~x3 ) | ( x1 & n1193 ) | ( ~x3 & n1193 ) ;
  assign n1195 = ~x1 & n1194 ;
  assign n1196 = x0 & n1195 ;
  assign n1197 = ( x13 & x17 ) | ( x13 & n239 ) | ( x17 & n239 ) ;
  assign n1198 = ~x13 & n1197 ;
  assign n1199 = x4 & ~x14 ;
  assign n1200 = ( ~x14 & n601 ) | ( ~x14 & n1199 ) | ( n601 & n1199 ) ;
  assign n1201 = x13 & ~n1200 ;
  assign n1202 = ~n129 & n239 ;
  assign n1203 = x13 | n1202 ;
  assign n1204 = ~n1201 & n1203 ;
  assign n1205 = ( x17 & x18 ) | ( x17 & n1204 ) | ( x18 & n1204 ) ;
  assign n1206 = ~x5 & n245 ;
  assign n1207 = ( x4 & ~x13 ) | ( x4 & n1206 ) | ( ~x13 & n1206 ) ;
  assign n1208 = ~x4 & n1207 ;
  assign n1209 = ~x17 & n1208 ;
  assign n1210 = ( n1204 & ~n1205 ) | ( n1204 & n1209 ) | ( ~n1205 & n1209 ) ;
  assign n1211 = ( x4 & x5 ) | ( x4 & ~n1210 ) | ( x5 & ~n1210 ) ;
  assign n1212 = n1198 & n1211 ;
  assign n1213 = ( n1198 & n1210 ) | ( n1198 & ~n1212 ) | ( n1210 & ~n1212 ) ;
  assign n1214 = x15 & n1213 ;
  assign n1215 = ( x17 & ~n95 ) | ( x17 & n931 ) | ( ~n95 & n931 ) ;
  assign n1216 = ( x5 & n190 ) | ( x5 & n1215 ) | ( n190 & n1215 ) ;
  assign n1217 = ~x5 & n1216 ;
  assign n1218 = n1214 | n1217 ;
  assign n1219 = ( ~x4 & n1214 ) | ( ~x4 & n1218 ) | ( n1214 & n1218 ) ;
  assign n1220 = ~x12 & n1219 ;
  assign n1221 = x15 & x40 ;
  assign n1222 = ( ~x14 & x17 ) | ( ~x14 & n1221 ) | ( x17 & n1221 ) ;
  assign n1223 = x14 & n1222 ;
  assign n1224 = x13 & n1223 ;
  assign n1225 = ( x5 & x12 ) | ( x5 & n1224 ) | ( x12 & n1224 ) ;
  assign n1226 = ~x5 & n1225 ;
  assign n1227 = n1220 | n1226 ;
  assign n1228 = ( ~x4 & n1220 ) | ( ~x4 & n1227 ) | ( n1220 & n1227 ) ;
  assign n1229 = ~x14 & n109 ;
  assign n1230 = ( x12 & x13 ) | ( x12 & n1229 ) | ( x13 & n1229 ) ;
  assign n1231 = ~x12 & n1230 ;
  assign n1232 = ( x3 & n118 ) | ( x3 & ~n1231 ) | ( n118 & ~n1231 ) ;
  assign n1233 = ( x3 & n118 ) | ( x3 & ~n1228 ) | ( n118 & ~n1228 ) ;
  assign n1234 = ( n1228 & ~n1232 ) | ( n1228 & n1233 ) | ( ~n1232 & n1233 ) ;
  assign n1235 = x1 & n1234 ;
  assign n1236 = x1 & ~x2 ;
  assign n1237 = ~x14 & n665 ;
  assign n1238 = ~n275 & n1237 ;
  assign n1239 = ( ~n109 & n1236 ) | ( ~n109 & n1238 ) | ( n1236 & n1238 ) ;
  assign n1240 = n109 & n1239 ;
  assign n1241 = ~x16 & n418 ;
  assign n1242 = n304 & n1241 ;
  assign n1243 = x13 | x17 ;
  assign n1244 = ( n95 & n558 ) | ( n95 & ~n1243 ) | ( n558 & ~n1243 ) ;
  assign n1245 = ( ~x12 & n558 ) | ( ~x12 & n1244 ) | ( n558 & n1244 ) ;
  assign n1246 = ( x16 & n931 ) | ( x16 & ~n1245 ) | ( n931 & ~n1245 ) ;
  assign n1247 = n1245 & n1246 ;
  assign n1248 = ( x4 & n1029 ) | ( x4 & n1247 ) | ( n1029 & n1247 ) ;
  assign n1249 = ~x4 & n1248 ;
  assign n1250 = ( x13 & x16 ) | ( x13 & n58 ) | ( x16 & n58 ) ;
  assign n1251 = ~x13 & n1250 ;
  assign n1252 = x37 & ~x38 ;
  assign n1253 = ~x39 & n1252 ;
  assign n1254 = ( x18 & n396 ) | ( x18 & n1253 ) | ( n396 & n1253 ) ;
  assign n1255 = ~n1253 & n1254 ;
  assign n1256 = x4 & ~n601 ;
  assign n1257 = ( n418 & n601 ) | ( n418 & n1256 ) | ( n601 & n1256 ) ;
  assign n1258 = ( x4 & x5 ) | ( x4 & ~n1257 ) | ( x5 & ~n1257 ) ;
  assign n1259 = n1255 & n1258 ;
  assign n1260 = ( n1255 & n1257 ) | ( n1255 & ~n1259 ) | ( n1257 & ~n1259 ) ;
  assign n1261 = ( x16 & ~n665 ) | ( x16 & n1260 ) | ( ~n665 & n1260 ) ;
  assign n1262 = n1260 & ~n1261 ;
  assign n1263 = ( x4 & x5 ) | ( x4 & ~n1262 ) | ( x5 & ~n1262 ) ;
  assign n1264 = n1251 & n1263 ;
  assign n1265 = ( n1251 & n1262 ) | ( n1251 & ~n1264 ) | ( n1262 & ~n1264 ) ;
  assign n1266 = ( ~x14 & n1249 ) | ( ~x14 & n1265 ) | ( n1249 & n1265 ) ;
  assign n1267 = x15 & ~n1266 ;
  assign n1268 = ( x15 & n1249 ) | ( x15 & ~n1267 ) | ( n1249 & ~n1267 ) ;
  assign n1269 = ~x3 & n1268 ;
  assign n1270 = x3 & ~x5 ;
  assign n1271 = ( x4 & n665 ) | ( x4 & n1270 ) | ( n665 & n1270 ) ;
  assign n1272 = ~x4 & n1271 ;
  assign n1273 = n1269 | n1272 ;
  assign n1274 = ( n1242 & n1269 ) | ( n1242 & n1273 ) | ( n1269 & n1273 ) ;
  assign n1275 = ( x1 & x2 ) | ( x1 & n1274 ) | ( x2 & n1274 ) ;
  assign n1276 = x5 & ~x12 ;
  assign n1277 = x1 & ~x4 ;
  assign n1278 = ( x3 & n1276 ) | ( x3 & n1277 ) | ( n1276 & n1277 ) ;
  assign n1279 = ~x3 & n1278 ;
  assign n1280 = x13 & n1279 ;
  assign n1281 = ( n304 & ~n1116 ) | ( n304 & n1280 ) | ( ~n1116 & n1280 ) ;
  assign n1282 = n1116 & n1281 ;
  assign n1283 = ~x2 & n1282 ;
  assign n1284 = ( n1274 & ~n1275 ) | ( n1274 & n1283 ) | ( ~n1275 & n1283 ) ;
  assign n1285 = n1240 | n1284 ;
  assign n1286 = ( n1234 & ~n1235 ) | ( n1234 & n1285 ) | ( ~n1235 & n1285 ) ;
  assign n1287 = ~x21 & x27 ;
  assign n1288 = ( x19 & x20 ) | ( x19 & n1287 ) | ( x20 & n1287 ) ;
  assign n1289 = ~x19 & n1288 ;
  assign n1290 = n1119 & n1289 ;
  assign n1291 = n155 | n608 ;
  assign n1292 = ( x1 & n515 ) | ( x1 & ~n1291 ) | ( n515 & ~n1291 ) ;
  assign n1293 = ~x1 & n1292 ;
  assign n1294 = ( x2 & ~n1290 ) | ( x2 & n1293 ) | ( ~n1290 & n1293 ) ;
  assign n1295 = n96 & n110 ;
  assign n1296 = x1 | n1295 ;
  assign n1297 = ( n138 & n1295 ) | ( n138 & n1296 ) | ( n1295 & n1296 ) ;
  assign n1298 = x13 & n1297 ;
  assign n1299 = ~x12 & n1298 ;
  assign n1300 = x2 & n1299 ;
  assign n1301 = ( n1290 & n1294 ) | ( n1290 & n1300 ) | ( n1294 & n1300 ) ;
  assign n1302 = n66 & n110 ;
  assign n1303 = ( ~x3 & x17 ) | ( ~x3 & n1302 ) | ( x17 & n1302 ) ;
  assign n1304 = x15 & ~x19 ;
  assign n1305 = ( n110 & ~n133 ) | ( n110 & n1304 ) | ( ~n133 & n1304 ) ;
  assign n1306 = x18 & n1305 ;
  assign n1307 = x4 & n1306 ;
  assign n1308 = x18 & n601 ;
  assign n1309 = n1305 & n1308 ;
  assign n1310 = ~x19 & x40 ;
  assign n1311 = ~x18 & n1310 ;
  assign n1312 = ~x5 & n1311 ;
  assign n1313 = n110 & n1312 ;
  assign n1314 = n1309 | n1313 ;
  assign n1315 = ~x4 & n1314 ;
  assign n1316 = n1307 | n1315 ;
  assign n1317 = ( x3 & x17 ) | ( x3 & n1316 ) | ( x17 & n1316 ) ;
  assign n1318 = n1303 & n1317 ;
  assign n1319 = n559 & n1318 ;
  assign n1320 = ( x20 & x22 ) | ( x20 & x23 ) | ( x22 & x23 ) ;
  assign n1321 = x24 & ~n1320 ;
  assign n1322 = ( x20 & x24 ) | ( x20 & ~n1321 ) | ( x24 & ~n1321 ) ;
  assign n1323 = x20 | x21 ;
  assign n1324 = x22 & x24 ;
  assign n1325 = x23 & n1324 ;
  assign n1326 = x20 | n1325 ;
  assign n1327 = x21 & ~n1326 ;
  assign n1328 = ( ~x21 & n1323 ) | ( ~x21 & n1327 ) | ( n1323 & n1327 ) ;
  assign n1329 = x21 | n1328 ;
  assign n1330 = ( n1322 & n1328 ) | ( n1322 & n1329 ) | ( n1328 & n1329 ) ;
  assign n1331 = ( x17 & n369 ) | ( x17 & ~n1330 ) | ( n369 & ~n1330 ) ;
  assign n1332 = n1330 & n1331 ;
  assign n1333 = ( x15 & x40 ) | ( x15 & n1332 ) | ( x40 & n1332 ) ;
  assign n1334 = ( n110 & ~n126 ) | ( n110 & n136 ) | ( ~n126 & n136 ) ;
  assign n1335 = ( x18 & n693 ) | ( x18 & ~n1334 ) | ( n693 & ~n1334 ) ;
  assign n1336 = ( x15 & ~x16 ) | ( x15 & x17 ) | ( ~x16 & x17 ) ;
  assign n1337 = ~x15 & n1336 ;
  assign n1338 = ( x17 & n694 ) | ( x17 & ~n1337 ) | ( n694 & ~n1337 ) ;
  assign n1339 = ( n1336 & n1337 ) | ( n1336 & ~n1338 ) | ( n1337 & ~n1338 ) ;
  assign n1340 = ~x18 & n1339 ;
  assign n1341 = ( n693 & ~n1335 ) | ( n693 & n1340 ) | ( ~n1335 & n1340 ) ;
  assign n1342 = x40 & n1341 ;
  assign n1343 = ( ~x15 & n1333 ) | ( ~x15 & n1342 ) | ( n1333 & n1342 ) ;
  assign n1344 = ( ~x21 & x23 ) | ( ~x21 & n1324 ) | ( x23 & n1324 ) ;
  assign n1345 = x21 & n1344 ;
  assign n1346 = x20 & n1345 ;
  assign n1347 = x18 & ~n1328 ;
  assign n1348 = ( ~n1345 & n1346 ) | ( ~n1345 & n1347 ) | ( n1346 & n1347 ) ;
  assign n1349 = ( ~x16 & n570 ) | ( ~x16 & n1348 ) | ( n570 & n1348 ) ;
  assign n1350 = ~n1348 & n1349 ;
  assign n1351 = ( x5 & n114 ) | ( x5 & ~n1350 ) | ( n114 & ~n1350 ) ;
  assign n1352 = ( x5 & n114 ) | ( x5 & ~n1343 ) | ( n114 & ~n1343 ) ;
  assign n1353 = ( n1343 & ~n1351 ) | ( n1343 & n1352 ) | ( ~n1351 & n1352 ) ;
  assign n1354 = x3 | n1353 ;
  assign n1355 = x5 & ~x27 ;
  assign n1356 = ( x4 & ~x27 ) | ( x4 & n1355 ) | ( ~x27 & n1355 ) ;
  assign n1357 = x20 & ~n972 ;
  assign n1358 = ~n1356 & n1357 ;
  assign n1359 = x27 & ~n561 ;
  assign n1360 = ~x24 & n1359 ;
  assign n1361 = x4 & n1360 ;
  assign n1362 = ( x24 & n561 ) | ( x24 & ~n1359 ) | ( n561 & ~n1359 ) ;
  assign n1363 = ( x23 & ~x24 ) | ( x23 & x25 ) | ( ~x24 & x25 ) ;
  assign n1364 = x23 & x27 ;
  assign n1365 = ( x24 & n1363 ) | ( x24 & n1364 ) | ( n1363 & n1364 ) ;
  assign n1366 = x22 & n1365 ;
  assign n1367 = ~x5 & n1366 ;
  assign n1368 = ( x5 & n1362 ) | ( x5 & ~n1367 ) | ( n1362 & ~n1367 ) ;
  assign n1369 = x22 & ~x24 ;
  assign n1370 = x5 & x27 ;
  assign n1371 = ( ~x22 & n1369 ) | ( ~x22 & n1370 ) | ( n1369 & n1370 ) ;
  assign n1372 = n1368 & ~n1371 ;
  assign n1373 = x4 | n1372 ;
  assign n1374 = ~n1361 & n1373 ;
  assign n1375 = ( n972 & ~n1357 ) | ( n972 & n1374 ) | ( ~n1357 & n1374 ) ;
  assign n1376 = ( x21 & n1358 ) | ( x21 & ~n1375 ) | ( n1358 & ~n1375 ) ;
  assign n1377 = ( x17 & n369 ) | ( x17 & ~n1376 ) | ( n369 & ~n1376 ) ;
  assign n1378 = n1376 & n1377 ;
  assign n1379 = ~x15 & n1378 ;
  assign n1380 = x3 & ~n1379 ;
  assign n1381 = n1354 & ~n1380 ;
  assign n1382 = ~x19 & n1381 ;
  assign n1383 = x15 & x18 ;
  assign n1384 = x17 & ~x39 ;
  assign n1385 = ( x17 & x18 ) | ( x17 & ~n1384 ) | ( x18 & ~n1384 ) ;
  assign n1386 = ( x15 & x18 ) | ( x15 & n1385 ) | ( x18 & n1385 ) ;
  assign n1387 = ( n1383 & n1385 ) | ( n1383 & ~n1386 ) | ( n1385 & ~n1386 ) ;
  assign n1388 = x40 & n1387 ;
  assign n1389 = x5 | n1388 ;
  assign n1390 = x15 & n416 ;
  assign n1391 = x5 & ~n1390 ;
  assign n1392 = n1389 & ~n1391 ;
  assign n1393 = ~x4 & n1392 ;
  assign n1394 = x4 & x15 ;
  assign n1395 = ( x5 & n416 ) | ( x5 & n1394 ) | ( n416 & n1394 ) ;
  assign n1396 = ~x5 & n1395 ;
  assign n1397 = ~n1393 & n1396 ;
  assign n1398 = ( n296 & n1393 ) | ( n296 & n1397 ) | ( n1393 & n1397 ) ;
  assign n1399 = n1382 | n1398 ;
  assign n1400 = ( ~x3 & n1382 ) | ( ~x3 & n1399 ) | ( n1382 & n1399 ) ;
  assign n1401 = ( ~n558 & n559 ) | ( ~n558 & n1400 ) | ( n559 & n1400 ) ;
  assign n1402 = ( x12 & n1319 ) | ( x12 & n1401 ) | ( n1319 & n1401 ) ;
  assign n1403 = ( x1 & ~x2 ) | ( x1 & n1402 ) | ( ~x2 & n1402 ) ;
  assign n1404 = x3 | n1295 ;
  assign n1405 = ( n138 & n1295 ) | ( n138 & n1404 ) | ( n1295 & n1404 ) ;
  assign n1406 = ( ~x3 & n138 ) | ( ~x3 & n1405 ) | ( n138 & n1405 ) ;
  assign n1407 = x4 & ~n1406 ;
  assign n1408 = ( x4 & n1405 ) | ( x4 & ~n1407 ) | ( n1405 & ~n1407 ) ;
  assign n1409 = x15 & ~n155 ;
  assign n1410 = ( x5 & ~n160 ) | ( x5 & n1409 ) | ( ~n160 & n1409 ) ;
  assign n1411 = n160 & n1410 ;
  assign n1412 = ~n1408 & n1411 ;
  assign n1413 = ( n665 & n1408 ) | ( n665 & n1412 ) | ( n1408 & n1412 ) ;
  assign n1414 = ( x1 & x2 ) | ( x1 & ~n1413 ) | ( x2 & ~n1413 ) ;
  assign n1415 = n1403 & ~n1414 ;
  assign n1416 = x19 & x40 ;
  assign n1417 = ~x18 & n1416 ;
  assign n1418 = n126 & n558 ;
  assign n1419 = ( n745 & ~n1417 ) | ( n745 & n1418 ) | ( ~n1417 & n1418 ) ;
  assign n1420 = n1417 & n1419 ;
  assign n1421 = x40 | n1420 ;
  assign n1422 = ( n129 & ~n1420 ) | ( n129 & n1421 ) | ( ~n1420 & n1421 ) ;
  assign n1423 = x2 | n1422 ;
  assign n1424 = ( ~x1 & x3 ) | ( ~x1 & n1423 ) | ( x3 & n1423 ) ;
  assign n1425 = x1 | n1424 ;
  assign n1426 = ( n1301 & ~n1415 ) | ( n1301 & n1425 ) | ( ~n1415 & n1425 ) ;
  assign n1427 = x14 & n1425 ;
  assign n1428 = ( ~n1301 & n1426 ) | ( ~n1301 & n1427 ) | ( n1426 & n1427 ) ;
  assign n1429 = ~n1286 & n1428 ;
  assign n1430 = x0 | n1429 ;
  assign n1431 = ~n1196 & n1430 ;
  assign n1432 = ~x11 & x36 ;
  assign n1433 = ( x11 & n1431 ) | ( x11 & ~n1432 ) | ( n1431 & ~n1432 ) ;
  assign n1434 = ( x9 & ~n1189 ) | ( x9 & n1433 ) | ( ~n1189 & n1433 ) ;
  assign n1435 = ( n1188 & ~n1189 ) | ( n1188 & n1434 ) | ( ~n1189 & n1434 ) ;
  assign n1436 = x12 & ~x15 ;
  assign n1437 = x13 & n1436 ;
  assign n1438 = x15 & x19 ;
  assign n1439 = ( ~x13 & x16 ) | ( ~x13 & n1438 ) | ( x16 & n1438 ) ;
  assign n1440 = x13 & n1439 ;
  assign n1441 = x13 | x18 ;
  assign n1442 = x12 & x18 ;
  assign n1443 = x13 & x19 ;
  assign n1444 = x12 & ~n1443 ;
  assign n1445 = ( n1441 & ~n1442 ) | ( n1441 & n1444 ) | ( ~n1442 & n1444 ) ;
  assign n1446 = x16 | n1445 ;
  assign n1447 = x15 | n1446 ;
  assign n1448 = ~x12 & n1447 ;
  assign n1449 = ( ~n1440 & n1447 ) | ( ~n1440 & n1448 ) | ( n1447 & n1448 ) ;
  assign n1450 = x17 | n1449 ;
  assign n1451 = ~n85 & n1450 ;
  assign n1452 = ( ~n1437 & n1450 ) | ( ~n1437 & n1451 ) | ( n1450 & n1451 ) ;
  assign n1453 = x14 & n1452 ;
  assign n1454 = ( ~x13 & x15 ) | ( ~x13 & x16 ) | ( x15 & x16 ) ;
  assign n1455 = x13 & n1454 ;
  assign n1456 = ( ~x15 & n1078 ) | ( ~x15 & n1455 ) | ( n1078 & n1455 ) ;
  assign n1457 = ( n1454 & n1455 ) | ( n1454 & n1456 ) | ( n1455 & n1456 ) ;
  assign n1458 = x12 & n1457 ;
  assign n1459 = x14 | n1458 ;
  assign n1460 = ~n1453 & n1459 ;
  assign n1461 = ( x36 & ~n748 ) | ( x36 & n1460 ) | ( ~n748 & n1460 ) ;
  assign n1462 = n1460 & ~n1461 ;
  assign n1463 = ~x9 & n1462 ;
  assign n1464 = ( x8 & ~x10 ) | ( x8 & n1463 ) | ( ~x10 & n1463 ) ;
  assign n1465 = ~x8 & n1464 ;
  assign n1466 = ~x4 & n1465 ;
  assign n1467 = ( x3 & ~x5 ) | ( x3 & n1466 ) | ( ~x5 & n1466 ) ;
  assign n1468 = ~x3 & n1467 ;
  assign n1469 = ~x1 & n1468 ;
  assign n1470 = ( x0 & ~x2 ) | ( x0 & n1469 ) | ( ~x2 & n1469 ) ;
  assign n1471 = ~x0 & n1470 ;
  assign n1472 = ( ~x18 & n84 ) | ( ~x18 & n878 ) | ( n84 & n878 ) ;
  assign n1473 = n304 & n1472 ;
  assign n1474 = ( x11 & n665 ) | ( x11 & n1473 ) | ( n665 & n1473 ) ;
  assign n1475 = ~x11 & n1474 ;
  assign n1476 = ~x8 & n1475 ;
  assign n1477 = ~x10 & n1476 ;
  assign n1478 = x3 & n1477 ;
  assign n1479 = ~x38 & n70 ;
  assign n1480 = x37 & n1479 ;
  assign n1481 = x17 & ~x19 ;
  assign n1482 = ( n416 & ~n878 ) | ( n416 & n1481 ) | ( ~n878 & n1481 ) ;
  assign n1483 = x13 & ~n665 ;
  assign n1484 = n1482 & n1483 ;
  assign n1485 = ( n95 & n665 ) | ( n95 & ~n1483 ) | ( n665 & ~n1483 ) ;
  assign n1486 = ( x12 & ~n1484 ) | ( x12 & n1485 ) | ( ~n1484 & n1485 ) ;
  assign n1487 = x14 & ~n1486 ;
  assign n1488 = n153 & n530 ;
  assign n1489 = n1487 | n1488 ;
  assign n1490 = ( n1480 & n1487 ) | ( n1480 & n1489 ) | ( n1487 & n1489 ) ;
  assign n1491 = ( x15 & ~x40 ) | ( x15 & n1490 ) | ( ~x40 & n1490 ) ;
  assign n1492 = x13 & x18 ;
  assign n1493 = x12 & ~x18 ;
  assign n1494 = x13 | x19 ;
  assign n1495 = x12 & n1494 ;
  assign n1496 = ( n1492 & n1493 ) | ( n1492 & ~n1495 ) | ( n1493 & ~n1495 ) ;
  assign n1497 = ( x39 & ~n1252 ) | ( x39 & n1496 ) | ( ~n1252 & n1496 ) ;
  assign n1498 = n1496 & ~n1497 ;
  assign n1499 = ~x17 & n1498 ;
  assign n1500 = ( x14 & x15 ) | ( x14 & n1499 ) | ( x15 & n1499 ) ;
  assign n1501 = ~x14 & n1500 ;
  assign n1502 = x40 & n1501 ;
  assign n1503 = ( n1490 & ~n1491 ) | ( n1490 & n1502 ) | ( ~n1491 & n1502 ) ;
  assign n1504 = ~x11 & n1503 ;
  assign n1505 = ( x10 & ~x16 ) | ( x10 & n1504 ) | ( ~x16 & n1504 ) ;
  assign n1506 = ~x10 & n1505 ;
  assign n1507 = x8 | n1506 ;
  assign n1508 = ~x3 & n1507 ;
  assign n1509 = n1478 | n1508 ;
  assign n1510 = x4 | x36 ;
  assign n1511 = ( x5 & n1509 ) | ( x5 & n1510 ) | ( n1509 & n1510 ) ;
  assign n1512 = n1509 & ~n1511 ;
  assign n1513 = ~x1 & n1512 ;
  assign n1514 = ( x0 & ~x2 ) | ( x0 & n1513 ) | ( ~x2 & n1513 ) ;
  assign n1515 = ~x0 & n1514 ;
  assign n1516 = x10 | n1515 ;
  assign n1517 = ( ~x8 & n1515 ) | ( ~x8 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = ~x9 & n1517 ;
  assign n1519 = n727 | n1518 ;
  assign n1520 = ( ~x8 & n1518 ) | ( ~x8 & n1519 ) | ( n1518 & n1519 ) ;
  assign n1521 = ~x12 & x14 ;
  assign n1522 = ( x14 & x15 ) | ( x14 & ~x16 ) | ( x15 & ~x16 ) ;
  assign n1523 = ( ~x12 & x15 ) | ( ~x12 & n1522 ) | ( x15 & n1522 ) ;
  assign n1524 = ( x15 & n1521 ) | ( x15 & ~n1523 ) | ( n1521 & ~n1523 ) ;
  assign n1525 = n1521 | n1524 ;
  assign n1526 = ( n1149 & n1524 ) | ( n1149 & n1525 ) | ( n1524 & n1525 ) ;
  assign n1527 = x13 | n1526 ;
  assign n1528 = x17 & n76 ;
  assign n1529 = x14 & n1528 ;
  assign n1530 = x12 & n1529 ;
  assign n1531 = x13 & ~n1530 ;
  assign n1532 = n1527 & ~n1531 ;
  assign n1533 = n110 & n416 ;
  assign n1534 = ( n1161 & n1532 ) | ( n1161 & n1533 ) | ( n1532 & n1533 ) ;
  assign n1535 = x12 & ~n1534 ;
  assign n1536 = ( x12 & n1532 ) | ( x12 & ~n1535 ) | ( n1532 & ~n1535 ) ;
  assign n1537 = ( x12 & n1121 ) | ( x12 & n1536 ) | ( n1121 & n1536 ) ;
  assign n1538 = x19 & ~n1537 ;
  assign n1539 = ( x19 & n1536 ) | ( x19 & ~n1538 ) | ( n1536 & ~n1538 ) ;
  assign n1540 = ~x10 & x40 ;
  assign n1541 = ( x11 & n1539 ) | ( x11 & ~n1540 ) | ( n1539 & ~n1540 ) ;
  assign n1542 = n1539 & ~n1541 ;
  assign n1543 = ( x5 & x8 ) | ( x5 & ~n1542 ) | ( x8 & ~n1542 ) ;
  assign n1544 = x5 & n1543 ;
  assign n1545 = x14 | n635 ;
  assign n1546 = ( ~x15 & x16 ) | ( ~x15 & x18 ) | ( x16 & x18 ) ;
  assign n1547 = ( x15 & ~x16 ) | ( x15 & x19 ) | ( ~x16 & x19 ) ;
  assign n1548 = n1546 & n1547 ;
  assign n1549 = ~x17 & n1548 ;
  assign n1550 = x14 & ~n1549 ;
  assign n1551 = n1545 & ~n1550 ;
  assign n1552 = x19 | n76 ;
  assign n1553 = x17 & ~n1552 ;
  assign n1554 = n635 | n1553 ;
  assign n1555 = ( n51 & n1553 ) | ( n51 & n1554 ) | ( n1553 & n1554 ) ;
  assign n1556 = n1156 & n1555 ;
  assign n1557 = x37 & n570 ;
  assign n1558 = x19 & n1557 ;
  assign n1559 = ( x17 & ~x39 ) | ( x17 & n1304 ) | ( ~x39 & n1304 ) ;
  assign n1560 = ~x17 & n1559 ;
  assign n1561 = ~x38 & n1560 ;
  assign n1562 = ( ~x38 & n1558 ) | ( ~x38 & n1561 ) | ( n1558 & n1561 ) ;
  assign n1563 = x16 | n1562 ;
  assign n1564 = ~x15 & n51 ;
  assign n1565 = x16 & ~n1564 ;
  assign n1566 = n1563 & ~n1565 ;
  assign n1567 = ( ~n190 & n1156 ) | ( ~n190 & n1566 ) | ( n1156 & n1566 ) ;
  assign n1568 = ( ~x13 & n1556 ) | ( ~x13 & n1567 ) | ( n1556 & n1567 ) ;
  assign n1569 = ~x18 & n1568 ;
  assign n1570 = x13 | n1569 ;
  assign n1571 = ( n1551 & n1569 ) | ( n1551 & n1570 ) | ( n1569 & n1570 ) ;
  assign n1572 = x12 & n1571 ;
  assign n1573 = x16 | n95 ;
  assign n1574 = x13 | n1573 ;
  assign n1575 = n745 & ~n1574 ;
  assign n1576 = n1147 & ~n1575 ;
  assign n1577 = x12 | n1576 ;
  assign n1578 = ~n1572 & n1577 ;
  assign n1579 = ( ~x11 & n1540 ) | ( ~x11 & n1578 ) | ( n1540 & n1578 ) ;
  assign n1580 = ~n1578 & n1579 ;
  assign n1581 = x5 | x8 ;
  assign n1582 = ( ~n1544 & n1580 ) | ( ~n1544 & n1581 ) | ( n1580 & n1581 ) ;
  assign n1583 = ~n1544 & n1582 ;
  assign n1584 = x3 | n1583 ;
  assign n1585 = ~x5 & n1477 ;
  assign n1586 = x3 & ~n1585 ;
  assign n1587 = n1584 & ~n1586 ;
  assign n1588 = x2 | x36 ;
  assign n1589 = ( x4 & n1587 ) | ( x4 & n1588 ) | ( n1587 & n1588 ) ;
  assign n1590 = n1587 & ~n1589 ;
  assign n1591 = ~x8 & x11 ;
  assign n1592 = x10 & n1591 ;
  assign n1593 = ( x0 & x1 ) | ( x0 & ~n1592 ) | ( x1 & ~n1592 ) ;
  assign n1594 = n1590 & n1593 ;
  assign n1595 = ( n1590 & n1592 ) | ( n1590 & ~n1594 ) | ( n1592 & ~n1594 ) ;
  assign n1596 = ~x9 & n1595 ;
  assign n1597 = n727 | n1596 ;
  assign n1598 = ( ~x8 & n1596 ) | ( ~x8 & n1597 ) | ( n1596 & n1597 ) ;
  assign n1599 = ( x3 & ~x14 ) | ( x3 & n661 ) | ( ~x14 & n661 ) ;
  assign n1600 = n109 & n665 ;
  assign n1601 = x5 & ~n1041 ;
  assign n1602 = x5 | n1044 ;
  assign n1603 = ( ~x5 & n1601 ) | ( ~x5 & n1602 ) | ( n1601 & n1602 ) ;
  assign n1604 = ( x21 & n592 ) | ( x21 & ~n1603 ) | ( n592 & ~n1603 ) ;
  assign n1605 = n1603 & n1604 ;
  assign n1606 = x17 & n1605 ;
  assign n1607 = ( x18 & x19 ) | ( x18 & n1606 ) | ( x19 & n1606 ) ;
  assign n1608 = ~x19 & n1607 ;
  assign n1609 = ( x13 & n1436 ) | ( x13 & n1608 ) | ( n1436 & n1608 ) ;
  assign n1610 = ~x13 & n1609 ;
  assign n1611 = ( n578 & ~n1600 ) | ( n578 & n1610 ) | ( ~n1600 & n1610 ) ;
  assign n1612 = ( ~n579 & n1600 ) | ( ~n579 & n1611 ) | ( n1600 & n1611 ) ;
  assign n1613 = ( x3 & x14 ) | ( x3 & ~n1612 ) | ( x14 & ~n1612 ) ;
  assign n1614 = n1599 & ~n1613 ;
  assign n1615 = x4 & n1614 ;
  assign n1616 = ( x16 & x17 ) | ( x16 & ~n952 ) | ( x17 & ~n952 ) ;
  assign n1617 = ( ~x15 & x16 ) | ( ~x15 & n952 ) | ( x16 & n952 ) ;
  assign n1618 = n1616 & ~n1617 ;
  assign n1619 = ( x15 & x19 ) | ( x15 & ~n322 ) | ( x19 & ~n322 ) ;
  assign n1620 = ( x16 & ~x18 ) | ( x16 & n1619 ) | ( ~x18 & n1619 ) ;
  assign n1621 = ~x19 & n1620 ;
  assign n1622 = ( x15 & n322 ) | ( x15 & ~n1621 ) | ( n322 & ~n1621 ) ;
  assign n1623 = ( x18 & n1620 ) | ( x18 & ~n1622 ) | ( n1620 & ~n1622 ) ;
  assign n1624 = ~x17 & n1623 ;
  assign n1625 = ( ~x15 & x18 ) | ( ~x15 & n736 ) | ( x18 & n736 ) ;
  assign n1626 = ( x15 & ~x19 ) | ( x15 & n1625 ) | ( ~x19 & n1625 ) ;
  assign n1627 = ( ~x15 & x19 ) | ( ~x15 & n1626 ) | ( x19 & n1626 ) ;
  assign n1628 = ( ~x18 & n1626 ) | ( ~x18 & n1627 ) | ( n1626 & n1627 ) ;
  assign n1629 = x16 & ~n1628 ;
  assign n1630 = x17 & ~n1629 ;
  assign n1631 = n1624 | n1630 ;
  assign n1632 = ~n1618 & n1631 ;
  assign n1633 = x14 | n1632 ;
  assign n1634 = ~n745 & n1633 ;
  assign n1635 = x13 | n1634 ;
  assign n1636 = x17 & n1573 ;
  assign n1637 = x14 & x15 ;
  assign n1638 = ( ~n1573 & n1636 ) | ( ~n1573 & n1637 ) | ( n1636 & n1637 ) ;
  assign n1639 = ~x29 & x31 ;
  assign n1640 = x29 & ~n972 ;
  assign n1641 = n1639 | n1640 ;
  assign n1642 = ( ~x14 & x15 ) | ( ~x14 & n1641 ) | ( x15 & n1641 ) ;
  assign n1643 = ( ~x16 & x18 ) | ( ~x16 & x19 ) | ( x18 & x19 ) ;
  assign n1644 = x17 & ~n1643 ;
  assign n1645 = ( x16 & ~x17 ) | ( x16 & n1643 ) | ( ~x17 & n1643 ) ;
  assign n1646 = ( ~x16 & n1644 ) | ( ~x16 & n1645 ) | ( n1644 & n1645 ) ;
  assign n1647 = ( x14 & x15 ) | ( x14 & n1646 ) | ( x15 & n1646 ) ;
  assign n1648 = n1642 | n1647 ;
  assign n1649 = ~n1638 & n1648 ;
  assign n1650 = x13 & ~n1649 ;
  assign n1651 = n1635 & ~n1650 ;
  assign n1652 = ( x12 & ~x40 ) | ( x12 & n1651 ) | ( ~x40 & n1651 ) ;
  assign n1653 = ( n76 & n190 ) | ( n76 & n192 ) | ( n190 & n192 ) ;
  assign n1654 = ( ~x14 & n190 ) | ( ~x14 & n1653 ) | ( n190 & n1653 ) ;
  assign n1655 = n952 | n1654 ;
  assign n1656 = ( ~x18 & x19 ) | ( ~x18 & n76 ) | ( x19 & n76 ) ;
  assign n1657 = ( ~x18 & n76 ) | ( ~x18 & n878 ) | ( n76 & n878 ) ;
  assign n1658 = ( x19 & ~n1656 ) | ( x19 & n1657 ) | ( ~n1656 & n1657 ) ;
  assign n1659 = x14 & n1658 ;
  assign n1660 = ~x13 & n1659 ;
  assign n1661 = ~x15 & x19 ;
  assign n1662 = x17 & n1661 ;
  assign n1663 = ~n136 & n1662 ;
  assign n1664 = ( n136 & n797 ) | ( n136 & n1663 ) | ( n797 & n1663 ) ;
  assign n1665 = ( x13 & x15 ) | ( x13 & x17 ) | ( x15 & x17 ) ;
  assign n1666 = ( ~x14 & x17 ) | ( ~x14 & n1665 ) | ( x17 & n1665 ) ;
  assign n1667 = x17 & ~n1666 ;
  assign n1668 = n1666 | n1667 ;
  assign n1669 = ( ~x17 & n1667 ) | ( ~x17 & n1668 ) | ( n1667 & n1668 ) ;
  assign n1670 = ( x16 & x18 ) | ( x16 & n1669 ) | ( x18 & n1669 ) ;
  assign n1671 = ( x14 & ~x17 ) | ( x14 & n66 ) | ( ~x17 & n66 ) ;
  assign n1672 = ( ~n66 & n276 ) | ( ~n66 & n1671 ) | ( n276 & n1671 ) ;
  assign n1673 = x13 & n1672 ;
  assign n1674 = x17 & n878 ;
  assign n1675 = n745 & n1674 ;
  assign n1676 = x13 | n1675 ;
  assign n1677 = ~n1673 & n1676 ;
  assign n1678 = ~x16 & n1677 ;
  assign n1679 = ( n1669 & ~n1670 ) | ( n1669 & n1678 ) | ( ~n1670 & n1678 ) ;
  assign n1680 = ( x14 & ~n1664 ) | ( x14 & n1679 ) | ( ~n1664 & n1679 ) ;
  assign n1681 = x13 | n1679 ;
  assign n1682 = ( n1664 & n1680 ) | ( n1664 & n1681 ) | ( n1680 & n1681 ) ;
  assign n1683 = n1660 | n1682 ;
  assign n1684 = ( ~n952 & n1655 ) | ( ~n952 & n1683 ) | ( n1655 & n1683 ) ;
  assign n1685 = ( x12 & x40 ) | ( x12 & n1684 ) | ( x40 & n1684 ) ;
  assign n1686 = ~n1652 & n1685 ;
  assign n1687 = x3 | n1686 ;
  assign n1688 = ( x21 & ~x22 ) | ( x21 & n629 ) | ( ~x22 & n629 ) ;
  assign n1689 = ( x21 & x22 ) | ( x21 & n624 ) | ( x22 & n624 ) ;
  assign n1690 = n1688 & n1689 ;
  assign n1691 = x18 & ~x20 ;
  assign n1692 = ( x19 & n1690 ) | ( x19 & n1691 ) | ( n1690 & n1691 ) ;
  assign n1693 = ~x19 & n1692 ;
  assign n1694 = ( x15 & n84 ) | ( x15 & n1693 ) | ( n84 & n1693 ) ;
  assign n1695 = ~x15 & n1694 ;
  assign n1696 = ( x12 & ~x13 ) | ( x12 & n661 ) | ( ~x13 & n661 ) ;
  assign n1697 = n1695 & ~n1696 ;
  assign n1698 = ( n661 & n1695 ) | ( n661 & ~n1697 ) | ( n1695 & ~n1697 ) ;
  assign n1699 = ~x14 & n1698 ;
  assign n1700 = x3 & ~n1699 ;
  assign n1701 = n1687 & ~n1700 ;
  assign n1702 = x5 | n1701 ;
  assign n1703 = ~x27 & n1357 ;
  assign n1704 = x24 | x27 ;
  assign n1705 = ( ~x24 & n624 ) | ( ~x24 & n1704 ) | ( n624 & n1704 ) ;
  assign n1706 = ~x22 & n1705 ;
  assign n1707 = ( x22 & ~n1366 ) | ( x22 & n1706 ) | ( ~n1366 & n1706 ) ;
  assign n1708 = ( n972 & ~n1357 ) | ( n972 & n1707 ) | ( ~n1357 & n1707 ) ;
  assign n1709 = ( x21 & n1703 ) | ( x21 & ~n1708 ) | ( n1703 & ~n1708 ) ;
  assign n1710 = ( x18 & n1481 ) | ( x18 & ~n1709 ) | ( n1481 & ~n1709 ) ;
  assign n1711 = n1709 & n1710 ;
  assign n1712 = ( x13 & n1436 ) | ( x13 & n1711 ) | ( n1436 & n1711 ) ;
  assign n1713 = ~x13 & n1712 ;
  assign n1714 = ( n578 & ~n1600 ) | ( n578 & n1713 ) | ( ~n1600 & n1713 ) ;
  assign n1715 = ( ~n579 & n1600 ) | ( ~n579 & n1714 ) | ( n1600 & n1714 ) ;
  assign n1716 = x3 & ~n1715 ;
  assign n1717 = ( x13 & x15 ) | ( x13 & n1573 ) | ( x15 & n1573 ) ;
  assign n1718 = x15 | x19 ;
  assign n1719 = ( ~x15 & x18 ) | ( ~x15 & n1718 ) | ( x18 & n1718 ) ;
  assign n1720 = ( ~x17 & x18 ) | ( ~x17 & n1718 ) | ( x18 & n1718 ) ;
  assign n1721 = ( n570 & ~n1719 ) | ( n570 & n1720 ) | ( ~n1719 & n1720 ) ;
  assign n1722 = x16 & n1721 ;
  assign n1723 = x13 & n1722 ;
  assign n1724 = ( ~n1573 & n1717 ) | ( ~n1573 & n1723 ) | ( n1717 & n1723 ) ;
  assign n1725 = ~x12 & n1724 ;
  assign n1726 = x3 | n1725 ;
  assign n1727 = ~n1716 & n1726 ;
  assign n1728 = ~x14 & n1727 ;
  assign n1729 = x5 & ~n1728 ;
  assign n1730 = n1702 & ~n1729 ;
  assign n1731 = x4 | n1730 ;
  assign n1732 = ( ~x4 & n1615 ) | ( ~x4 & n1731 ) | ( n1615 & n1731 ) ;
  assign n1733 = x2 | n1732 ;
  assign n1734 = ~n76 & n153 ;
  assign n1735 = x20 & n1287 ;
  assign n1736 = n1674 & n1735 ;
  assign n1737 = ~x13 & n90 ;
  assign n1738 = ( x3 & ~n76 ) | ( x3 & n1737 ) | ( ~n76 & n1737 ) ;
  assign n1739 = ~x3 & n1738 ;
  assign n1740 = n661 | n1739 ;
  assign n1741 = ( n661 & n1736 ) | ( n661 & n1740 ) | ( n1736 & n1740 ) ;
  assign n1742 = ~x24 & x27 ;
  assign n1743 = ~x19 & n477 ;
  assign n1744 = ~x20 & n1743 ;
  assign n1745 = n1742 & n1744 ;
  assign n1746 = ( x21 & x22 ) | ( x21 & n1745 ) | ( x22 & n1745 ) ;
  assign n1747 = ~x22 & n1746 ;
  assign n1748 = ( ~n275 & n1741 ) | ( ~n275 & n1747 ) | ( n1741 & n1747 ) ;
  assign n1749 = n1734 & ~n1748 ;
  assign n1750 = ( n1734 & n1741 ) | ( n1734 & ~n1749 ) | ( n1741 & ~n1749 ) ;
  assign n1751 = ~x14 & n1750 ;
  assign n1752 = x2 & ~n1751 ;
  assign n1753 = n1733 & ~n1752 ;
  assign n1754 = ( ~x0 & x1 ) | ( ~x0 & n1753 ) | ( x1 & n1753 ) ;
  assign n1755 = n635 & n1078 ;
  assign n1756 = x5 | n123 ;
  assign n1757 = x4 & ~n1756 ;
  assign n1758 = n1755 & ~n1757 ;
  assign n1759 = ( ~x18 & n135 ) | ( ~x18 & n136 ) | ( n135 & n136 ) ;
  assign n1760 = ~n135 & n1759 ;
  assign n1761 = ~x3 & n1760 ;
  assign n1762 = ( x2 & ~x4 ) | ( x2 & n1761 ) | ( ~x4 & n1761 ) ;
  assign n1763 = ~x2 & n1762 ;
  assign n1764 = n140 | n1763 ;
  assign n1765 = ( n1755 & ~n1758 ) | ( n1755 & n1764 ) | ( ~n1758 & n1764 ) ;
  assign n1766 = ( x14 & ~n665 ) | ( x14 & n1765 ) | ( ~n665 & n1765 ) ;
  assign n1767 = n1765 & ~n1766 ;
  assign n1768 = ( x0 & x1 ) | ( x0 & ~n1767 ) | ( x1 & ~n1767 ) ;
  assign n1769 = n1754 & ~n1768 ;
  assign n1770 = ( x3 & ~n129 ) | ( x3 & n165 ) | ( ~n129 & n165 ) ;
  assign n1771 = n70 & n136 ;
  assign n1772 = ( ~x3 & n165 ) | ( ~x3 & n1771 ) | ( n165 & n1771 ) ;
  assign n1773 = ~n1770 & n1772 ;
  assign n1774 = ( ~n129 & n165 ) | ( ~n129 & n1773 ) | ( n165 & n1773 ) ;
  assign n1775 = x16 & n1774 ;
  assign n1776 = ( x4 & n169 ) | ( x4 & ~n1573 ) | ( n169 & ~n1573 ) ;
  assign n1777 = ~x4 & n1776 ;
  assign n1778 = n1775 | n1777 ;
  assign n1779 = ( ~x3 & n1775 ) | ( ~x3 & n1778 ) | ( n1775 & n1778 ) ;
  assign n1780 = ( x14 & ~n665 ) | ( x14 & n1779 ) | ( ~n665 & n1779 ) ;
  assign n1781 = n1779 & ~n1780 ;
  assign n1782 = x0 & ~x2 ;
  assign n1783 = ( x1 & n1781 ) | ( x1 & n1782 ) | ( n1781 & n1782 ) ;
  assign n1784 = ~x1 & n1783 ;
  assign n1785 = ~n1769 & n1784 ;
  assign n1786 = ( ~n848 & n1769 ) | ( ~n848 & n1785 ) | ( n1769 & n1785 ) ;
  assign n1787 = ~x9 & n1786 ;
  assign n1788 = ( x8 & ~x10 ) | ( x8 & n1787 ) | ( ~x10 & n1787 ) ;
  assign n1789 = ~x8 & n1788 ;
  assign n1790 = n153 & n416 ;
  assign n1791 = ( ~n418 & n1674 ) | ( ~n418 & n1790 ) | ( n1674 & n1790 ) ;
  assign n1792 = n665 | n1790 ;
  assign n1793 = ( n418 & n1791 ) | ( n418 & n1792 ) | ( n1791 & n1792 ) ;
  assign n1794 = ( x36 & ~n332 ) | ( x36 & n1793 ) | ( ~n332 & n1793 ) ;
  assign n1795 = n1793 & ~n1794 ;
  assign n1796 = ( x11 & n304 ) | ( x11 & n1795 ) | ( n304 & n1795 ) ;
  assign n1797 = ~x11 & n1796 ;
  assign n1798 = ~x9 & n1797 ;
  assign n1799 = ( x8 & ~x10 ) | ( x8 & n1798 ) | ( ~x10 & n1798 ) ;
  assign n1800 = ~x8 & n1799 ;
  assign n1801 = ~x4 & n1800 ;
  assign n1802 = ( x3 & ~x5 ) | ( x3 & n1801 ) | ( ~x5 & n1801 ) ;
  assign n1803 = ~x3 & n1802 ;
  assign n1804 = ~x1 & n1803 ;
  assign n1805 = ( x0 & ~x2 ) | ( x0 & n1804 ) | ( ~x2 & n1804 ) ;
  assign n1806 = ~x0 & n1805 ;
  assign n1807 = x8 & ~x9 ;
  assign n1808 = ~x36 & n1807 ;
  assign n1809 = ~x4 & n1808 ;
  assign n1810 = ( x3 & ~x5 ) | ( x3 & n1809 ) | ( ~x5 & n1809 ) ;
  assign n1811 = ~x3 & n1810 ;
  assign n1812 = ~x1 & n1811 ;
  assign n1813 = ( x0 & ~x2 ) | ( x0 & n1812 ) | ( ~x2 & n1812 ) ;
  assign n1814 = ~x0 & n1813 ;
  assign n1815 = ~n123 & n515 ;
  assign n1816 = ( x0 & x4 ) | ( x0 & n1815 ) | ( x4 & n1815 ) ;
  assign n1817 = ~x4 & n1816 ;
  assign n1818 = x21 & x22 ;
  assign n1819 = ~x23 & n1742 ;
  assign n1820 = n1818 & n1819 ;
  assign n1821 = n1744 & n1820 ;
  assign n1822 = x13 & x15 ;
  assign n1823 = ~x22 & x24 ;
  assign n1824 = x24 & ~n1823 ;
  assign n1825 = x26 & n1824 ;
  assign n1826 = ( x22 & n1823 ) | ( x22 & ~n1825 ) | ( n1823 & ~n1825 ) ;
  assign n1827 = ( x23 & n1823 ) | ( x23 & n1826 ) | ( n1823 & n1826 ) ;
  assign n1828 = x27 & n1827 ;
  assign n1829 = x22 & ~x23 ;
  assign n1830 = n1041 & ~n1829 ;
  assign n1831 = ~n1828 & n1830 ;
  assign n1832 = ( ~x20 & n918 ) | ( ~x20 & n1323 ) | ( n918 & n1323 ) ;
  assign n1833 = ( n918 & ~n1831 ) | ( n918 & n1832 ) | ( ~n1831 & n1832 ) ;
  assign n1834 = x18 & ~n1833 ;
  assign n1835 = x13 | n1834 ;
  assign n1836 = x12 & n1835 ;
  assign n1837 = ( n1436 & n1822 ) | ( n1436 & ~n1836 ) | ( n1822 & ~n1836 ) ;
  assign n1838 = x5 | n1837 ;
  assign n1839 = x27 & n1357 ;
  assign n1840 = ( x22 & ~x24 ) | ( x22 & x27 ) | ( ~x24 & x27 ) ;
  assign n1841 = ~x22 & n1840 ;
  assign n1842 = ( ~x23 & n1840 ) | ( ~x23 & n1841 ) | ( n1840 & n1841 ) ;
  assign n1843 = ( ~n972 & n1357 ) | ( ~n972 & n1842 ) | ( n1357 & n1842 ) ;
  assign n1844 = ( x21 & n1839 ) | ( x21 & n1843 ) | ( n1839 & n1843 ) ;
  assign n1845 = ~x13 & x18 ;
  assign n1846 = ( x15 & n1844 ) | ( x15 & ~n1845 ) | ( n1844 & ~n1845 ) ;
  assign n1847 = n1844 & ~n1846 ;
  assign n1848 = x12 & n1847 ;
  assign n1849 = x5 & ~n1848 ;
  assign n1850 = n1838 & ~n1849 ;
  assign n1851 = x4 | n1850 ;
  assign n1852 = ~x24 & n1829 ;
  assign n1853 = ~x20 & n1852 ;
  assign n1854 = x21 & n1853 ;
  assign n1855 = ( ~x21 & n1323 ) | ( ~x21 & n1854 ) | ( n1323 & n1854 ) ;
  assign n1856 = ( x5 & n562 ) | ( x5 & ~n1041 ) | ( n562 & ~n1041 ) ;
  assign n1857 = ~x5 & n1856 ;
  assign n1858 = ~n1855 & n1857 ;
  assign n1859 = x18 & x27 ;
  assign n1860 = ( n1855 & n1858 ) | ( n1855 & n1859 ) | ( n1858 & n1859 ) ;
  assign n1861 = ~x13 & n1860 ;
  assign n1862 = ~x15 & n1861 ;
  assign n1863 = x12 & n1862 ;
  assign n1864 = x4 & ~n1863 ;
  assign n1865 = n1851 & ~n1864 ;
  assign n1866 = ( ~x17 & x19 ) | ( ~x17 & n1865 ) | ( x19 & n1865 ) ;
  assign n1867 = x5 | x12 ;
  assign n1868 = n70 & n1822 ;
  assign n1869 = ( x4 & ~n1867 ) | ( x4 & n1868 ) | ( ~n1867 & n1868 ) ;
  assign n1870 = ~x4 & n1869 ;
  assign n1871 = x17 & n1870 ;
  assign n1872 = ( n1865 & ~n1866 ) | ( n1865 & n1871 ) | ( ~n1866 & n1871 ) ;
  assign n1873 = ~x14 & n1872 ;
  assign n1874 = ~x16 & n1873 ;
  assign n1875 = x3 & n1874 ;
  assign n1876 = ~x12 & n487 ;
  assign n1877 = ~x15 & n1330 ;
  assign n1878 = x17 & ~n1877 ;
  assign n1879 = ( n1438 & n1481 ) | ( n1438 & ~n1878 ) | ( n1481 & ~n1878 ) ;
  assign n1880 = ( x5 & ~x15 ) | ( x5 & x17 ) | ( ~x15 & x17 ) ;
  assign n1881 = ( x15 & ~x19 ) | ( x15 & n1880 ) | ( ~x19 & n1880 ) ;
  assign n1882 = ( x5 & x15 ) | ( x5 & ~n1881 ) | ( x15 & ~n1881 ) ;
  assign n1883 = n1880 | n1882 ;
  assign n1884 = ~x19 & n1883 ;
  assign n1885 = ( ~n1881 & n1883 ) | ( ~n1881 & n1884 ) | ( n1883 & n1884 ) ;
  assign n1886 = x40 & ~n1885 ;
  assign n1887 = ( n601 & n1879 ) | ( n601 & n1886 ) | ( n1879 & n1886 ) ;
  assign n1888 = ( x12 & ~x18 ) | ( x12 & n1887 ) | ( ~x18 & n1887 ) ;
  assign n1889 = x5 & ~x19 ;
  assign n1890 = ( x15 & x17 ) | ( x15 & n1889 ) | ( x17 & n1889 ) ;
  assign n1891 = ~x15 & n1890 ;
  assign n1892 = x37 & ~x39 ;
  assign n1893 = ( x17 & ~x37 ) | ( x17 & n1892 ) | ( ~x37 & n1892 ) ;
  assign n1894 = ( ~x15 & x17 ) | ( ~x15 & n1893 ) | ( x17 & n1893 ) ;
  assign n1895 = ( n136 & ~n1893 ) | ( n136 & n1894 ) | ( ~n1893 & n1894 ) ;
  assign n1896 = x19 | n1895 ;
  assign n1897 = ( x15 & x19 ) | ( x15 & n693 ) | ( x19 & n693 ) ;
  assign n1898 = ( x17 & ~x19 ) | ( x17 & n1897 ) | ( ~x19 & n1897 ) ;
  assign n1899 = ( x15 & x17 ) | ( x15 & ~n1897 ) | ( x17 & ~n1897 ) ;
  assign n1900 = n1898 & ~n1899 ;
  assign n1901 = n1562 | n1900 ;
  assign n1902 = ( ~n1895 & n1896 ) | ( ~n1895 & n1901 ) | ( n1896 & n1901 ) ;
  assign n1903 = ( ~x5 & n1891 ) | ( ~x5 & n1902 ) | ( n1891 & n1902 ) ;
  assign n1904 = x40 & ~n1903 ;
  assign n1905 = ( x40 & n1891 ) | ( x40 & ~n1904 ) | ( n1891 & ~n1904 ) ;
  assign n1906 = ( x12 & x18 ) | ( x12 & n1905 ) | ( x18 & n1905 ) ;
  assign n1907 = n1888 & n1906 ;
  assign n1908 = ( ~x18 & n70 ) | ( ~x18 & n693 ) | ( n70 & n693 ) ;
  assign n1909 = ( x17 & n1674 ) | ( x17 & n1908 ) | ( n1674 & n1908 ) ;
  assign n1910 = ~x15 & n1909 ;
  assign n1911 = ( x5 & x12 ) | ( x5 & n1910 ) | ( x12 & n1910 ) ;
  assign n1912 = ~x5 & n1911 ;
  assign n1913 = x15 | n95 ;
  assign n1914 = ( x5 & x12 ) | ( x5 & ~n1913 ) | ( x12 & ~n1913 ) ;
  assign n1915 = ( n325 & n1867 ) | ( n325 & ~n1914 ) | ( n1867 & ~n1914 ) ;
  assign n1916 = n1912 | n1915 ;
  assign n1917 = ( n1002 & n1912 ) | ( n1002 & ~n1916 ) | ( n1912 & ~n1916 ) ;
  assign n1918 = ( ~n1876 & n1907 ) | ( ~n1876 & n1917 ) | ( n1907 & n1917 ) ;
  assign n1919 = x16 & ~n1917 ;
  assign n1920 = ( n1876 & n1918 ) | ( n1876 & ~n1919 ) | ( n1918 & ~n1919 ) ;
  assign n1921 = x14 | n1920 ;
  assign n1922 = n83 & ~n1573 ;
  assign n1923 = ~x17 & n878 ;
  assign n1924 = ( x5 & ~n76 ) | ( x5 & n1923 ) | ( ~n76 & n1923 ) ;
  assign n1925 = ~x5 & n1924 ;
  assign n1926 = x5 & n76 ;
  assign n1927 = ( x5 & n1149 ) | ( x5 & n1926 ) | ( n1149 & n1926 ) ;
  assign n1928 = n1925 | n1927 ;
  assign n1929 = ( n1573 & n1922 ) | ( n1573 & ~n1928 ) | ( n1922 & ~n1928 ) ;
  assign n1930 = ~x12 & n1929 ;
  assign n1931 = x12 & ~n169 ;
  assign n1932 = n1930 | n1931 ;
  assign n1933 = x40 & ~n1932 ;
  assign n1934 = x14 & ~n1933 ;
  assign n1935 = n1921 & ~n1934 ;
  assign n1936 = ( x4 & x13 ) | ( x4 & n1935 ) | ( x13 & n1935 ) ;
  assign n1937 = ~x17 & n76 ;
  assign n1938 = n110 & n1078 ;
  assign n1939 = n1533 | n1938 ;
  assign n1940 = ( n76 & ~n1937 ) | ( n76 & n1939 ) | ( ~n1937 & n1939 ) ;
  assign n1941 = x14 & n1940 ;
  assign n1942 = x12 & n1941 ;
  assign n1943 = ( ~x5 & x40 ) | ( ~x5 & n1942 ) | ( x40 & n1942 ) ;
  assign n1944 = ( x18 & ~n110 ) | ( x18 & n161 ) | ( ~n110 & n161 ) ;
  assign n1945 = x17 & ~n156 ;
  assign n1946 = ( n156 & n1944 ) | ( n156 & ~n1945 ) | ( n1944 & ~n1945 ) ;
  assign n1947 = x12 & n1946 ;
  assign n1948 = x12 | x15 ;
  assign n1949 = ( ~x12 & n1947 ) | ( ~x12 & n1948 ) | ( n1947 & n1948 ) ;
  assign n1950 = x14 & n1949 ;
  assign n1951 = ( x12 & ~x17 ) | ( x12 & x18 ) | ( ~x17 & x18 ) ;
  assign n1952 = ( x12 & x16 ) | ( x12 & x17 ) | ( x16 & x17 ) ;
  assign n1953 = n1951 | n1952 ;
  assign n1954 = x15 & n1953 ;
  assign n1955 = x12 & x29 ;
  assign n1956 = x18 & ~n1643 ;
  assign n1957 = ( ~x17 & x19 ) | ( ~x17 & n1956 ) | ( x19 & n1956 ) ;
  assign n1958 = ( ~n1643 & n1956 ) | ( ~n1643 & n1957 ) | ( n1956 & n1957 ) ;
  assign n1959 = ~x12 & n1958 ;
  assign n1960 = ( x12 & ~n1955 ) | ( x12 & n1959 ) | ( ~n1955 & n1959 ) ;
  assign n1961 = x15 | n1960 ;
  assign n1962 = ( ~x15 & n1954 ) | ( ~x15 & n1961 ) | ( n1954 & n1961 ) ;
  assign n1963 = x14 | n1962 ;
  assign n1964 = ( ~x14 & n1950 ) | ( ~x14 & n1963 ) | ( n1950 & n1963 ) ;
  assign n1965 = ( x5 & x40 ) | ( x5 & n1964 ) | ( x40 & n1964 ) ;
  assign n1966 = n1943 & n1965 ;
  assign n1967 = ( x5 & ~x12 ) | ( x5 & n1966 ) | ( ~x12 & n1966 ) ;
  assign n1968 = n1473 & ~n1967 ;
  assign n1969 = ( n1473 & n1966 ) | ( n1473 & ~n1968 ) | ( n1966 & ~n1968 ) ;
  assign n1970 = x13 & n1969 ;
  assign n1971 = x40 & ~n1970 ;
  assign n1972 = ( x5 & ~n1970 ) | ( x5 & n1971 ) | ( ~n1970 & n1971 ) ;
  assign n1973 = x4 | n1972 ;
  assign n1974 = ( ~n1935 & n1936 ) | ( ~n1935 & n1973 ) | ( n1936 & n1973 ) ;
  assign n1975 = ( ~x19 & n570 ) | ( ~x19 & n1348 ) | ( n570 & n1348 ) ;
  assign n1976 = ~n1348 & n1975 ;
  assign n1977 = ( x12 & x13 ) | ( x12 & x19 ) | ( x13 & x19 ) ;
  assign n1978 = ( x13 & ~x17 ) | ( x13 & n1977 ) | ( ~x17 & n1977 ) ;
  assign n1979 = x13 & ~n1978 ;
  assign n1980 = n1978 | n1979 ;
  assign n1981 = ( ~x13 & n1979 ) | ( ~x13 & n1980 ) | ( n1979 & n1980 ) ;
  assign n1982 = ( x15 & x18 ) | ( x15 & ~n1981 ) | ( x18 & ~n1981 ) ;
  assign n1983 = n418 & n665 ;
  assign n1984 = x15 & n1983 ;
  assign n1985 = ( n1981 & n1982 ) | ( n1981 & n1984 ) | ( n1982 & n1984 ) ;
  assign n1986 = ( x12 & ~x13 ) | ( x12 & n1985 ) | ( ~x13 & n1985 ) ;
  assign n1987 = n1976 & ~n1986 ;
  assign n1988 = ( n1976 & n1985 ) | ( n1976 & ~n1987 ) | ( n1985 & ~n1987 ) ;
  assign n1989 = ( x16 & ~n1199 ) | ( x16 & n1988 ) | ( ~n1199 & n1988 ) ;
  assign n1990 = n1988 & ~n1989 ;
  assign n1991 = n1974 & ~n1990 ;
  assign n1992 = x3 | n1991 ;
  assign n1993 = ~n1875 & n1992 ;
  assign n1994 = x2 | n1993 ;
  assign n1995 = x14 | n76 ;
  assign n1996 = n153 & ~n1995 ;
  assign n1997 = ~n129 & n1996 ;
  assign n1998 = ( x2 & x3 ) | ( x2 & n1997 ) | ( x3 & n1997 ) ;
  assign n1999 = ~x3 & n1998 ;
  assign n2000 = n1994 & ~n1999 ;
  assign n2001 = ( ~n1821 & n1994 ) | ( ~n1821 & n2000 ) | ( n1994 & n2000 ) ;
  assign n2002 = x0 | n2001 ;
  assign n2003 = ~x13 & n85 ;
  assign n2004 = ~n276 & n2003 ;
  assign n2005 = n2002 & ~n2004 ;
  assign n2006 = ( ~n1817 & n2002 ) | ( ~n1817 & n2005 ) | ( n2002 & n2005 ) ;
  assign n2007 = x1 & ~x36 ;
  assign n2008 = ( ~x36 & n2006 ) | ( ~x36 & n2007 ) | ( n2006 & n2007 ) ;
  assign n2009 = x11 & ~n2008 ;
  assign n2010 = x9 | x10 ;
  assign n2011 = ( n2008 & n2009 ) | ( n2008 & ~n2010 ) | ( n2009 & ~n2010 ) ;
  assign n2012 = ~n1814 & n2011 ;
  assign n2013 = ( x8 & ~n1814 ) | ( x8 & n2012 ) | ( ~n1814 & n2012 ) ;
  assign n2014 = ( x15 & x20 ) | ( x15 & x21 ) | ( x20 & x21 ) ;
  assign n2015 = x29 & ~n2014 ;
  assign n2016 = ( x15 & x29 ) | ( x15 & ~n2015 ) | ( x29 & ~n2015 ) ;
  assign n2017 = x14 & ~x18 ;
  assign n2018 = ( ~n190 & n1845 ) | ( ~n190 & n2017 ) | ( n1845 & n2017 ) ;
  assign n2019 = ( x17 & ~n94 ) | ( x17 & n2018 ) | ( ~n94 & n2018 ) ;
  assign n2020 = n2018 & ~n2019 ;
  assign n2021 = ( x13 & ~x14 ) | ( x13 & n2020 ) | ( ~x14 & n2020 ) ;
  assign n2022 = n2016 | n2021 ;
  assign n2023 = ( ~n2016 & n2020 ) | ( ~n2016 & n2022 ) | ( n2020 & n2022 ) ;
  assign n2024 = x12 & ~n2023 ;
  assign n2025 = x13 & n1637 ;
  assign n2026 = x12 | n2025 ;
  assign n2027 = ~n2024 & n2026 ;
  assign n2028 = ( x36 & ~n748 ) | ( x36 & n2027 ) | ( ~n748 & n2027 ) ;
  assign n2029 = n2027 & ~n2028 ;
  assign n2030 = ~x9 & n2029 ;
  assign n2031 = ( x8 & ~x10 ) | ( x8 & n2030 ) | ( ~x10 & n2030 ) ;
  assign n2032 = ~x8 & n2031 ;
  assign n2033 = ~x4 & n2032 ;
  assign n2034 = ( x3 & ~x5 ) | ( x3 & n2033 ) | ( ~x5 & n2033 ) ;
  assign n2035 = ~x3 & n2034 ;
  assign n2036 = ~x1 & n2035 ;
  assign n2037 = ( x0 & ~x2 ) | ( x0 & n2036 ) | ( ~x2 & n2036 ) ;
  assign n2038 = ~x0 & n2037 ;
  assign n2039 = x3 | n1867 ;
  assign n2040 = ( x0 & n1236 ) | ( x0 & ~n2039 ) | ( n1236 & ~n2039 ) ;
  assign n2041 = ~x0 & n2040 ;
  assign n2042 = x13 & n2041 ;
  assign n2043 = ( n43 & n94 ) | ( n43 & n2042 ) | ( n94 & n2042 ) ;
  assign n2044 = ~n43 & n2043 ;
  assign n2045 = ( x18 & n70 ) | ( x18 & n396 ) | ( n70 & n396 ) ;
  assign n2046 = ( x2 & x5 ) | ( x2 & ~n1742 ) | ( x5 & ~n1742 ) ;
  assign n2047 = x2 & n2046 ;
  assign n2048 = ( x40 & n310 ) | ( x40 & ~n2047 ) | ( n310 & ~n2047 ) ;
  assign n2049 = ~n2047 & n2048 ;
  assign n2050 = ~x2 & x23 ;
  assign n2051 = ( x22 & ~n601 ) | ( x22 & n2050 ) | ( ~n601 & n2050 ) ;
  assign n2052 = n601 & n2051 ;
  assign n2053 = n561 & ~n2052 ;
  assign n2054 = ( n2049 & n2052 ) | ( n2049 & ~n2053 ) | ( n2052 & ~n2053 ) ;
  assign n2055 = x20 | n2054 ;
  assign n2056 = ~x2 & n601 ;
  assign n2057 = x20 & ~n2056 ;
  assign n2058 = n2055 & ~n2057 ;
  assign n2059 = x21 & n2058 ;
  assign n2060 = x20 & n601 ;
  assign n2061 = ~x21 & n2060 ;
  assign n2062 = n2059 | n2061 ;
  assign n2063 = ( ~x2 & n2059 ) | ( ~x2 & n2062 ) | ( n2059 & n2062 ) ;
  assign n2064 = x18 & ~n2063 ;
  assign n2065 = x18 | n443 ;
  assign n2066 = ~n2064 & n2065 ;
  assign n2067 = ( ~x17 & x19 ) | ( ~x17 & n2066 ) | ( x19 & n2066 ) ;
  assign n2068 = ~x2 & n1417 ;
  assign n2069 = ~x5 & n2068 ;
  assign n2070 = x17 & n2069 ;
  assign n2071 = ( n2066 & ~n2067 ) | ( n2066 & n2070 ) | ( ~n2067 & n2070 ) ;
  assign n2072 = ( x2 & x5 ) | ( x2 & ~n2071 ) | ( x5 & ~n2071 ) ;
  assign n2073 = n2045 & n2072 ;
  assign n2074 = ( n2045 & n2071 ) | ( n2045 & ~n2073 ) | ( n2071 & ~n2073 ) ;
  assign n2075 = x15 | n2074 ;
  assign n2076 = x5 & x19 ;
  assign n2077 = x17 & ~x40 ;
  assign n2078 = ~x5 & x17 ;
  assign n2079 = ( n2076 & ~n2077 ) | ( n2076 & n2078 ) | ( ~n2077 & n2078 ) ;
  assign n2080 = ( ~x19 & n2076 ) | ( ~x19 & n2079 ) | ( n2076 & n2079 ) ;
  assign n2081 = x18 & ~n2080 ;
  assign n2082 = ( ~x17 & x19 ) | ( ~x17 & x40 ) | ( x19 & x40 ) ;
  assign n2083 = ~x19 & n2082 ;
  assign n2084 = ( x17 & n2082 ) | ( x17 & n2083 ) | ( n2082 & n2083 ) ;
  assign n2085 = ~x5 & n2084 ;
  assign n2086 = x18 | n2085 ;
  assign n2087 = ~n2081 & n2086 ;
  assign n2088 = ~x2 & n2087 ;
  assign n2089 = x15 & ~n2088 ;
  assign n2090 = n2075 & ~n2089 ;
  assign n2091 = x12 & n2090 ;
  assign n2092 = n1876 | n2091 ;
  assign n2093 = ( ~x2 & n2091 ) | ( ~x2 & n2092 ) | ( n2091 & n2092 ) ;
  assign n2094 = ~x16 & n2093 ;
  assign n2095 = n1917 | n2094 ;
  assign n2096 = ( ~x2 & n2094 ) | ( ~x2 & n2095 ) | ( n2094 & n2095 ) ;
  assign n2097 = x13 | n2096 ;
  assign n2098 = ( x5 & x17 ) | ( x5 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n2099 = ( ~x18 & x40 ) | ( ~x18 & n2098 ) | ( x40 & n2098 ) ;
  assign n2100 = n2098 | n2099 ;
  assign n2101 = ~n418 & n2100 ;
  assign n2102 = ( ~x16 & n946 ) | ( ~x16 & n2101 ) | ( n946 & n2101 ) ;
  assign n2103 = x15 & ~n2102 ;
  assign n2104 = ( x15 & n946 ) | ( x15 & ~n2103 ) | ( n946 & ~n2103 ) ;
  assign n2105 = x19 & n2104 ;
  assign n2106 = x19 & n601 ;
  assign n2107 = ~x18 & n2106 ;
  assign n2108 = x15 & n2107 ;
  assign n2109 = ( x16 & x17 ) | ( x16 & n2108 ) | ( x17 & n2108 ) ;
  assign n2110 = ~x17 & n2109 ;
  assign n2111 = x5 & n418 ;
  assign n2112 = ( x15 & x16 ) | ( x15 & n2111 ) | ( x16 & n2111 ) ;
  assign n2113 = ~x16 & n2112 ;
  assign n2114 = ( x15 & x17 ) | ( x15 & x18 ) | ( x17 & x18 ) ;
  assign n2115 = x15 & n2114 ;
  assign n2116 = x15 | x18 ;
  assign n2117 = ( x16 & n2115 ) | ( x16 & ~n2116 ) | ( n2115 & ~n2116 ) ;
  assign n2118 = n2115 | n2117 ;
  assign n2119 = ( ~x5 & n2113 ) | ( ~x5 & n2118 ) | ( n2113 & n2118 ) ;
  assign n2120 = x40 & ~n2119 ;
  assign n2121 = ( x40 & n2113 ) | ( x40 & ~n2120 ) | ( n2113 & ~n2120 ) ;
  assign n2122 = n2110 | n2121 ;
  assign n2123 = ( n2104 & ~n2105 ) | ( n2104 & n2122 ) | ( ~n2105 & n2122 ) ;
  assign n2124 = x12 | n2123 ;
  assign n2125 = ~x22 & x29 ;
  assign n2126 = x23 & n2125 ;
  assign n2127 = ( x40 & n972 ) | ( x40 & ~n2126 ) | ( n972 & ~n2126 ) ;
  assign n2128 = ( n1221 & n2126 ) | ( n1221 & n2127 ) | ( n2126 & n2127 ) ;
  assign n2129 = ~x5 & n2128 ;
  assign n2130 = x12 & ~n2129 ;
  assign n2131 = n2124 & ~n2130 ;
  assign n2132 = ~x2 & n2131 ;
  assign n2133 = x13 & ~n2132 ;
  assign n2134 = n2097 & ~n2133 ;
  assign n2135 = x3 | n2134 ;
  assign n2136 = ( ~x18 & n562 ) | ( ~x18 & n624 ) | ( n562 & n624 ) ;
  assign n2137 = n1829 & ~n2136 ;
  assign n2138 = ( x18 & ~n1829 ) | ( x18 & n2137 ) | ( ~n1829 & n2137 ) ;
  assign n2139 = x13 | n2138 ;
  assign n2140 = x12 & n2139 ;
  assign n2141 = ( n1436 & n1822 ) | ( n1436 & ~n2140 ) | ( n1822 & ~n2140 ) ;
  assign n2142 = ( ~x17 & x19 ) | ( ~x17 & n2141 ) | ( x19 & n2141 ) ;
  assign n2143 = x15 & n70 ;
  assign n2144 = n665 & n2143 ;
  assign n2145 = x17 & n2144 ;
  assign n2146 = ( n2141 & ~n2142 ) | ( n2141 & n2145 ) | ( ~n2142 & n2145 ) ;
  assign n2147 = ~x5 & n2146 ;
  assign n2148 = ~x16 & n2147 ;
  assign n2149 = ~x2 & n2148 ;
  assign n2150 = x3 & ~n2149 ;
  assign n2151 = n2135 & ~n2150 ;
  assign n2152 = ( x0 & ~x1 ) | ( x0 & n2151 ) | ( ~x1 & n2151 ) ;
  assign n2153 = n1079 & ~n1573 ;
  assign n2154 = ~n1082 & n2153 ;
  assign n2155 = ( n665 & n1082 ) | ( n665 & n2154 ) | ( n1082 & n2154 ) ;
  assign n2156 = n1088 & ~n2155 ;
  assign n2157 = ( ~n310 & n2155 ) | ( ~n310 & n2156 ) | ( n2155 & n2156 ) ;
  assign n2158 = ( x0 & x1 ) | ( x0 & ~n2157 ) | ( x1 & ~n2157 ) ;
  assign n2159 = n2152 & ~n2158 ;
  assign n2160 = ( x13 & ~n165 ) | ( x13 & n576 ) | ( ~n165 & n576 ) ;
  assign n2161 = n165 & n2160 ;
  assign n2162 = ~x2 & n2161 ;
  assign n2163 = ( x1 & ~x3 ) | ( x1 & n2162 ) | ( ~x3 & n2162 ) ;
  assign n2164 = ~x1 & n2163 ;
  assign n2165 = x0 & n2164 ;
  assign n2166 = ~x3 & x4 ;
  assign n2167 = ( x13 & n872 ) | ( x13 & n1436 ) | ( n872 & n1436 ) ;
  assign n2168 = ~x13 & n2167 ;
  assign n2169 = ( n578 & ~n1600 ) | ( n578 & n2168 ) | ( ~n1600 & n2168 ) ;
  assign n2170 = ( ~n579 & n1600 ) | ( ~n579 & n2169 ) | ( n1600 & n2169 ) ;
  assign n2171 = ( ~x1 & x2 ) | ( ~x1 & n2170 ) | ( x2 & n2170 ) ;
  assign n2172 = ( x1 & x2 ) | ( x1 & ~n661 ) | ( x2 & ~n661 ) ;
  assign n2173 = n2171 & ~n2172 ;
  assign n2174 = ( x1 & ~n140 ) | ( x1 & n665 ) | ( ~n140 & n665 ) ;
  assign n2175 = n140 & n2174 ;
  assign n2176 = n2173 | n2175 ;
  assign n2177 = ( ~x3 & x4 ) | ( ~x3 & n2176 ) | ( x4 & n2176 ) ;
  assign n2178 = ( n2166 & n2176 ) | ( n2166 & ~n2177 ) | ( n2176 & ~n2177 ) ;
  assign n2179 = ~x17 & n235 ;
  assign n2180 = ( x13 & n66 ) | ( x13 & n2179 ) | ( n66 & n2179 ) ;
  assign n2181 = ~x13 & n2180 ;
  assign n2182 = ( x2 & x17 ) | ( x2 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n2183 = ( ~x2 & x3 ) | ( ~x2 & n2182 ) | ( x3 & n2182 ) ;
  assign n2184 = ( x3 & x17 ) | ( x3 & ~n2182 ) | ( x17 & ~n2182 ) ;
  assign n2185 = n2183 & ~n2184 ;
  assign n2186 = n123 & ~n2185 ;
  assign n2187 = ( n1674 & n2185 ) | ( n1674 & ~n2186 ) | ( n2185 & ~n2186 ) ;
  assign n2188 = ( ~x12 & n2181 ) | ( ~x12 & n2187 ) | ( n2181 & n2187 ) ;
  assign n2189 = x13 & ~n2188 ;
  assign n2190 = ( x13 & n2181 ) | ( x13 & ~n2189 ) | ( n2181 & ~n2189 ) ;
  assign n2191 = ( ~x15 & x16 ) | ( ~x15 & n2190 ) | ( x16 & n2190 ) ;
  assign n2192 = ( x24 & x27 ) | ( x24 & ~n561 ) | ( x27 & ~n561 ) ;
  assign n2193 = ( x3 & ~x27 ) | ( x3 & n2192 ) | ( ~x27 & n2192 ) ;
  assign n2194 = ( x3 & x24 ) | ( x3 & ~n2192 ) | ( x24 & ~n2192 ) ;
  assign n2195 = n2193 & ~n2194 ;
  assign n2196 = ~x3 & x22 ;
  assign n2197 = n629 & n2196 ;
  assign n2198 = ~n2195 & n2197 ;
  assign n2199 = ( n562 & n2195 ) | ( n562 & n2198 ) | ( n2195 & n2198 ) ;
  assign n2200 = x18 & ~n2199 ;
  assign n2201 = x3 | x18 ;
  assign n2202 = ( ~x18 & n2200 ) | ( ~x18 & n2201 ) | ( n2200 & n2201 ) ;
  assign n2203 = ( ~x19 & n570 ) | ( ~x19 & n2202 ) | ( n570 & n2202 ) ;
  assign n2204 = ~n2202 & n2203 ;
  assign n2205 = ~x13 & n2204 ;
  assign n2206 = ( x2 & x12 ) | ( x2 & n2205 ) | ( x12 & n2205 ) ;
  assign n2207 = ~x2 & n2206 ;
  assign n2208 = ~x16 & n2207 ;
  assign n2209 = ( n2190 & ~n2191 ) | ( n2190 & n2208 ) | ( ~n2191 & n2208 ) ;
  assign n2210 = ( x2 & n578 ) | ( x2 & n2209 ) | ( n578 & n2209 ) ;
  assign n2211 = x3 & ~n2210 ;
  assign n2212 = ( x3 & n2209 ) | ( x3 & ~n2211 ) | ( n2209 & ~n2211 ) ;
  assign n2213 = x1 | n2212 ;
  assign n2214 = ( x3 & ~n140 ) | ( x3 & n665 ) | ( ~n140 & n665 ) ;
  assign n2215 = n140 & n2214 ;
  assign n2216 = x2 & n2215 ;
  assign n2217 = x1 & ~n2216 ;
  assign n2218 = n2213 & ~n2217 ;
  assign n2219 = ~x4 & n2218 ;
  assign n2220 = ( x16 & ~n95 ) | ( x16 & n296 ) | ( ~n95 & n296 ) ;
  assign n2221 = x15 & ~n2220 ;
  assign n2222 = x15 | n809 ;
  assign n2223 = ~n2221 & n2222 ;
  assign n2224 = ~x4 & x13 ;
  assign n2225 = ( x12 & n2223 ) | ( x12 & ~n2224 ) | ( n2223 & ~n2224 ) ;
  assign n2226 = n2223 & ~n2225 ;
  assign n2227 = x1 & ~x3 ;
  assign n2228 = ( x2 & n2226 ) | ( x2 & n2227 ) | ( n2226 & n2227 ) ;
  assign n2229 = ~x2 & n2228 ;
  assign n2230 = x13 | n76 ;
  assign n2231 = ( x1 & x12 ) | ( x1 & ~n2230 ) | ( x12 & ~n2230 ) ;
  assign n2232 = ~x1 & n2231 ;
  assign n2233 = ( x1 & x13 ) | ( x1 & n1760 ) | ( x13 & n1760 ) ;
  assign n2234 = x13 & n140 ;
  assign n2235 = ( ~x1 & n2233 ) | ( ~x1 & n2234 ) | ( n2233 & n2234 ) ;
  assign n2236 = ~x12 & n2235 ;
  assign n2237 = n1736 | n2236 ;
  assign n2238 = ( n2232 & n2236 ) | ( n2232 & n2237 ) | ( n2236 & n2237 ) ;
  assign n2239 = ( x2 & x4 ) | ( x2 & n2238 ) | ( x4 & n2238 ) ;
  assign n2240 = ( x3 & ~x4 ) | ( x3 & n2239 ) | ( ~x4 & n2239 ) ;
  assign n2241 = ( x2 & x3 ) | ( x2 & ~n2239 ) | ( x3 & ~n2239 ) ;
  assign n2242 = n2240 & ~n2241 ;
  assign n2243 = n2229 | n2242 ;
  assign n2244 = ( n2218 & ~n2219 ) | ( n2218 & n2243 ) | ( ~n2219 & n2243 ) ;
  assign n2245 = n2178 | n2244 ;
  assign n2246 = ~x0 & n2245 ;
  assign n2247 = n2165 | n2246 ;
  assign n2248 = ( ~n2044 & n2159 ) | ( ~n2044 & n2247 ) | ( n2159 & n2247 ) ;
  assign n2249 = x4 & ~n2247 ;
  assign n2250 = ( n2044 & n2248 ) | ( n2044 & ~n2249 ) | ( n2248 & ~n2249 ) ;
  assign n2251 = ~x14 & n2250 ;
  assign n2252 = ( x4 & ~x5 ) | ( x4 & x40 ) | ( ~x5 & x40 ) ;
  assign n2253 = ( x13 & x18 ) | ( x13 & n76 ) | ( x18 & n76 ) ;
  assign n2254 = ( x12 & ~x13 ) | ( x12 & n2253 ) | ( ~x13 & n2253 ) ;
  assign n2255 = ( x12 & x18 ) | ( x12 & ~n2253 ) | ( x18 & ~n2253 ) ;
  assign n2256 = n2254 & ~n2255 ;
  assign n2257 = x12 | n608 ;
  assign n2258 = n1165 & ~n2257 ;
  assign n2259 = x17 | n2258 ;
  assign n2260 = ( n2256 & n2258 ) | ( n2256 & n2259 ) | ( n2258 & n2259 ) ;
  assign n2261 = ~x5 & n2260 ;
  assign n2262 = ( x15 & ~x16 ) | ( x15 & n1880 ) | ( ~x16 & n1880 ) ;
  assign n2263 = ( x5 & x15 ) | ( x5 & ~n2262 ) | ( x15 & ~n2262 ) ;
  assign n2264 = n1880 & n2263 ;
  assign n2265 = x16 & ~n2264 ;
  assign n2266 = ( n2262 & ~n2264 ) | ( n2262 & n2265 ) | ( ~n2264 & n2265 ) ;
  assign n2267 = ( x12 & ~x18 ) | ( x12 & n2266 ) | ( ~x18 & n2266 ) ;
  assign n2268 = ( ~x13 & x18 ) | ( ~x13 & n2267 ) | ( x18 & n2267 ) ;
  assign n2269 = ( ~x12 & x13 ) | ( ~x12 & n2267 ) | ( x13 & n2267 ) ;
  assign n2270 = n2268 | n2269 ;
  assign n2271 = ( x5 & x12 ) | ( x5 & ~x17 ) | ( x12 & ~x17 ) ;
  assign n2272 = ( ~x12 & x13 ) | ( ~x12 & n2271 ) | ( x13 & n2271 ) ;
  assign n2273 = ( x5 & x13 ) | ( x5 & ~n2271 ) | ( x13 & ~n2271 ) ;
  assign n2274 = n2272 & ~n2273 ;
  assign n2275 = x15 & ~n2274 ;
  assign n2276 = ~x13 & n1276 ;
  assign n2277 = n84 & n2276 ;
  assign n2278 = x15 | n2277 ;
  assign n2279 = ~n2275 & n2278 ;
  assign n2280 = n2270 & ~n2279 ;
  assign n2281 = ( ~n2260 & n2261 ) | ( ~n2260 & n2280 ) | ( n2261 & n2280 ) ;
  assign n2282 = ( ~x12 & x13 ) | ( ~x12 & x15 ) | ( x13 & x15 ) ;
  assign n2283 = x15 & ~n2282 ;
  assign n2284 = ( ~x16 & x17 ) | ( ~x16 & x19 ) | ( x17 & x19 ) ;
  assign n2285 = ( x17 & x18 ) | ( x17 & x19 ) | ( x18 & x19 ) ;
  assign n2286 = n2284 & ~n2285 ;
  assign n2287 = ( x13 & n2283 ) | ( x13 & n2286 ) | ( n2283 & n2286 ) ;
  assign n2288 = ( ~n2282 & n2283 ) | ( ~n2282 & n2287 ) | ( n2283 & n2287 ) ;
  assign n2289 = n878 & ~n2257 ;
  assign n2290 = ~n159 & n2289 ;
  assign n2291 = x5 & x12 ;
  assign n2292 = ( x13 & x15 ) | ( x13 & n2291 ) | ( x15 & n2291 ) ;
  assign n2293 = ~x15 & n2292 ;
  assign n2294 = n127 & n2293 ;
  assign n2295 = ( ~n2288 & n2290 ) | ( ~n2288 & n2294 ) | ( n2290 & n2294 ) ;
  assign n2296 = x5 & ~n2294 ;
  assign n2297 = ( n2288 & n2295 ) | ( n2288 & ~n2296 ) | ( n2295 & ~n2296 ) ;
  assign n2298 = n2281 & n2297 ;
  assign n2299 = ( n239 & ~n2281 ) | ( n239 & n2298 ) | ( ~n2281 & n2298 ) ;
  assign n2300 = ~x4 & n2299 ;
  assign n2301 = ( x5 & n2252 ) | ( x5 & ~n2300 ) | ( n2252 & ~n2300 ) ;
  assign n2302 = x2 | n2301 ;
  assign n2303 = ( ~x1 & x3 ) | ( ~x1 & n2302 ) | ( x3 & n2302 ) ;
  assign n2304 = x1 | n2303 ;
  assign n2305 = ~n2251 & n2304 ;
  assign n2306 = ( x0 & ~n2251 ) | ( x0 & n2305 ) | ( ~n2251 & n2305 ) ;
  assign n2307 = x36 & n2306 ;
  assign n2308 = x10 | x11 ;
  assign n2309 = ( n2306 & ~n2307 ) | ( n2306 & n2308 ) | ( ~n2307 & n2308 ) ;
  assign n2310 = x0 | x1 ;
  assign n2311 = n129 | n2310 ;
  assign n2312 = ( n123 & n1808 ) | ( n123 & ~n2311 ) | ( n1808 & ~n2311 ) ;
  assign n2313 = ~n123 & n2312 ;
  assign n2314 = ( ~x9 & x10 ) | ( ~x9 & n2313 ) | ( x10 & n2313 ) ;
  assign n2315 = x8 & ~n2313 ;
  assign n2316 = ( x9 & n2314 ) | ( x9 & ~n2315 ) | ( n2314 & ~n2315 ) ;
  assign n2317 = ( x8 & x9 ) | ( x8 & ~n2316 ) | ( x9 & ~n2316 ) ;
  assign n2318 = ~n2309 & n2317 ;
  assign n2319 = ( n2309 & ~n2316 ) | ( n2309 & n2318 ) | ( ~n2316 & n2318 ) ;
  assign n2320 = x13 & n1779 ;
  assign n2321 = ~x12 & n2320 ;
  assign n2322 = ~x1 & n2321 ;
  assign n2323 = ~x2 & n2322 ;
  assign n2324 = x0 & n2323 ;
  assign n2325 = x3 & n661 ;
  assign n2326 = ~x22 & n1742 ;
  assign n2327 = n562 & n2326 ;
  assign n2328 = n153 & n2327 ;
  assign n2329 = ( x15 & n477 ) | ( x15 & n2328 ) | ( n477 & n2328 ) ;
  assign n2330 = ~x15 & n2329 ;
  assign n2331 = ( ~x5 & n1600 ) | ( ~x5 & n2330 ) | ( n1600 & n2330 ) ;
  assign n2332 = x20 & x27 ;
  assign n2333 = ( x18 & x21 ) | ( x18 & n2332 ) | ( x21 & n2332 ) ;
  assign n2334 = ~x21 & n2333 ;
  assign n2335 = n570 & n2334 ;
  assign n2336 = n153 & n2335 ;
  assign n2337 = ( x5 & n1600 ) | ( x5 & n2336 ) | ( n1600 & n2336 ) ;
  assign n2338 = n2331 | n2337 ;
  assign n2339 = ( x16 & x19 ) | ( x16 & n2338 ) | ( x19 & n2338 ) ;
  assign n2340 = x15 & n1078 ;
  assign n2341 = ( x12 & x13 ) | ( x12 & n2340 ) | ( x13 & n2340 ) ;
  assign n2342 = ~x12 & n2341 ;
  assign n2343 = ~x16 & n2342 ;
  assign n2344 = ( n2338 & ~n2339 ) | ( n2338 & n2343 ) | ( ~n2339 & n2343 ) ;
  assign n2345 = n578 | n2344 ;
  assign n2346 = ~x3 & n2345 ;
  assign n2347 = n2325 | n2346 ;
  assign n2348 = x2 & n2347 ;
  assign n2349 = x3 | x5 ;
  assign n2350 = ( ~x17 & n1311 ) | ( ~x17 & n2349 ) | ( n1311 & n2349 ) ;
  assign n2351 = x3 & x18 ;
  assign n2352 = ( ~x5 & x18 ) | ( ~x5 & n601 ) | ( x18 & n601 ) ;
  assign n2353 = ( x3 & x18 ) | ( x3 & n2352 ) | ( x18 & n2352 ) ;
  assign n2354 = ( n2351 & n2352 ) | ( n2351 & ~n2353 ) | ( n2352 & ~n2353 ) ;
  assign n2355 = x19 & n2354 ;
  assign n2356 = x17 & n2355 ;
  assign n2357 = ( n1311 & ~n2350 ) | ( n1311 & n2356 ) | ( ~n2350 & n2356 ) ;
  assign n2358 = ( x3 & ~x17 ) | ( x3 & n1312 ) | ( ~x17 & n1312 ) ;
  assign n2359 = ~x3 & n2358 ;
  assign n2360 = ~n2357 & n2359 ;
  assign n2361 = x13 & x16 ;
  assign n2362 = ( n2357 & n2360 ) | ( n2357 & n2361 ) | ( n2360 & n2361 ) ;
  assign n2363 = ( x12 & ~x15 ) | ( x12 & n2362 ) | ( ~x15 & n2362 ) ;
  assign n2364 = ~x29 & x40 ;
  assign n2365 = ( x5 & x13 ) | ( x5 & n2364 ) | ( x13 & n2364 ) ;
  assign n2366 = ~x5 & n2365 ;
  assign n2367 = x3 & n2366 ;
  assign n2368 = x13 & x40 ;
  assign n2369 = ( x5 & x29 ) | ( x5 & n2368 ) | ( x29 & n2368 ) ;
  assign n2370 = ~x5 & n2369 ;
  assign n2371 = ( x3 & ~x20 ) | ( x3 & n2370 ) | ( ~x20 & n2370 ) ;
  assign n2372 = x21 & ~n1053 ;
  assign n2373 = ( x21 & n1828 ) | ( x21 & n2372 ) | ( n1828 & n2372 ) ;
  assign n2374 = x17 & n2373 ;
  assign n2375 = ( x18 & x19 ) | ( x18 & n2374 ) | ( x19 & n2374 ) ;
  assign n2376 = ~x19 & n2375 ;
  assign n2377 = x5 & ~x16 ;
  assign n2378 = ( x13 & n2376 ) | ( x13 & n2377 ) | ( n2376 & n2377 ) ;
  assign n2379 = ~x13 & n2378 ;
  assign n2380 = ( x3 & x20 ) | ( x3 & ~n2379 ) | ( x20 & ~n2379 ) ;
  assign n2381 = n2371 & ~n2380 ;
  assign n2382 = ( x22 & x23 ) | ( x22 & x40 ) | ( x23 & x40 ) ;
  assign n2383 = ~x21 & x40 ;
  assign n2384 = ( ~x22 & n2382 ) | ( ~x22 & n2383 ) | ( n2382 & n2383 ) ;
  assign n2385 = x29 & n2384 ;
  assign n2386 = ( x5 & x13 ) | ( x5 & n2385 ) | ( x13 & n2385 ) ;
  assign n2387 = ~x5 & n2386 ;
  assign n2388 = ( x3 & x20 ) | ( x3 & n2387 ) | ( x20 & n2387 ) ;
  assign n2389 = ( x3 & x13 ) | ( x3 & n2377 ) | ( x13 & n2377 ) ;
  assign n2390 = ~x13 & n2389 ;
  assign n2391 = x19 | x27 ;
  assign n2392 = x21 | n2391 ;
  assign n2393 = n477 & ~n2392 ;
  assign n2394 = n2390 & n2393 ;
  assign n2395 = x20 & n2394 ;
  assign n2396 = ( ~x3 & n2388 ) | ( ~x3 & n2395 ) | ( n2388 & n2395 ) ;
  assign n2397 = n2381 | n2396 ;
  assign n2398 = ( n2366 & ~n2367 ) | ( n2366 & n2397 ) | ( ~n2367 & n2397 ) ;
  assign n2399 = ( x12 & x15 ) | ( x12 & ~n2398 ) | ( x15 & ~n2398 ) ;
  assign n2400 = n2363 & ~n2399 ;
  assign n2401 = x3 & ~n1416 ;
  assign n2402 = ( ~n95 & n1416 ) | ( ~n95 & n2401 ) | ( n1416 & n2401 ) ;
  assign n2403 = x16 & n2402 ;
  assign n2404 = x18 & n1416 ;
  assign n2405 = ( x3 & x17 ) | ( x3 & n2404 ) | ( x17 & n2404 ) ;
  assign n2406 = ~x3 & n2405 ;
  assign n2407 = x3 & ~n1310 ;
  assign n2408 = ( ~n95 & n1310 ) | ( ~n95 & n2407 ) | ( n1310 & n2407 ) ;
  assign n2409 = n2406 | n2408 ;
  assign n2410 = ~x16 & n2409 ;
  assign n2411 = n2403 | n2410 ;
  assign n2412 = x5 | n2411 ;
  assign n2413 = ( x3 & x16 ) | ( x3 & x19 ) | ( x16 & x19 ) ;
  assign n2414 = ( x18 & n134 ) | ( x18 & ~n2413 ) | ( n134 & ~n2413 ) ;
  assign n2415 = x17 | n2414 ;
  assign n2416 = x5 & n2415 ;
  assign n2417 = n2412 & ~n2416 ;
  assign n2418 = ~x12 & x15 ;
  assign n2419 = ( x13 & ~n2417 ) | ( x13 & n2418 ) | ( ~n2417 & n2418 ) ;
  assign n2420 = n2417 & n2419 ;
  assign n2421 = n2400 | n2420 ;
  assign n2422 = ~x2 & n2421 ;
  assign n2423 = n2348 | n2422 ;
  assign n2424 = ( ~x1 & x4 ) | ( ~x1 & n2423 ) | ( x4 & n2423 ) ;
  assign n2425 = ( x1 & x4 ) | ( x1 & ~n661 ) | ( x4 & ~n661 ) ;
  assign n2426 = n2424 & ~n2425 ;
  assign n2427 = n667 | n2426 ;
  assign n2428 = ~x0 & n2427 ;
  assign n2429 = n2324 | n2428 ;
  assign n2430 = ( x14 & x36 ) | ( x14 & n2429 ) | ( x36 & n2429 ) ;
  assign n2431 = ( x15 & n277 ) | ( x15 & n1661 ) | ( n277 & n1661 ) ;
  assign n2432 = x14 & ~x17 ;
  assign n2433 = ( x16 & n2431 ) | ( x16 & n2432 ) | ( n2431 & n2432 ) ;
  assign n2434 = ~x16 & n2433 ;
  assign n2435 = x13 & n2434 ;
  assign n2436 = ( x5 & x12 ) | ( x5 & n2435 ) | ( x12 & n2435 ) ;
  assign n2437 = ~x5 & n2436 ;
  assign n2438 = ~x3 & n2437 ;
  assign n2439 = ( x2 & ~x4 ) | ( x2 & n2438 ) | ( ~x4 & n2438 ) ;
  assign n2440 = ~x2 & n2439 ;
  assign n2441 = ~x0 & n2440 ;
  assign n2442 = ~x1 & n2441 ;
  assign n2443 = ~x36 & n2442 ;
  assign n2444 = ( n2429 & ~n2430 ) | ( n2429 & n2443 ) | ( ~n2430 & n2443 ) ;
  assign n2445 = ~x10 & n2444 ;
  assign n2446 = ( x9 & ~x11 ) | ( x9 & n2445 ) | ( ~x11 & n2445 ) ;
  assign n2447 = ~x9 & n2446 ;
  assign n2448 = ~x8 & n2447 ;
  assign n2449 = ( x16 & ~x17 ) | ( x16 & x18 ) | ( ~x17 & x18 ) ;
  assign n2450 = ( x16 & x18 ) | ( x16 & ~n2449 ) | ( x18 & ~n2449 ) ;
  assign n2451 = ( x15 & ~x17 ) | ( x15 & n2450 ) | ( ~x17 & n2450 ) ;
  assign n2452 = ~x13 & x40 ;
  assign n2453 = ( x19 & ~n2451 ) | ( x19 & n2452 ) | ( ~n2451 & n2452 ) ;
  assign n2454 = n2451 & n2453 ;
  assign n2455 = ( x3 & n515 ) | ( x3 & n2454 ) | ( n515 & n2454 ) ;
  assign n2456 = ~x3 & n2455 ;
  assign n2457 = x2 & n2456 ;
  assign n2458 = x2 | n601 ;
  assign n2459 = x3 | n2458 ;
  assign n2460 = ( x18 & ~n136 ) | ( x18 & n2459 ) | ( ~n136 & n2459 ) ;
  assign n2461 = n2459 & ~n2460 ;
  assign n2462 = n559 & n2461 ;
  assign n2463 = n136 & n244 ;
  assign n2464 = ( x5 & ~n1709 ) | ( x5 & n2351 ) | ( ~n1709 & n2351 ) ;
  assign n2465 = n1709 & n2464 ;
  assign n2466 = ( x2 & x17 ) | ( x2 & n2465 ) | ( x17 & n2465 ) ;
  assign n2467 = ~x2 & x18 ;
  assign n2468 = x18 & ~n2467 ;
  assign n2469 = n1735 & n2468 ;
  assign n2470 = ( x40 & ~n2467 ) | ( x40 & n2468 ) | ( ~n2467 & n2468 ) ;
  assign n2471 = ( ~x2 & n2469 ) | ( ~x2 & n2470 ) | ( n2469 & n2470 ) ;
  assign n2472 = ~x5 & n2471 ;
  assign n2473 = ~x3 & n2472 ;
  assign n2474 = x17 & n2473 ;
  assign n2475 = ( ~x2 & n2466 ) | ( ~x2 & n2474 ) | ( n2466 & n2474 ) ;
  assign n2476 = ~x15 & n2475 ;
  assign n2477 = x2 | n2349 ;
  assign n2478 = ~n2476 & n2477 ;
  assign n2479 = ( n2463 & n2476 ) | ( n2463 & ~n2478 ) | ( n2476 & ~n2478 ) ;
  assign n2480 = ( ~n558 & n559 ) | ( ~n558 & n2479 ) | ( n559 & n2479 ) ;
  assign n2481 = ( x12 & n2462 ) | ( x12 & n2480 ) | ( n2462 & n2480 ) ;
  assign n2482 = ( x16 & ~x19 ) | ( x16 & n2481 ) | ( ~x19 & n2481 ) ;
  assign n2483 = x2 & n1600 ;
  assign n2484 = ( x5 & ~x15 ) | ( x5 & n1270 ) | ( ~x15 & n1270 ) ;
  assign n2485 = ( x5 & ~x40 ) | ( x5 & n1270 ) | ( ~x40 & n1270 ) ;
  assign n2486 = ( x40 & ~n2484 ) | ( x40 & n2485 ) | ( ~n2484 & n2485 ) ;
  assign n2487 = ( ~x13 & x17 ) | ( ~x13 & n2486 ) | ( x17 & n2486 ) ;
  assign n2488 = x40 & ~n2349 ;
  assign n2489 = ( x15 & x17 ) | ( x15 & n2488 ) | ( x17 & n2488 ) ;
  assign n2490 = ~x15 & n2489 ;
  assign n2491 = x13 & n2490 ;
  assign n2492 = ( n2486 & ~n2487 ) | ( n2486 & n2491 ) | ( ~n2487 & n2491 ) ;
  assign n2493 = ~x12 & n2492 ;
  assign n2494 = ( x17 & x40 ) | ( x17 & n618 ) | ( x40 & n618 ) ;
  assign n2495 = ( ~n618 & n1221 ) | ( ~n618 & n2494 ) | ( n1221 & n2494 ) ;
  assign n2496 = ~x13 & n2495 ;
  assign n2497 = ( x5 & x12 ) | ( x5 & n2496 ) | ( x12 & n2496 ) ;
  assign n2498 = ~x5 & n2497 ;
  assign n2499 = n2493 | n2498 ;
  assign n2500 = ( ~x3 & n2493 ) | ( ~x3 & n2499 ) | ( n2493 & n2499 ) ;
  assign n2501 = ~x18 & n2500 ;
  assign n2502 = ( x15 & ~n185 ) | ( x15 & n244 ) | ( ~n185 & n244 ) ;
  assign n2503 = ~x13 & n2502 ;
  assign n2504 = ( x5 & x12 ) | ( x5 & n2503 ) | ( x12 & n2503 ) ;
  assign n2505 = ~x5 & n2504 ;
  assign n2506 = n2501 | n2505 ;
  assign n2507 = ( ~x3 & n2501 ) | ( ~x3 & n2506 ) | ( n2501 & n2506 ) ;
  assign n2508 = x2 | n2507 ;
  assign n2509 = ( ~x2 & n2483 ) | ( ~x2 & n2508 ) | ( n2483 & n2508 ) ;
  assign n2510 = ( x16 & x19 ) | ( x16 & ~n2509 ) | ( x19 & ~n2509 ) ;
  assign n2511 = n2482 & ~n2510 ;
  assign n2512 = x19 & n479 ;
  assign n2513 = ~x12 & n2512 ;
  assign n2514 = ( ~x2 & x13 ) | ( ~x2 & n2513 ) | ( x13 & n2513 ) ;
  assign n2515 = ( x16 & x17 ) | ( x16 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n2516 = ( ~x17 & n133 ) | ( ~x17 & n2515 ) | ( n133 & n2515 ) ;
  assign n2517 = ~x12 & n2516 ;
  assign n2518 = ~x22 & x23 ;
  assign n2519 = x21 & x29 ;
  assign n2520 = ( x22 & n2518 ) | ( x22 & n2519 ) | ( n2518 & n2519 ) ;
  assign n2521 = x20 & n2520 ;
  assign n2522 = x12 & ~n2521 ;
  assign n2523 = n2517 | n2522 ;
  assign n2524 = ~x15 & n2523 ;
  assign n2525 = ( x17 & ~x18 ) | ( x17 & x19 ) | ( ~x18 & x19 ) ;
  assign n2526 = ~x17 & n2525 ;
  assign n2527 = ( ~x16 & x18 ) | ( ~x16 & n2526 ) | ( x18 & n2526 ) ;
  assign n2528 = ( n2525 & n2526 ) | ( n2525 & n2527 ) | ( n2526 & n2527 ) ;
  assign n2529 = ~x12 & n2528 ;
  assign n2530 = x15 & ~n2529 ;
  assign n2531 = n2524 | n2530 ;
  assign n2532 = x40 & ~n2531 ;
  assign n2533 = ( x5 & n1270 ) | ( x5 & ~n2513 ) | ( n1270 & ~n2513 ) ;
  assign n2534 = ( x5 & n1270 ) | ( x5 & ~n2532 ) | ( n1270 & ~n2532 ) ;
  assign n2535 = ( n2532 & ~n2533 ) | ( n2532 & n2534 ) | ( ~n2533 & n2534 ) ;
  assign n2536 = ( x2 & x13 ) | ( x2 & n2535 ) | ( x13 & n2535 ) ;
  assign n2537 = n2514 & n2536 ;
  assign n2538 = n2511 | n2537 ;
  assign n2539 = ( n2456 & ~n2457 ) | ( n2456 & n2538 ) | ( ~n2457 & n2538 ) ;
  assign n2540 = ( ~x1 & x4 ) | ( ~x1 & n2539 ) | ( x4 & n2539 ) ;
  assign n2541 = x3 & n443 ;
  assign n2542 = ( n661 & n1734 ) | ( n661 & n1747 ) | ( n1734 & n1747 ) ;
  assign n2543 = n2541 & ~n2542 ;
  assign n2544 = ( n661 & n2541 ) | ( n661 & ~n2543 ) | ( n2541 & ~n2543 ) ;
  assign n2545 = ( x1 & x4 ) | ( x1 & ~n2544 ) | ( x4 & ~n2544 ) ;
  assign n2546 = n2540 & ~n2545 ;
  assign n2547 = ( ~x13 & x16 ) | ( ~x13 & x17 ) | ( x16 & x17 ) ;
  assign n2548 = n66 & n2547 ;
  assign n2549 = ( x13 & n66 ) | ( x13 & ~n2548 ) | ( n66 & ~n2548 ) ;
  assign n2550 = ~x12 & n2549 ;
  assign n2551 = ~x18 & n1643 ;
  assign n2552 = ( x17 & ~x19 ) | ( x17 & n2551 ) | ( ~x19 & n2551 ) ;
  assign n2553 = ( n1643 & n2551 ) | ( n1643 & n2552 ) | ( n2551 & n2552 ) ;
  assign n2554 = n127 | n2553 ;
  assign n2555 = x13 & ~n2554 ;
  assign n2556 = x12 & ~n2555 ;
  assign n2557 = n2550 | n2556 ;
  assign n2558 = ( x15 & ~x40 ) | ( x15 & n2557 ) | ( ~x40 & n2557 ) ;
  assign n2559 = n1165 & ~n1437 ;
  assign n2560 = ( x12 & x16 ) | ( x12 & ~x17 ) | ( x16 & ~x17 ) ;
  assign n2561 = ( ~x12 & x13 ) | ( ~x12 & n2560 ) | ( x13 & n2560 ) ;
  assign n2562 = ( ~x13 & x17 ) | ( ~x13 & n2560 ) | ( x17 & n2560 ) ;
  assign n2563 = n2561 & n2562 ;
  assign n2564 = ~x15 & n2563 ;
  assign n2565 = x12 | x13 ;
  assign n2566 = ( x12 & ~x15 ) | ( x12 & x17 ) | ( ~x15 & x17 ) ;
  assign n2567 = ( x13 & ~x15 ) | ( x13 & n2566 ) | ( ~x15 & n2566 ) ;
  assign n2568 = ( x15 & ~n2565 ) | ( x15 & n2567 ) | ( ~n2565 & n2567 ) ;
  assign n2569 = n2564 | n2568 ;
  assign n2570 = ( n1165 & ~n2559 ) | ( n1165 & n2569 ) | ( ~n2559 & n2569 ) ;
  assign n2571 = x40 & n2570 ;
  assign n2572 = ( n2557 & ~n2558 ) | ( n2557 & n2571 ) | ( ~n2558 & n2571 ) ;
  assign n2573 = ( x4 & n1029 ) | ( x4 & n2572 ) | ( n1029 & n2572 ) ;
  assign n2574 = ~x4 & n2573 ;
  assign n2575 = ~x2 & n2574 ;
  assign n2576 = ( x1 & ~x3 ) | ( x1 & n2575 ) | ( ~x3 & n2575 ) ;
  assign n2577 = ~x1 & n2576 ;
  assign n2578 = ( ~n667 & n2546 ) | ( ~n667 & n2577 ) | ( n2546 & n2577 ) ;
  assign n2579 = x14 & ~n2577 ;
  assign n2580 = ( n667 & n2578 ) | ( n667 & ~n2579 ) | ( n2578 & ~n2579 ) ;
  assign n2581 = x0 | n2580 ;
  assign n2582 = ( x4 & n169 ) | ( x4 & n1078 ) | ( n169 & n1078 ) ;
  assign n2583 = ~x4 & n2582 ;
  assign n2584 = x16 & n501 ;
  assign n2585 = ( x16 & n2583 ) | ( x16 & n2584 ) | ( n2583 & n2584 ) ;
  assign n2586 = n1777 & ~n2585 ;
  assign n2587 = ( n215 & n2585 ) | ( n215 & n2586 ) | ( n2585 & n2586 ) ;
  assign n2588 = ~x3 & n2587 ;
  assign n2589 = ( x2 & ~x12 ) | ( x2 & n2588 ) | ( ~x12 & n2588 ) ;
  assign n2590 = ~x2 & n2589 ;
  assign n2591 = ~x1 & n2590 ;
  assign n2592 = x0 & ~n2591 ;
  assign n2593 = n2581 & ~n2592 ;
  assign n2594 = ( x11 & n391 ) | ( x11 & n2593 ) | ( n391 & n2593 ) ;
  assign n2595 = n2593 & ~n2594 ;
  assign n2596 = ~x8 & n2595 ;
  assign n2597 = ~x9 & n2596 ;
  assign n2598 = x11 & n1111 ;
  assign n2599 = x1 & ~x10 ;
  assign n2600 = ( x8 & n1767 ) | ( x8 & n2599 ) | ( n1767 & n2599 ) ;
  assign n2601 = ~x8 & n2600 ;
  assign n2602 = x13 & ~x18 ;
  assign n2603 = ~x13 & x19 ;
  assign n2604 = x12 & ~n2603 ;
  assign n2605 = ( n1442 & n2602 ) | ( n1442 & ~n2604 ) | ( n2602 & ~n2604 ) ;
  assign n2606 = x15 & n2605 ;
  assign n2607 = ~x17 & n2606 ;
  assign n2608 = x13 | n1348 ;
  assign n2609 = x12 & n2608 ;
  assign n2610 = ( n1436 & n1822 ) | ( n1436 & ~n2609 ) | ( n1822 & ~n2609 ) ;
  assign n2611 = ( ~x17 & x19 ) | ( ~x17 & n2610 ) | ( x19 & n2610 ) ;
  assign n2612 = ( n2145 & n2610 ) | ( n2145 & ~n2611 ) | ( n2610 & ~n2611 ) ;
  assign n2613 = ( n578 & ~n2607 ) | ( n578 & n2612 ) | ( ~n2607 & n2612 ) ;
  assign n2614 = ( ~n579 & n2607 ) | ( ~n579 & n2613 ) | ( n2607 & n2613 ) ;
  assign n2615 = ~x14 & n2614 ;
  assign n2616 = x4 & ~x10 ;
  assign n2617 = ( x8 & n2615 ) | ( x8 & n2616 ) | ( n2615 & n2616 ) ;
  assign n2618 = ~x8 & n2617 ;
  assign n2619 = x37 | x39 ;
  assign n2620 = x38 | n2619 ;
  assign n2621 = x19 & ~n2620 ;
  assign n2622 = ( ~n95 & n2620 ) | ( ~n95 & n2621 ) | ( n2620 & n2621 ) ;
  assign n2623 = ( x12 & x16 ) | ( x12 & n2622 ) | ( x16 & n2622 ) ;
  assign n2624 = ( ~x16 & n558 ) | ( ~x16 & n2623 ) | ( n558 & n2623 ) ;
  assign n2625 = ( x12 & x13 ) | ( x12 & ~n159 ) | ( x13 & ~n159 ) ;
  assign n2626 = ( x12 & x13 ) | ( x12 & x18 ) | ( x13 & x18 ) ;
  assign n2627 = x13 | n2626 ;
  assign n2628 = ( x12 & ~n2620 ) | ( x12 & n2626 ) | ( ~n2620 & n2626 ) ;
  assign n2629 = x13 & n2628 ;
  assign n2630 = n2627 & ~n2629 ;
  assign n2631 = ( x16 & n2625 ) | ( x16 & ~n2630 ) | ( n2625 & ~n2630 ) ;
  assign n2632 = ~x17 & n2631 ;
  assign n2633 = ( x17 & n2625 ) | ( x17 & n2632 ) | ( n2625 & n2632 ) ;
  assign n2634 = ( x18 & ~n1328 ) | ( x18 & n1481 ) | ( ~n1328 & n1481 ) ;
  assign n2635 = n1328 & n2634 ;
  assign n2636 = x24 & x28 ;
  assign n2637 = ( ~x13 & x25 ) | ( ~x13 & n2636 ) | ( x25 & n2636 ) ;
  assign n2638 = x13 & n2637 ;
  assign n2639 = ( x13 & x16 ) | ( x13 & ~n2638 ) | ( x16 & ~n2638 ) ;
  assign n2640 = n2635 & n2639 ;
  assign n2641 = ( n2635 & n2638 ) | ( n2635 & ~n2640 ) | ( n2638 & ~n2640 ) ;
  assign n2642 = x23 & n1818 ;
  assign n2643 = ( x20 & n624 ) | ( x20 & n2642 ) | ( n624 & n2642 ) ;
  assign n2644 = ~x20 & n2643 ;
  assign n2645 = ~x16 & n2644 ;
  assign n2646 = ( x13 & n1674 ) | ( x13 & n2645 ) | ( n1674 & n2645 ) ;
  assign n2647 = ~x13 & n2646 ;
  assign n2648 = ( x13 & ~x24 ) | ( x13 & n2647 ) | ( ~x24 & n2647 ) ;
  assign n2649 = x28 & ~n2648 ;
  assign n2650 = ( x28 & n2647 ) | ( x28 & ~n2649 ) | ( n2647 & ~n2649 ) ;
  assign n2651 = ( ~x22 & x24 ) | ( ~x22 & n1364 ) | ( x24 & n1364 ) ;
  assign n2652 = x22 & n2651 ;
  assign n2653 = ( x19 & ~x20 ) | ( x19 & n2652 ) | ( ~x20 & n2652 ) ;
  assign n2654 = x19 | x21 ;
  assign n2655 = ( x20 & n2653 ) | ( x20 & n2654 ) | ( n2653 & n2654 ) ;
  assign n2656 = n369 & ~n2655 ;
  assign n2657 = ( x13 & x24 ) | ( x13 & x25 ) | ( x24 & x25 ) ;
  assign n2658 = x13 & ~x28 ;
  assign n2659 = ( ~x25 & n2657 ) | ( ~x25 & n2658 ) | ( n2657 & n2658 ) ;
  assign n2660 = ( ~x17 & n2656 ) | ( ~x17 & n2659 ) | ( n2656 & n2659 ) ;
  assign n2661 = x13 & ~n2659 ;
  assign n2662 = ( n2656 & ~n2660 ) | ( n2656 & n2661 ) | ( ~n2660 & n2661 ) ;
  assign n2663 = ( x12 & n2650 ) | ( x12 & ~n2662 ) | ( n2650 & ~n2662 ) ;
  assign n2664 = ~n2641 & n2663 ;
  assign n2665 = ( x12 & n2641 ) | ( x12 & n2664 ) | ( n2641 & n2664 ) ;
  assign n2666 = ( x15 & n1948 ) | ( x15 & ~n2665 ) | ( n1948 & ~n2665 ) ;
  assign n2667 = ( n2624 & n2633 ) | ( n2624 & n2666 ) | ( n2633 & n2666 ) ;
  assign n2668 = ~x15 & n2666 ;
  assign n2669 = ( ~n2624 & n2667 ) | ( ~n2624 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2670 = ~x14 & n2669 ;
  assign n2671 = ( x8 & ~x40 ) | ( x8 & n2670 ) | ( ~x40 & n2670 ) ;
  assign n2672 = ~x8 & x10 ;
  assign n2673 = ( n2670 & ~n2671 ) | ( n2670 & n2672 ) | ( ~n2671 & n2672 ) ;
  assign n2674 = ( x4 & x5 ) | ( x4 & ~n2673 ) | ( x5 & ~n2673 ) ;
  assign n2675 = x16 | n1718 ;
  assign n2676 = ( x12 & x14 ) | ( x12 & ~x40 ) | ( x14 & ~x40 ) ;
  assign n2677 = x14 & ~n2676 ;
  assign n2678 = ( x12 & n635 ) | ( x12 & n2677 ) | ( n635 & n2677 ) ;
  assign n2679 = ( ~n2676 & n2677 ) | ( ~n2676 & n2678 ) | ( n2677 & n2678 ) ;
  assign n2680 = ( x12 & ~x14 ) | ( x12 & n2679 ) | ( ~x14 & n2679 ) ;
  assign n2681 = n2675 | n2680 ;
  assign n2682 = ( ~n2675 & n2679 ) | ( ~n2675 & n2681 ) | ( n2679 & n2681 ) ;
  assign n2683 = ~x18 & n2682 ;
  assign n2684 = x12 & x14 ;
  assign n2685 = x14 & ~n2684 ;
  assign n2686 = x40 & n2685 ;
  assign n2687 = ~x19 & n1330 ;
  assign n2688 = ( ~n2684 & n2685 ) | ( ~n2684 & n2687 ) | ( n2685 & n2687 ) ;
  assign n2689 = ( x12 & n2686 ) | ( x12 & n2688 ) | ( n2686 & n2688 ) ;
  assign n2690 = ( x15 & ~x16 ) | ( x15 & n2689 ) | ( ~x16 & n2689 ) ;
  assign n2691 = ( x12 & x19 ) | ( x12 & n2677 ) | ( x19 & n2677 ) ;
  assign n2692 = ( ~n2676 & n2677 ) | ( ~n2676 & n2691 ) | ( n2677 & n2691 ) ;
  assign n2693 = ( x15 & x16 ) | ( x15 & ~n2692 ) | ( x16 & ~n2692 ) ;
  assign n2694 = n2690 & ~n2693 ;
  assign n2695 = ( x12 & x15 ) | ( x12 & n2677 ) | ( x15 & n2677 ) ;
  assign n2696 = ( ~n2676 & n2677 ) | ( ~n2676 & n2695 ) | ( n2677 & n2695 ) ;
  assign n2697 = x16 & n2696 ;
  assign n2698 = n2694 | n2697 ;
  assign n2699 = x18 & n2698 ;
  assign n2700 = n2683 | n2699 ;
  assign n2701 = x17 & n2700 ;
  assign n2702 = ~x16 & n66 ;
  assign n2703 = x12 & n2702 ;
  assign n2704 = n304 & n2703 ;
  assign n2705 = x40 | n2704 ;
  assign n2706 = ( n1524 & n2704 ) | ( n1524 & n2705 ) | ( n2704 & n2705 ) ;
  assign n2707 = x17 | n2706 ;
  assign n2708 = ( ~x17 & n2701 ) | ( ~x17 & n2707 ) | ( n2701 & n2707 ) ;
  assign n2709 = ~x13 & n2708 ;
  assign n2710 = ( x40 & n797 ) | ( x40 & n1221 ) | ( n797 & n1221 ) ;
  assign n2711 = x12 & x17 ;
  assign n2712 = ( x14 & ~n2710 ) | ( x14 & n2711 ) | ( ~n2710 & n2711 ) ;
  assign n2713 = n2710 & n2712 ;
  assign n2714 = x15 & ~n373 ;
  assign n2715 = ~n796 & n2714 ;
  assign n2716 = ~x12 & n1116 ;
  assign n2717 = n304 & n2716 ;
  assign n2718 = x16 & n745 ;
  assign n2719 = ( x12 & ~n244 ) | ( x12 & n2718 ) | ( ~n244 & n2718 ) ;
  assign n2720 = n244 & n2719 ;
  assign n2721 = n2717 | n2720 ;
  assign n2722 = ( ~n2713 & n2715 ) | ( ~n2713 & n2721 ) | ( n2715 & n2721 ) ;
  assign n2723 = n2713 | n2722 ;
  assign n2724 = ( x15 & x18 ) | ( x15 & ~x19 ) | ( x18 & ~x19 ) ;
  assign n2725 = ( ~x15 & x16 ) | ( ~x15 & n2724 ) | ( x16 & n2724 ) ;
  assign n2726 = ( x18 & ~x19 ) | ( x18 & n2725 ) | ( ~x19 & n2725 ) ;
  assign n2727 = ~n2724 & n2726 ;
  assign n2728 = ( ~n2725 & n2726 ) | ( ~n2725 & n2727 ) | ( n2726 & n2727 ) ;
  assign n2729 = ~x12 & x17 ;
  assign n2730 = ( x14 & n2728 ) | ( x14 & ~n2729 ) | ( n2728 & ~n2729 ) ;
  assign n2731 = n2728 & ~n2730 ;
  assign n2732 = x14 & n110 ;
  assign n2733 = x12 & n2732 ;
  assign n2734 = ( ~n95 & n2731 ) | ( ~n95 & n2733 ) | ( n2731 & n2733 ) ;
  assign n2735 = n1416 & ~n2734 ;
  assign n2736 = ( n1416 & n2731 ) | ( n1416 & ~n2735 ) | ( n2731 & ~n2735 ) ;
  assign n2737 = n2723 | n2736 ;
  assign n2738 = x13 & n2737 ;
  assign n2739 = n2709 | n2738 ;
  assign n2740 = x5 & ~x8 ;
  assign n2741 = ( x10 & n2739 ) | ( x10 & ~n2740 ) | ( n2739 & ~n2740 ) ;
  assign n2742 = n2739 & ~n2741 ;
  assign n2743 = ~x4 & n2742 ;
  assign n2744 = ( n2673 & n2674 ) | ( n2673 & ~n2743 ) | ( n2674 & ~n2743 ) ;
  assign n2745 = ~x12 & n1822 ;
  assign n2746 = ( x4 & ~x19 ) | ( x4 & n2745 ) | ( ~x19 & n2745 ) ;
  assign n2747 = ( x4 & x15 ) | ( x4 & ~x18 ) | ( x15 & ~x18 ) ;
  assign n2748 = x21 & n1046 ;
  assign n2749 = ~x20 & n2748 ;
  assign n2750 = ( x15 & x18 ) | ( x15 & ~n2749 ) | ( x18 & ~n2749 ) ;
  assign n2751 = n2747 | n2750 ;
  assign n2752 = x13 | n2751 ;
  assign n2753 = x12 & ~n2752 ;
  assign n2754 = ~x19 & n2753 ;
  assign n2755 = ( ~x4 & n2746 ) | ( ~x4 & n2754 ) | ( n2746 & n2754 ) ;
  assign n2756 = x15 & n665 ;
  assign n2757 = ( x4 & n70 ) | ( x4 & n2756 ) | ( n70 & n2756 ) ;
  assign n2758 = ~x4 & n2757 ;
  assign n2759 = ~n2755 & n2758 ;
  assign n2760 = ( n84 & n2755 ) | ( n84 & n2759 ) | ( n2755 & n2759 ) ;
  assign n2761 = ( x5 & ~x14 ) | ( x5 & n2760 ) | ( ~x14 & n2760 ) ;
  assign n2762 = ( x21 & n561 ) | ( x21 & ~n1705 ) | ( n561 & ~n1705 ) ;
  assign n2763 = x21 & n1366 ;
  assign n2764 = ( ~n561 & n2762 ) | ( ~n561 & n2763 ) | ( n2762 & n2763 ) ;
  assign n2765 = ( ~x19 & x20 ) | ( ~x19 & n2764 ) | ( x20 & n2764 ) ;
  assign n2766 = ~x19 & n1061 ;
  assign n2767 = ( ~x20 & n2765 ) | ( ~x20 & n2766 ) | ( n2765 & n2766 ) ;
  assign n2768 = x18 & n2767 ;
  assign n2769 = ( x15 & x17 ) | ( x15 & n2768 ) | ( x17 & n2768 ) ;
  assign n2770 = ~x15 & n2769 ;
  assign n2771 = ~x13 & n2770 ;
  assign n2772 = ( x4 & x12 ) | ( x4 & n2771 ) | ( x12 & n2771 ) ;
  assign n2773 = ~x4 & n2772 ;
  assign n2774 = ( n573 & n578 ) | ( n573 & ~n2773 ) | ( n578 & ~n2773 ) ;
  assign n2775 = ( ~n579 & n2773 ) | ( ~n579 & n2774 ) | ( n2773 & n2774 ) ;
  assign n2776 = ~x14 & n2775 ;
  assign n2777 = ( ~x5 & n2761 ) | ( ~x5 & n2776 ) | ( n2761 & n2776 ) ;
  assign n2778 = x3 & ~x10 ;
  assign n2779 = ( x8 & n2777 ) | ( x8 & n2778 ) | ( n2777 & n2778 ) ;
  assign n2780 = ~x8 & n2779 ;
  assign n2781 = ( n2618 & n2744 ) | ( n2618 & ~n2780 ) | ( n2744 & ~n2780 ) ;
  assign n2782 = x3 & ~n2780 ;
  assign n2783 = ( ~n2618 & n2781 ) | ( ~n2618 & n2782 ) | ( n2781 & n2782 ) ;
  assign n2784 = ( x1 & x2 ) | ( x1 & ~n2783 ) | ( x2 & ~n2783 ) ;
  assign n2785 = ( x19 & n562 ) | ( x19 & n1360 ) | ( n562 & n1360 ) ;
  assign n2786 = ~x19 & n2785 ;
  assign n2787 = x18 & n2786 ;
  assign n2788 = ( x16 & x17 ) | ( x16 & n2787 ) | ( x17 & n2787 ) ;
  assign n2789 = ~x16 & n2788 ;
  assign n2790 = ( x13 & n1436 ) | ( x13 & n2789 ) | ( n1436 & n2789 ) ;
  assign n2791 = ~x13 & n2790 ;
  assign n2792 = ~x4 & n2791 ;
  assign n2793 = ( x3 & ~x5 ) | ( x3 & n2792 ) | ( ~x5 & n2792 ) ;
  assign n2794 = ~x3 & n2793 ;
  assign n2795 = ~x14 & n1741 ;
  assign n2796 = ( ~x14 & n2794 ) | ( ~x14 & n2795 ) | ( n2794 & n2795 ) ;
  assign n2797 = x2 & ~x10 ;
  assign n2798 = ( x8 & n2796 ) | ( x8 & n2797 ) | ( n2796 & n2797 ) ;
  assign n2799 = ~x8 & n2798 ;
  assign n2800 = ~x1 & n2799 ;
  assign n2801 = ( n2783 & n2784 ) | ( n2783 & ~n2800 ) | ( n2784 & ~n2800 ) ;
  assign n2802 = ~x14 & n158 ;
  assign n2803 = ( ~x14 & n2321 ) | ( ~x14 & n2802 ) | ( n2321 & n2802 ) ;
  assign n2804 = ~x8 & n2803 ;
  assign n2805 = ( x2 & ~x10 ) | ( x2 & n2804 ) | ( ~x10 & n2804 ) ;
  assign n2806 = ~x2 & n2805 ;
  assign n2807 = ~x1 & n2806 ;
  assign n2808 = x0 & n2807 ;
  assign n2809 = ( n2601 & n2801 ) | ( n2601 & ~n2808 ) | ( n2801 & ~n2808 ) ;
  assign n2810 = x0 & ~n2808 ;
  assign n2811 = ( ~n2601 & n2809 ) | ( ~n2601 & n2810 ) | ( n2809 & n2810 ) ;
  assign n2812 = ( x11 & x36 ) | ( x11 & ~n2811 ) | ( x36 & ~n2811 ) ;
  assign n2813 = ~x8 & x36 ;
  assign n2814 = ( ~x8 & x10 ) | ( ~x8 & n2813 ) | ( x10 & n2813 ) ;
  assign n2815 = ~x11 & n2814 ;
  assign n2816 = ( n2811 & n2812 ) | ( n2811 & ~n2815 ) | ( n2812 & ~n2815 ) ;
  assign n2817 = x9 & ~x11 ;
  assign n2818 = ( x8 & x10 ) | ( x8 & n2817 ) | ( x10 & n2817 ) ;
  assign n2819 = ~x8 & n2818 ;
  assign n2820 = ( n2598 & n2816 ) | ( n2598 & ~n2819 ) | ( n2816 & ~n2819 ) ;
  assign n2821 = x9 & ~n2819 ;
  assign n2822 = ( ~n2598 & n2820 ) | ( ~n2598 & n2821 ) | ( n2820 & n2821 ) ;
  assign n2823 = x9 & ~x10 ;
  assign n2824 = x9 & ~n2823 ;
  assign n2825 = ~x11 & n2824 ;
  assign n2826 = ~x38 & x40 ;
  assign n2827 = ( x39 & n1496 ) | ( x39 & ~n2826 ) | ( n1496 & ~n2826 ) ;
  assign n2828 = n1496 & ~n2827 ;
  assign n2829 = ~x36 & n2828 ;
  assign n2830 = ( x17 & ~x37 ) | ( x17 & n2829 ) | ( ~x37 & n2829 ) ;
  assign n2831 = ~x17 & n2830 ;
  assign n2832 = ~x16 & n2831 ;
  assign n2833 = ( x14 & x15 ) | ( x14 & n2832 ) | ( x15 & n2832 ) ;
  assign n2834 = ~x14 & n2833 ;
  assign n2835 = ~x10 & n2834 ;
  assign n2836 = ~x11 & n2835 ;
  assign n2837 = ~x4 & n2836 ;
  assign n2838 = ( x3 & ~x5 ) | ( x3 & n2837 ) | ( ~x5 & n2837 ) ;
  assign n2839 = ~x3 & n2838 ;
  assign n2840 = ~x1 & n2839 ;
  assign n2841 = ( x0 & ~x2 ) | ( x0 & n2840 ) | ( ~x2 & n2840 ) ;
  assign n2842 = ~x0 & n2841 ;
  assign n2843 = ( n2823 & ~n2824 ) | ( n2823 & n2842 ) | ( ~n2824 & n2842 ) ;
  assign n2844 = ( x10 & ~n2825 ) | ( x10 & n2843 ) | ( ~n2825 & n2843 ) ;
  assign n2845 = ~x8 & n2844 ;
  assign n2846 = ~x1 & n2803 ;
  assign n2847 = ~x2 & n2846 ;
  assign n2848 = x0 & n2847 ;
  assign n2849 = x3 & n2777 ;
  assign n2850 = x4 & n2615 ;
  assign n2851 = ( x12 & ~x19 ) | ( x12 & n1822 ) | ( ~x19 & n1822 ) ;
  assign n2852 = x18 | n1330 ;
  assign n2853 = ( n608 & ~n1330 ) | ( n608 & n2852 ) | ( ~n1330 & n2852 ) ;
  assign n2854 = ( x12 & x19 ) | ( x12 & n2853 ) | ( x19 & n2853 ) ;
  assign n2855 = n2851 & ~n2854 ;
  assign n2856 = n2144 | n2855 ;
  assign n2857 = ( x16 & ~x17 ) | ( x16 & n2856 ) | ( ~x17 & n2856 ) ;
  assign n2858 = ~x16 & n2607 ;
  assign n2859 = ( n2856 & ~n2857 ) | ( n2856 & n2858 ) | ( ~n2857 & n2858 ) ;
  assign n2860 = ( ~x12 & n1722 ) | ( ~x12 & n2859 ) | ( n1722 & n2859 ) ;
  assign n2861 = x13 & ~n2860 ;
  assign n2862 = ( x13 & n2859 ) | ( x13 & ~n2861 ) | ( n2859 & ~n2861 ) ;
  assign n2863 = ( x14 & ~n601 ) | ( x14 & n2862 ) | ( ~n601 & n2862 ) ;
  assign n2864 = ( x15 & x17 ) | ( x15 & ~n66 ) | ( x17 & ~n66 ) ;
  assign n2865 = ( n66 & n635 ) | ( n66 & n2864 ) | ( n635 & n2864 ) ;
  assign n2866 = ~x13 & n2865 ;
  assign n2867 = x12 & n2866 ;
  assign n2868 = ( ~x5 & x40 ) | ( ~x5 & n2867 ) | ( x40 & n2867 ) ;
  assign n2869 = ~x13 & x17 ;
  assign n2870 = ( ~x13 & x16 ) | ( ~x13 & n2869 ) | ( x16 & n2869 ) ;
  assign n2871 = n66 & n2729 ;
  assign n2872 = x13 & n2871 ;
  assign n2873 = ( x17 & x18 ) | ( x17 & n474 ) | ( x18 & n474 ) ;
  assign n2874 = ~x13 & n2873 ;
  assign n2875 = ( x12 & n2872 ) | ( x12 & ~n2874 ) | ( n2872 & ~n2874 ) ;
  assign n2876 = x16 | n2875 ;
  assign n2877 = x16 & ~n558 ;
  assign n2878 = n2876 & ~n2877 ;
  assign n2879 = ( x12 & n2870 ) | ( x12 & n2878 ) | ( n2870 & n2878 ) ;
  assign n2880 = ( x13 & x17 ) | ( x13 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n2881 = ~n2547 & n2880 ;
  assign n2882 = ( x12 & ~n2878 ) | ( x12 & n2881 ) | ( ~n2878 & n2881 ) ;
  assign n2883 = ~n2879 & n2882 ;
  assign n2884 = x15 & ~n2883 ;
  assign n2885 = x13 | n952 ;
  assign n2886 = ( ~n126 & n952 ) | ( ~n126 & n2885 ) | ( n952 & n2885 ) ;
  assign n2887 = ~n952 & n2886 ;
  assign n2888 = ( ~x13 & n2361 ) | ( ~x13 & n2887 ) | ( n2361 & n2887 ) ;
  assign n2889 = x12 | n2888 ;
  assign n2890 = x16 & x19 ;
  assign n2891 = ( x16 & x19 ) | ( x16 & ~n77 ) | ( x19 & ~n77 ) ;
  assign n2892 = ( n84 & ~n2890 ) | ( n84 & n2891 ) | ( ~n2890 & n2891 ) ;
  assign n2893 = ~x39 & n418 ;
  assign n2894 = n2892 & n2893 ;
  assign n2895 = ( ~n135 & n2892 ) | ( ~n135 & n2894 ) | ( n2892 & n2894 ) ;
  assign n2896 = ~x13 & n2895 ;
  assign n2897 = x12 & ~n2896 ;
  assign n2898 = n2889 & ~n2897 ;
  assign n2899 = ~x15 & n2898 ;
  assign n2900 = ( x15 & ~n2884 ) | ( x15 & n2899 ) | ( ~n2884 & n2899 ) ;
  assign n2901 = ( x5 & x40 ) | ( x5 & ~n2900 ) | ( x40 & ~n2900 ) ;
  assign n2902 = n2868 & n2901 ;
  assign n2903 = ~x14 & n2902 ;
  assign n2904 = ( n2862 & ~n2863 ) | ( n2862 & n2903 ) | ( ~n2863 & n2903 ) ;
  assign n2905 = x5 & ~x40 ;
  assign n2906 = ( ~x12 & x13 ) | ( ~x12 & n2566 ) | ( x13 & n2566 ) ;
  assign n2907 = ( ~x13 & x15 ) | ( ~x13 & n2566 ) | ( x15 & n2566 ) ;
  assign n2908 = n2906 & n2907 ;
  assign n2909 = ( x5 & ~x12 ) | ( x5 & x13 ) | ( ~x12 & x13 ) ;
  assign n2910 = ( x13 & ~x15 ) | ( x13 & n2909 ) | ( ~x15 & n2909 ) ;
  assign n2911 = n2909 & n2910 ;
  assign n2912 = n153 | n2911 ;
  assign n2913 = ( ~n2564 & n2908 ) | ( ~n2564 & n2912 ) | ( n2908 & n2912 ) ;
  assign n2914 = ~x5 & n2912 ;
  assign n2915 = ( ~n2908 & n2913 ) | ( ~n2908 & n2914 ) | ( n2913 & n2914 ) ;
  assign n2916 = x5 & n1533 ;
  assign n2917 = n558 & n2916 ;
  assign n2918 = ( x5 & x12 ) | ( x5 & x13 ) | ( x12 & x13 ) ;
  assign n2919 = ( n2294 & n2565 ) | ( n2294 & ~n2918 ) | ( n2565 & ~n2918 ) ;
  assign n2920 = n2917 | n2919 ;
  assign n2921 = n2915 & ~n2920 ;
  assign n2922 = x14 & ~n2921 ;
  assign n2923 = x40 & ~n2922 ;
  assign n2924 = n2905 | n2923 ;
  assign n2925 = ~n2904 & n2924 ;
  assign n2926 = x4 | n2925 ;
  assign n2927 = ~n2850 & n2926 ;
  assign n2928 = ~x3 & n2927 ;
  assign n2929 = ( x3 & ~n2849 ) | ( x3 & n2928 ) | ( ~n2849 & n2928 ) ;
  assign n2930 = ( x1 & ~x2 ) | ( x1 & n2929 ) | ( ~x2 & n2929 ) ;
  assign n2931 = ( x1 & x2 ) | ( x1 & ~n2796 ) | ( x2 & ~n2796 ) ;
  assign n2932 = n2930 | n2931 ;
  assign n2933 = x1 & n1767 ;
  assign n2934 = n2932 & ~n2933 ;
  assign n2935 = x0 | n2934 ;
  assign n2936 = ~n2848 & n2935 ;
  assign n2937 = ~x36 & n2936 ;
  assign n2938 = x11 & ~n2937 ;
  assign n2939 = ( ~n2010 & n2937 ) | ( ~n2010 & n2938 ) | ( n2937 & n2938 ) ;
  assign n2940 = ~n1814 & n2939 ;
  assign n2941 = ( x8 & ~n1814 ) | ( x8 & n2940 ) | ( ~n1814 & n2940 ) ;
  assign n2942 = x19 & n196 ;
  assign n2943 = ~x16 & n2942 ;
  assign n2944 = ( x15 & ~x18 ) | ( x15 & n2943 ) | ( ~x18 & n2943 ) ;
  assign n2945 = ~x15 & n2944 ;
  assign n2946 = ( x13 & n383 ) | ( x13 & n2945 ) | ( n383 & n2945 ) ;
  assign n2947 = ~x13 & n2946 ;
  assign n2948 = ~x10 & n2947 ;
  assign n2949 = ~x11 & n2948 ;
  assign n2950 = ~x8 & n2949 ;
  assign n2951 = ( x5 & ~x9 ) | ( x5 & n2950 ) | ( ~x9 & n2950 ) ;
  assign n2952 = ~x5 & n2951 ;
  assign n2953 = ~x3 & n2952 ;
  assign n2954 = ( x2 & ~x4 ) | ( x2 & n2953 ) | ( ~x4 & n2953 ) ;
  assign n2955 = ~x2 & n2954 ;
  assign n2956 = ~x0 & n2955 ;
  assign n2957 = ~x1 & n2956 ;
  assign n2958 = ~x4 & n2949 ;
  assign n2959 = ( x3 & ~x5 ) | ( x3 & n2958 ) | ( ~x5 & n2958 ) ;
  assign n2960 = ~x3 & n2959 ;
  assign n2961 = ~x1 & n2960 ;
  assign n2962 = ( x0 & ~x2 ) | ( x0 & n2961 ) | ( ~x2 & n2961 ) ;
  assign n2963 = ~x0 & n2962 ;
  assign n2964 = x10 & ~n2963 ;
  assign n2965 = x8 | x9 ;
  assign n2966 = ( n2963 & n2964 ) | ( n2963 & ~n2965 ) | ( n2964 & ~n2965 ) ;
  assign n2967 = x17 | n373 ;
  assign n2968 = x13 | n2967 ;
  assign n2969 = ( ~x12 & n1573 ) | ( ~x12 & n2968 ) | ( n1573 & n2968 ) ;
  assign n2970 = n1573 & ~n2969 ;
  assign n2971 = ( n2666 & n2668 ) | ( n2666 & n2970 ) | ( n2668 & n2970 ) ;
  assign n2972 = ~x14 & n2971 ;
  assign n2973 = ( x8 & ~x40 ) | ( x8 & n2972 ) | ( ~x40 & n2972 ) ;
  assign n2974 = ( n2672 & n2972 ) | ( n2672 & ~n2973 ) | ( n2972 & ~n2973 ) ;
  assign n2975 = ( x4 & x5 ) | ( x4 & ~n2974 ) | ( x5 & ~n2974 ) ;
  assign n2976 = ( ~n2743 & n2974 ) | ( ~n2743 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2977 = ( n2618 & ~n2780 ) | ( n2618 & n2976 ) | ( ~n2780 & n2976 ) ;
  assign n2978 = ( ~n2618 & n2782 ) | ( ~n2618 & n2977 ) | ( n2782 & n2977 ) ;
  assign n2979 = ( x1 & x2 ) | ( x1 & ~n2978 ) | ( x2 & ~n2978 ) ;
  assign n2980 = ( ~n2800 & n2978 ) | ( ~n2800 & n2979 ) | ( n2978 & n2979 ) ;
  assign n2981 = ( n2601 & ~n2808 ) | ( n2601 & n2980 ) | ( ~n2808 & n2980 ) ;
  assign n2982 = ( ~n2601 & n2810 ) | ( ~n2601 & n2981 ) | ( n2810 & n2981 ) ;
  assign n2983 = ( x11 & x36 ) | ( x11 & ~n2982 ) | ( x36 & ~n2982 ) ;
  assign n2984 = ( ~n2815 & n2982 ) | ( ~n2815 & n2983 ) | ( n2982 & n2983 ) ;
  assign n2985 = ( n2598 & ~n2819 ) | ( n2598 & n2984 ) | ( ~n2819 & n2984 ) ;
  assign n2986 = ( ~n2598 & n2821 ) | ( ~n2598 & n2985 ) | ( n2821 & n2985 ) ;
  assign n2987 = ( ~x8 & x9 ) | ( ~x8 & x10 ) | ( x9 & x10 ) ;
  assign n2988 = ( x8 & x9 ) | ( x8 & ~x11 ) | ( x9 & ~x11 ) ;
  assign n2989 = n2987 & ~n2988 ;
  assign n2990 = ( ~x10 & n2987 ) | ( ~x10 & n2989 ) | ( n2987 & n2989 ) ;
  assign n2991 = ( x15 & ~x40 ) | ( x15 & n1132 ) | ( ~x40 & n1132 ) ;
  assign n2992 = ( x15 & x40 ) | ( x15 & n66 ) | ( x40 & n66 ) ;
  assign n2993 = ~n2991 & n2992 ;
  assign n2994 = ~x17 & n2993 ;
  assign n2995 = ( x16 & ~x36 ) | ( x16 & n2994 ) | ( ~x36 & n2994 ) ;
  assign n2996 = ~x16 & n2995 ;
  assign n2997 = ( x13 & n383 ) | ( x13 & n2996 ) | ( n383 & n2996 ) ;
  assign n2998 = ~x13 & n2997 ;
  assign n2999 = ~x10 & n2998 ;
  assign n3000 = ( x5 & ~x11 ) | ( x5 & n2999 ) | ( ~x11 & n2999 ) ;
  assign n3001 = ~x5 & n3000 ;
  assign n3002 = ~x3 & n3001 ;
  assign n3003 = ( x2 & ~x4 ) | ( x2 & n3002 ) | ( ~x4 & n3002 ) ;
  assign n3004 = ~x2 & n3003 ;
  assign n3005 = ( x0 & x1 ) | ( x0 & ~x10 ) | ( x1 & ~x10 ) ;
  assign n3006 = n3004 & n3005 ;
  assign n3007 = ( x10 & n3004 ) | ( x10 & ~n3006 ) | ( n3004 & ~n3006 ) ;
  assign n3008 = ( x8 & x9 ) | ( x8 & n3007 ) | ( x9 & n3007 ) ;
  assign n3009 = ( n728 & n3007 ) | ( n728 & ~n3008 ) | ( n3007 & ~n3008 ) ;
  assign n3010 = ~x10 & x36 ;
  assign n3011 = ( x8 & ~x11 ) | ( x8 & n3010 ) | ( ~x11 & n3010 ) ;
  assign n3012 = ~x8 & n3011 ;
  assign n3013 = ~x10 & n1767 ;
  assign n3014 = ( x8 & ~x11 ) | ( x8 & n3013 ) | ( ~x11 & n3013 ) ;
  assign n3015 = ~x8 & n3014 ;
  assign n3016 = x1 & n3015 ;
  assign n3017 = ~x10 & n2796 ;
  assign n3018 = ( x8 & ~x11 ) | ( x8 & n3017 ) | ( ~x11 & n3017 ) ;
  assign n3019 = ~x8 & n3018 ;
  assign n3020 = x2 & n3019 ;
  assign n3021 = ~x10 & n2615 ;
  assign n3022 = ( x8 & ~x11 ) | ( x8 & n3021 ) | ( ~x11 & n3021 ) ;
  assign n3023 = ~x8 & n3022 ;
  assign n3024 = x4 & n3023 ;
  assign n3025 = ( x12 & n1253 ) | ( x12 & n2626 ) | ( n1253 & n2626 ) ;
  assign n3026 = x13 & n3025 ;
  assign n3027 = n2627 & ~n3026 ;
  assign n3028 = ( x16 & n2625 ) | ( x16 & ~n3027 ) | ( n2625 & ~n3027 ) ;
  assign n3029 = ~x17 & n3028 ;
  assign n3030 = ( x17 & n2625 ) | ( x17 & n3029 ) | ( n2625 & n3029 ) ;
  assign n3031 = ( x13 & n1573 ) | ( x13 & ~n3030 ) | ( n1573 & ~n3030 ) ;
  assign n3032 = ~x12 & n3030 ;
  assign n3033 = ( n1573 & ~n3031 ) | ( n1573 & n3032 ) | ( ~n3031 & n3032 ) ;
  assign n3034 = ( ~x14 & x15 ) | ( ~x14 & n3033 ) | ( x15 & n3033 ) ;
  assign n3035 = x14 | n2666 ;
  assign n3036 = ( n3033 & ~n3034 ) | ( n3033 & n3035 ) | ( ~n3034 & n3035 ) ;
  assign n3037 = ( x11 & ~x14 ) | ( x11 & n3036 ) | ( ~x14 & n3036 ) ;
  assign n3038 = x40 & ~n3037 ;
  assign n3039 = ( x11 & x40 ) | ( x11 & ~n3038 ) | ( x40 & ~n3038 ) ;
  assign n3040 = ( x5 & ~x10 ) | ( x5 & n3039 ) | ( ~x10 & n3039 ) ;
  assign n3041 = ( x10 & ~n1103 ) | ( x10 & n3040 ) | ( ~n1103 & n3040 ) ;
  assign n3042 = x8 | x11 ;
  assign n3043 = ( x10 & n2739 ) | ( x10 & n3042 ) | ( n2739 & n3042 ) ;
  assign n3044 = n2739 & ~n3043 ;
  assign n3045 = x5 & n3044 ;
  assign n3046 = n3041 & ~n3045 ;
  assign n3047 = x4 | n3046 ;
  assign n3048 = ~n3024 & n3047 ;
  assign n3049 = ( x2 & ~x3 ) | ( x2 & n3048 ) | ( ~x3 & n3048 ) ;
  assign n3050 = ~x10 & n2777 ;
  assign n3051 = ( x8 & ~x11 ) | ( x8 & n3050 ) | ( ~x11 & n3050 ) ;
  assign n3052 = ~x8 & n3051 ;
  assign n3053 = ( x2 & x3 ) | ( x2 & ~n3052 ) | ( x3 & ~n3052 ) ;
  assign n3054 = n3049 | n3053 ;
  assign n3055 = ~n3020 & n3054 ;
  assign n3056 = x1 | n3055 ;
  assign n3057 = ~n3016 & n3056 ;
  assign n3058 = ( x0 & x36 ) | ( x0 & ~n3057 ) | ( x36 & ~n3057 ) ;
  assign n3059 = ~x10 & n2803 ;
  assign n3060 = ( x8 & ~x11 ) | ( x8 & n3059 ) | ( ~x11 & n3059 ) ;
  assign n3061 = ~x8 & n3060 ;
  assign n3062 = ( x1 & n1782 ) | ( x1 & n3061 ) | ( n1782 & n3061 ) ;
  assign n3063 = ~x1 & n3062 ;
  assign n3064 = ~x36 & n3063 ;
  assign n3065 = ( n3057 & n3058 ) | ( n3057 & ~n3064 ) | ( n3058 & ~n3064 ) ;
  assign n3066 = ( ~n2819 & n3012 ) | ( ~n2819 & n3065 ) | ( n3012 & n3065 ) ;
  assign n3067 = ( n2821 & ~n3012 ) | ( n2821 & n3066 ) | ( ~n3012 & n3066 ) ;
  assign n3068 = ~x17 & n2655 ;
  assign n3069 = ( n369 & ~n2655 ) | ( n369 & n3068 ) | ( ~n2655 & n3068 ) ;
  assign n3070 = x13 & ~n3069 ;
  assign n3071 = n2650 | n2659 ;
  assign n3072 = ( n3069 & n3070 ) | ( n3069 & ~n3071 ) | ( n3070 & ~n3071 ) ;
  assign n3073 = ( x12 & n2641 ) | ( x12 & n3072 ) | ( n2641 & n3072 ) ;
  assign n3074 = ~n2641 & n3073 ;
  assign n3075 = ( x14 & ~x15 ) | ( x14 & n3074 ) | ( ~x15 & n3074 ) ;
  assign n3076 = ~x16 & n1908 ;
  assign n3077 = ~x17 & n3076 ;
  assign n3078 = ( ~x13 & n3030 ) | ( ~x13 & n3077 ) | ( n3030 & n3077 ) ;
  assign n3079 = ( n3032 & ~n3077 ) | ( n3032 & n3078 ) | ( ~n3077 & n3078 ) ;
  assign n3080 = ( x14 & x15 ) | ( x14 & n3079 ) | ( x15 & n3079 ) ;
  assign n3081 = n3075 | n3080 ;
  assign n3082 = ( x11 & ~x14 ) | ( x11 & n3081 ) | ( ~x14 & n3081 ) ;
  assign n3083 = x40 & ~n3082 ;
  assign n3084 = ( x11 & x40 ) | ( x11 & ~n3083 ) | ( x40 & ~n3083 ) ;
  assign n3085 = ( x5 & ~x10 ) | ( x5 & n3084 ) | ( ~x10 & n3084 ) ;
  assign n3086 = ( x10 & ~n1103 ) | ( x10 & n3085 ) | ( ~n1103 & n3085 ) ;
  assign n3087 = ~n3045 & n3086 ;
  assign n3088 = x4 | n3087 ;
  assign n3089 = ~n3024 & n3088 ;
  assign n3090 = ( x2 & ~x3 ) | ( x2 & n3089 ) | ( ~x3 & n3089 ) ;
  assign n3091 = n3053 | n3090 ;
  assign n3092 = ~n3020 & n3091 ;
  assign n3093 = x1 | n3092 ;
  assign n3094 = ~n3016 & n3093 ;
  assign n3095 = ( x0 & x36 ) | ( x0 & ~n3094 ) | ( x36 & ~n3094 ) ;
  assign n3096 = ( ~n3064 & n3094 ) | ( ~n3064 & n3095 ) | ( n3094 & n3095 ) ;
  assign n3097 = ( ~n2819 & n3012 ) | ( ~n2819 & n3096 ) | ( n3012 & n3096 ) ;
  assign n3098 = ( n2821 & ~n3012 ) | ( n2821 & n3097 ) | ( ~n3012 & n3097 ) ;
  assign n3099 = ~x15 & x18 ;
  assign n3100 = ~x19 & n693 ;
  assign n3101 = ( x15 & x19 ) | ( x15 & n3100 ) | ( x19 & n3100 ) ;
  assign n3102 = ( x15 & ~x18 ) | ( x15 & n3101 ) | ( ~x18 & n3101 ) ;
  assign n3103 = ( n3099 & ~n3101 ) | ( n3099 & n3102 ) | ( ~n3101 & n3102 ) ;
  assign n3104 = ( x36 & ~n396 ) | ( x36 & n3103 ) | ( ~n396 & n3103 ) ;
  assign n3105 = n3103 & ~n3104 ;
  assign n3106 = ~x14 & n3105 ;
  assign n3107 = ( x13 & ~x16 ) | ( x13 & n3106 ) | ( ~x16 & n3106 ) ;
  assign n3108 = ~x13 & n3107 ;
  assign n3109 = ( x10 & n198 ) | ( x10 & n3108 ) | ( n198 & n3108 ) ;
  assign n3110 = ~x10 & n3109 ;
  assign n3111 = ~x8 & n3110 ;
  assign n3112 = ( x5 & ~x9 ) | ( x5 & n3111 ) | ( ~x9 & n3111 ) ;
  assign n3113 = ~x5 & n3112 ;
  assign n3114 = ~x3 & n3113 ;
  assign n3115 = ( x2 & ~x4 ) | ( x2 & n3114 ) | ( ~x4 & n3114 ) ;
  assign n3116 = ~x2 & n3115 ;
  assign n3117 = ~x0 & n3116 ;
  assign n3118 = ~x1 & n3117 ;
  assign n3119 = ~x3 & n927 ;
  assign n3120 = ( x0 & x2 ) | ( x0 & n3119 ) | ( x2 & n3119 ) ;
  assign n3121 = ~x0 & n3120 ;
  assign n3122 = x26 & ~n212 ;
  assign n3123 = ( x15 & x26 ) | ( x15 & ~n3122 ) | ( x26 & ~n3122 ) ;
  assign n3124 = ( x28 & n58 ) | ( x28 & ~n3123 ) | ( n58 & ~n3123 ) ;
  assign n3125 = n3123 & n3124 ;
  assign n3126 = ~x0 & x3 ;
  assign n3127 = x3 & ~n3126 ;
  assign n3128 = n165 & n3127 ;
  assign n3129 = ( x18 & x19 ) | ( x18 & ~x40 ) | ( x19 & ~x40 ) ;
  assign n3130 = n2082 & ~n3129 ;
  assign n3131 = ~x15 & n3130 ;
  assign n3132 = ( ~n3126 & n3127 ) | ( ~n3126 & n3131 ) | ( n3127 & n3131 ) ;
  assign n3133 = ( ~x0 & n3128 ) | ( ~x0 & n3132 ) | ( n3128 & n3132 ) ;
  assign n3134 = ( x12 & ~x16 ) | ( x12 & n3133 ) | ( ~x16 & n3133 ) ;
  assign n3135 = x3 & ~x19 ;
  assign n3136 = x18 & ~x40 ;
  assign n3137 = ( ~x18 & x19 ) | ( ~x18 & n3136 ) | ( x19 & n3136 ) ;
  assign n3138 = ( ~x3 & x19 ) | ( ~x3 & n3137 ) | ( x19 & n3137 ) ;
  assign n3139 = ( n3135 & ~n3137 ) | ( n3135 & n3138 ) | ( ~n3137 & n3138 ) ;
  assign n3140 = ( x15 & n84 ) | ( x15 & ~n3139 ) | ( n84 & ~n3139 ) ;
  assign n3141 = n3139 & n3140 ;
  assign n3142 = ~x0 & n3141 ;
  assign n3143 = ~x12 & n3142 ;
  assign n3144 = ( n3133 & ~n3134 ) | ( n3133 & n3143 ) | ( ~n3134 & n3143 ) ;
  assign n3145 = ( x0 & x3 ) | ( x0 & ~n3144 ) | ( x3 & ~n3144 ) ;
  assign n3146 = n3125 & n3145 ;
  assign n3147 = ( n3125 & n3144 ) | ( n3125 & ~n3146 ) | ( n3144 & ~n3146 ) ;
  assign n3148 = x13 & n3147 ;
  assign n3149 = ~x23 & n1818 ;
  assign n3150 = ( x20 & n624 ) | ( x20 & n3149 ) | ( n624 & n3149 ) ;
  assign n3151 = ~x20 & n3150 ;
  assign n3152 = ( x15 & x16 ) | ( x15 & n952 ) | ( x16 & n952 ) ;
  assign n3153 = ~n525 & n3152 ;
  assign n3154 = ~x3 & n3153 ;
  assign n3155 = x3 & ~x16 ;
  assign n3156 = ( x15 & n878 ) | ( x15 & n3155 ) | ( n878 & n3155 ) ;
  assign n3157 = ~x15 & n3156 ;
  assign n3158 = n3154 | n3157 ;
  assign n3159 = ( n3151 & n3154 ) | ( n3151 & n3158 ) | ( n3154 & n3158 ) ;
  assign n3160 = ( x12 & n2869 ) | ( x12 & ~n3159 ) | ( n2869 & ~n3159 ) ;
  assign n3161 = n3159 & n3160 ;
  assign n3162 = n3148 | n3161 ;
  assign n3163 = ( ~x0 & n3148 ) | ( ~x0 & n3162 ) | ( n3148 & n3162 ) ;
  assign n3164 = ~x5 & n3163 ;
  assign n3165 = ( x23 & ~x24 ) | ( x23 & x27 ) | ( ~x24 & x27 ) ;
  assign n3166 = ( ~x24 & x26 ) | ( ~x24 & n3165 ) | ( x26 & n3165 ) ;
  assign n3167 = n3165 & n3166 ;
  assign n3168 = n624 | n3167 ;
  assign n3169 = ( n1053 & n1054 ) | ( n1053 & n3168 ) | ( n1054 & n3168 ) ;
  assign n3170 = ( n972 & ~n1357 ) | ( n972 & n3169 ) | ( ~n1357 & n3169 ) ;
  assign n3171 = ( x21 & n1703 ) | ( x21 & ~n3170 ) | ( n1703 & ~n3170 ) ;
  assign n3172 = ( x18 & n1481 ) | ( x18 & ~n3171 ) | ( n1481 & ~n3171 ) ;
  assign n3173 = n3171 & n3172 ;
  assign n3174 = ~x15 & n3173 ;
  assign n3175 = ( x13 & ~x16 ) | ( x13 & n3174 ) | ( ~x16 & n3174 ) ;
  assign n3176 = ~x13 & n3175 ;
  assign n3177 = x3 & x12 ;
  assign n3178 = ( x5 & ~n3176 ) | ( x5 & n3177 ) | ( ~n3176 & n3177 ) ;
  assign n3179 = n3176 & n3178 ;
  assign n3180 = n3164 | n3179 ;
  assign n3181 = ( ~x0 & n3164 ) | ( ~x0 & n3180 ) | ( n3164 & n3180 ) ;
  assign n3182 = ( x2 & x14 ) | ( x2 & n3181 ) | ( x14 & n3181 ) ;
  assign n3183 = x14 & x16 ;
  assign n3184 = ( x15 & ~n396 ) | ( x15 & n3183 ) | ( ~n396 & n3183 ) ;
  assign n3185 = n396 & n3184 ;
  assign n3186 = x13 & n3185 ;
  assign n3187 = ( x5 & x12 ) | ( x5 & n3186 ) | ( x12 & n3186 ) ;
  assign n3188 = ~x5 & n3187 ;
  assign n3189 = ~x0 & n3188 ;
  assign n3190 = ~x3 & n3189 ;
  assign n3191 = ~x2 & n3190 ;
  assign n3192 = ( n3181 & ~n3182 ) | ( n3181 & n3191 ) | ( ~n3182 & n3191 ) ;
  assign n3193 = ~x20 & n1481 ;
  assign n3194 = n1820 & n3193 ;
  assign n3195 = ( x3 & x15 ) | ( x3 & n3194 ) | ( x15 & n3194 ) ;
  assign n3196 = ~x15 & n3195 ;
  assign n3197 = ( ~x3 & n51 ) | ( ~x3 & n3196 ) | ( n51 & n3196 ) ;
  assign n3198 = x15 & ~n3197 ;
  assign n3199 = ( x15 & n3196 ) | ( x15 & ~n3198 ) | ( n3196 & ~n3198 ) ;
  assign n3200 = ~x14 & x18 ;
  assign n3201 = ( x16 & n3199 ) | ( x16 & ~n3200 ) | ( n3199 & ~n3200 ) ;
  assign n3202 = n3199 & ~n3201 ;
  assign n3203 = x5 & n3202 ;
  assign n3204 = ( x12 & x13 ) | ( x12 & n3203 ) | ( x13 & n3203 ) ;
  assign n3205 = ~x13 & n3204 ;
  assign n3206 = ~x2 & x4 ;
  assign n3207 = ( x0 & n3205 ) | ( x0 & n3206 ) | ( n3205 & n3206 ) ;
  assign n3208 = ~x0 & n3207 ;
  assign n3209 = ( ~n3121 & n3192 ) | ( ~n3121 & n3208 ) | ( n3192 & n3208 ) ;
  assign n3210 = x4 & ~n3208 ;
  assign n3211 = ( n3121 & n3209 ) | ( n3121 & ~n3210 ) | ( n3209 & ~n3210 ) ;
  assign n3212 = ( x11 & n391 ) | ( x11 & n3211 ) | ( n391 & n3211 ) ;
  assign n3213 = n3211 & ~n3212 ;
  assign n3214 = ~x8 & n3213 ;
  assign n3215 = ( x1 & ~x9 ) | ( x1 & n3214 ) | ( ~x9 & n3214 ) ;
  assign n3216 = ~x1 & n3215 ;
  assign n3217 = x5 & n250 ;
  assign n3218 = ( x4 & ~n1996 ) | ( x4 & n3217 ) | ( ~n1996 & n3217 ) ;
  assign n3219 = n1996 & n3218 ;
  assign n3220 = ( x36 & n1821 ) | ( x36 & ~n3219 ) | ( n1821 & ~n3219 ) ;
  assign n3221 = ( x13 & x15 ) | ( x13 & n239 ) | ( x15 & n239 ) ;
  assign n3222 = ~x13 & n3221 ;
  assign n3223 = x33 & x40 ;
  assign n3224 = ( ~x32 & x34 ) | ( ~x32 & n3223 ) | ( x34 & n3223 ) ;
  assign n3225 = x32 & n3224 ;
  assign n3226 = x30 & n3225 ;
  assign n3227 = ( x5 & x13 ) | ( x5 & n3226 ) | ( x13 & n3226 ) ;
  assign n3228 = ~x5 & n3227 ;
  assign n3229 = x15 & n487 ;
  assign n3230 = ( ~x19 & n123 ) | ( ~x19 & n3229 ) | ( n123 & n3229 ) ;
  assign n3231 = ~x3 & x27 ;
  assign n3232 = ( ~x5 & n561 ) | ( ~x5 & n3231 ) | ( n561 & n3231 ) ;
  assign n3233 = ~n561 & n3232 ;
  assign n3234 = ( ~x2 & x24 ) | ( ~x2 & n3233 ) | ( x24 & n3233 ) ;
  assign n3235 = x22 & ~x27 ;
  assign n3236 = ( x23 & n2541 ) | ( x23 & n3235 ) | ( n2541 & n3235 ) ;
  assign n3237 = ~x23 & n3236 ;
  assign n3238 = ~x24 & n3237 ;
  assign n3239 = ( n3233 & ~n3234 ) | ( n3233 & n3238 ) | ( ~n3234 & n3238 ) ;
  assign n3240 = x27 & n2541 ;
  assign n3241 = ( x24 & ~n1829 ) | ( x24 & n3240 ) | ( ~n1829 & n3240 ) ;
  assign n3242 = n1829 & n3241 ;
  assign n3243 = ~n3239 & n3242 ;
  assign n3244 = ( n562 & n3239 ) | ( n562 & n3243 ) | ( n3239 & n3243 ) ;
  assign n3245 = x2 & x5 ;
  assign n3246 = ( x3 & n1735 ) | ( x3 & n3245 ) | ( n1735 & n3245 ) ;
  assign n3247 = ~x3 & n3246 ;
  assign n3248 = ~x15 & n3247 ;
  assign n3249 = ( ~x15 & n3244 ) | ( ~x15 & n3248 ) | ( n3244 & n3248 ) ;
  assign n3250 = ~x19 & n3249 ;
  assign n3251 = ( ~n123 & n3230 ) | ( ~n123 & n3250 ) | ( n3230 & n3250 ) ;
  assign n3252 = ( x17 & x18 ) | ( x17 & ~n3251 ) | ( x18 & ~n3251 ) ;
  assign n3253 = n1416 & ~n2477 ;
  assign n3254 = ( x15 & x18 ) | ( x15 & n3253 ) | ( x18 & n3253 ) ;
  assign n3255 = ~x18 & n3254 ;
  assign n3256 = x17 & n3255 ;
  assign n3257 = ( n3251 & n3252 ) | ( n3251 & n3256 ) | ( n3252 & n3256 ) ;
  assign n3258 = ~n123 & n169 ;
  assign n3259 = ( n416 & n3257 ) | ( n416 & n3258 ) | ( n3257 & n3258 ) ;
  assign n3260 = n1310 & ~n3259 ;
  assign n3261 = ( n1310 & n3257 ) | ( n1310 & ~n3260 ) | ( n3257 & ~n3260 ) ;
  assign n3262 = ( x13 & x16 ) | ( x13 & n3261 ) | ( x16 & n3261 ) ;
  assign n3263 = n71 & ~n123 ;
  assign n3264 = ( n83 & n1417 ) | ( n83 & ~n3263 ) | ( n1417 & ~n3263 ) ;
  assign n3265 = n1417 & ~n3264 ;
  assign n3266 = ~x13 & n3265 ;
  assign n3267 = ( n3261 & ~n3262 ) | ( n3261 & n3266 ) | ( ~n3262 & n3266 ) ;
  assign n3268 = ( x2 & x3 ) | ( x2 & ~n3267 ) | ( x3 & ~n3267 ) ;
  assign n3269 = n3228 & n3268 ;
  assign n3270 = ( n3228 & n3267 ) | ( n3228 & ~n3269 ) | ( n3267 & ~n3269 ) ;
  assign n3271 = ~x14 & n3270 ;
  assign n3272 = n2477 & ~n3271 ;
  assign n3273 = ( n3222 & n3271 ) | ( n3222 & ~n3272 ) | ( n3271 & ~n3272 ) ;
  assign n3274 = ( x4 & ~x12 ) | ( x4 & n3273 ) | ( ~x12 & n3273 ) ;
  assign n3275 = x40 & n1161 ;
  assign n3276 = x15 & n3275 ;
  assign n3277 = ~n1867 & n3276 ;
  assign n3278 = ~n123 & n3277 ;
  assign n3279 = ~x4 & n3278 ;
  assign n3280 = ( n3273 & ~n3274 ) | ( n3273 & n3279 ) | ( ~n3274 & n3279 ) ;
  assign n3281 = ~x36 & n3280 ;
  assign n3282 = ( n1821 & ~n3220 ) | ( n1821 & n3281 ) | ( ~n3220 & n3281 ) ;
  assign n3283 = ~x10 & n3282 ;
  assign n3284 = ( x9 & ~x11 ) | ( x9 & n3283 ) | ( ~x11 & n3283 ) ;
  assign n3285 = ~x9 & n3284 ;
  assign n3286 = ~x1 & n3285 ;
  assign n3287 = ( x0 & ~x8 ) | ( x0 & n3286 ) | ( ~x8 & n3286 ) ;
  assign n3288 = ~x0 & n3287 ;
  assign n3289 = x13 | x14 ;
  assign n3290 = x12 & ~n3289 ;
  assign n3291 = ( x3 & ~n156 ) | ( x3 & n3290 ) | ( ~n156 & n3290 ) ;
  assign n3292 = n156 & n3291 ;
  assign n3293 = x14 & ~n2549 ;
  assign n3294 = ( x16 & ~n66 ) | ( x16 & n71 ) | ( ~n66 & n71 ) ;
  assign n3295 = x13 & ~n3294 ;
  assign n3296 = x14 | n3295 ;
  assign n3297 = ~n3293 & n3296 ;
  assign n3298 = ( x12 & ~x15 ) | ( x12 & n3297 ) | ( ~x15 & n3297 ) ;
  assign n3299 = ( x14 & ~n952 ) | ( x14 & n1140 ) | ( ~n952 & n1140 ) ;
  assign n3300 = n952 & n3299 ;
  assign n3301 = ( x13 & n231 ) | ( x13 & ~n689 ) | ( n231 & ~n689 ) ;
  assign n3302 = ~x13 & n3301 ;
  assign n3303 = ~x14 & x20 ;
  assign n3304 = x13 & n3303 ;
  assign n3305 = x29 & n3304 ;
  assign n3306 = ( x23 & ~n1818 ) | ( x23 & n3305 ) | ( ~n1818 & n3305 ) ;
  assign n3307 = n1818 & n3306 ;
  assign n3308 = ( x14 & ~n1165 ) | ( x14 & n3307 ) | ( ~n1165 & n3307 ) ;
  assign n3309 = x13 & ~n3307 ;
  assign n3310 = ( n1165 & n3308 ) | ( n1165 & ~n3309 ) | ( n3308 & ~n3309 ) ;
  assign n3311 = ( ~n3300 & n3302 ) | ( ~n3300 & n3310 ) | ( n3302 & n3310 ) ;
  assign n3312 = x17 | n3310 ;
  assign n3313 = ( n3300 & n3311 ) | ( n3300 & n3312 ) | ( n3311 & n3312 ) ;
  assign n3314 = ( x12 & x15 ) | ( x12 & ~n3313 ) | ( x15 & ~n3313 ) ;
  assign n3315 = n3298 & ~n3314 ;
  assign n3316 = ( n153 & n160 ) | ( n153 & n3315 ) | ( n160 & n3315 ) ;
  assign n3317 = n304 & ~n3316 ;
  assign n3318 = ( n304 & n3315 ) | ( n304 & ~n3317 ) | ( n3315 & ~n3317 ) ;
  assign n3319 = ( ~x3 & n3292 ) | ( ~x3 & n3318 ) | ( n3292 & n3318 ) ;
  assign n3320 = x40 & ~n3319 ;
  assign n3321 = ( x40 & n3292 ) | ( x40 & ~n3320 ) | ( n3292 & ~n3320 ) ;
  assign n3322 = ( ~x0 & x5 ) | ( ~x0 & n3321 ) | ( x5 & n3321 ) ;
  assign n3323 = ~x3 & n239 ;
  assign n3324 = ~x12 & n3323 ;
  assign n3325 = ( x24 & x26 ) | ( x24 & ~x27 ) | ( x26 & ~x27 ) ;
  assign n3326 = ( x24 & x25 ) | ( x24 & x27 ) | ( x25 & x27 ) ;
  assign n3327 = n3325 & n3326 ;
  assign n3328 = x23 & n3327 ;
  assign n3329 = x22 & n3328 ;
  assign n3330 = ( x20 & x21 ) | ( x20 & n3329 ) | ( x21 & n3329 ) ;
  assign n3331 = ~x20 & n3330 ;
  assign n3332 = x3 & n3331 ;
  assign n3333 = ( x12 & x14 ) | ( x12 & n3332 ) | ( x14 & n3332 ) ;
  assign n3334 = ~x14 & n3333 ;
  assign n3335 = ( x3 & n1416 ) | ( x3 & n1521 ) | ( n1416 & n1521 ) ;
  assign n3336 = ~x3 & n3335 ;
  assign n3337 = ( ~n3324 & n3334 ) | ( ~n3324 & n3336 ) | ( n3334 & n3336 ) ;
  assign n3338 = x19 & ~n3336 ;
  assign n3339 = ( n3324 & n3337 ) | ( n3324 & ~n3338 ) | ( n3337 & ~n3338 ) ;
  assign n3340 = x15 | n3339 ;
  assign n3341 = ~x3 & n2692 ;
  assign n3342 = x15 & ~n3341 ;
  assign n3343 = n3340 & ~n3342 ;
  assign n3344 = x16 | n3343 ;
  assign n3345 = ~x3 & n2696 ;
  assign n3346 = x16 & ~n3345 ;
  assign n3347 = n3344 & ~n3346 ;
  assign n3348 = x18 & ~n3347 ;
  assign n3349 = ~x3 & n2679 ;
  assign n3350 = x18 | n3349 ;
  assign n3351 = ~n3348 & n3350 ;
  assign n3352 = ( x13 & ~x17 ) | ( x13 & n3351 ) | ( ~x17 & n3351 ) ;
  assign n3353 = ( x17 & ~n345 ) | ( x17 & n1524 ) | ( ~n345 & n1524 ) ;
  assign n3354 = n1524 & ~n3353 ;
  assign n3355 = ~x13 & n3354 ;
  assign n3356 = ( n3351 & ~n3352 ) | ( n3351 & n3355 ) | ( ~n3352 & n3355 ) ;
  assign n3357 = ( x14 & ~n1940 ) | ( x14 & n2368 ) | ( ~n1940 & n2368 ) ;
  assign n3358 = n1940 & n3357 ;
  assign n3359 = ( ~x3 & n3356 ) | ( ~x3 & n3358 ) | ( n3356 & n3358 ) ;
  assign n3360 = x12 & ~n3359 ;
  assign n3361 = ( x12 & n3356 ) | ( x12 & ~n3360 ) | ( n3356 & ~n3360 ) ;
  assign n3362 = ( x0 & x5 ) | ( x0 & ~n3361 ) | ( x5 & ~n3361 ) ;
  assign n3363 = n3322 & ~n3362 ;
  assign n3364 = ~x3 & n154 ;
  assign n3365 = x0 & n3364 ;
  assign n3366 = n77 & n3365 ;
  assign n3367 = ( x14 & ~n76 ) | ( x14 & n3366 ) | ( ~n76 & n3366 ) ;
  assign n3368 = ~x14 & n3367 ;
  assign n3369 = ~n3363 & n3368 ;
  assign n3370 = ( ~n848 & n3363 ) | ( ~n848 & n3369 ) | ( n3363 & n3369 ) ;
  assign n3371 = ~x9 & n3370 ;
  assign n3372 = ( x8 & ~x10 ) | ( x8 & n3371 ) | ( ~x10 & n3371 ) ;
  assign n3373 = ~x8 & n3372 ;
  assign n3374 = ~x2 & n3373 ;
  assign n3375 = ( x1 & ~x4 ) | ( x1 & n3374 ) | ( ~x4 & n3374 ) ;
  assign n3376 = ~x1 & n3375 ;
  assign n3377 = ~x5 & n564 ;
  assign n3378 = x20 | n3377 ;
  assign n3379 = ( ~x21 & n3377 ) | ( ~x21 & n3378 ) | ( n3377 & n3378 ) ;
  assign n3380 = x27 & n3379 ;
  assign n3381 = ~x3 & n3380 ;
  assign n3382 = ~x4 & n3381 ;
  assign n3383 = x2 & n3382 ;
  assign n3384 = x3 & n631 ;
  assign n3385 = x23 & x26 ;
  assign n3386 = ( ~x22 & x24 ) | ( ~x22 & n3385 ) | ( x24 & n3385 ) ;
  assign n3387 = x22 & n3386 ;
  assign n3388 = x27 & n3387 ;
  assign n3389 = x24 | n561 ;
  assign n3390 = ~x27 & n3389 ;
  assign n3391 = n3388 | n3390 ;
  assign n3392 = ( x3 & ~n631 ) | ( x3 & n3391 ) | ( ~n631 & n3391 ) ;
  assign n3393 = x3 | x40 ;
  assign n3394 = ( n3384 & ~n3392 ) | ( n3384 & n3393 ) | ( ~n3392 & n3393 ) ;
  assign n3395 = ~x5 & n3394 ;
  assign n3396 = ~x3 & x23 ;
  assign n3397 = x23 & ~n3396 ;
  assign n3398 = n3327 & n3397 ;
  assign n3399 = ( n1742 & ~n3396 ) | ( n1742 & n3397 ) | ( ~n3396 & n3397 ) ;
  assign n3400 = ( ~x3 & n3398 ) | ( ~x3 & n3399 ) | ( n3398 & n3399 ) ;
  assign n3401 = x22 & ~n3400 ;
  assign n3402 = ~x3 & n1742 ;
  assign n3403 = x22 | n3402 ;
  assign n3404 = ~n3401 & n3403 ;
  assign n3405 = ~x26 & x27 ;
  assign n3406 = ( ~x24 & x27 ) | ( ~x24 & n3405 ) | ( x27 & n3405 ) ;
  assign n3407 = ( x23 & n1705 ) | ( x23 & ~n2518 ) | ( n1705 & ~n2518 ) ;
  assign n3408 = ( ~x23 & n2518 ) | ( ~x23 & n3406 ) | ( n2518 & n3406 ) ;
  assign n3409 = ( ~n3406 & n3407 ) | ( ~n3406 & n3408 ) | ( n3407 & n3408 ) ;
  assign n3410 = ~n3404 & n3409 ;
  assign n3411 = x5 & ~n3410 ;
  assign n3412 = n3395 | n3411 ;
  assign n3413 = x4 | n3412 ;
  assign n3414 = x5 & ~n561 ;
  assign n3415 = x3 & ~n561 ;
  assign n3416 = ( ~x3 & x5 ) | ( ~x3 & n561 ) | ( x5 & n561 ) ;
  assign n3417 = ( ~n3414 & n3415 ) | ( ~n3414 & n3416 ) | ( n3415 & n3416 ) ;
  assign n3418 = ~x24 & n3417 ;
  assign n3419 = ~x22 & n1270 ;
  assign n3420 = x24 & ~n3419 ;
  assign n3421 = n3418 | n3420 ;
  assign n3422 = x27 & ~n3421 ;
  assign n3423 = x4 & ~n3422 ;
  assign n3424 = n3413 & ~n3423 ;
  assign n3425 = ( x20 & ~x21 ) | ( x20 & n3424 ) | ( ~x21 & n3424 ) ;
  assign n3426 = x40 & ~n155 ;
  assign n3427 = ( x5 & x20 ) | ( x5 & n3426 ) | ( x20 & n3426 ) ;
  assign n3428 = ~x5 & n3427 ;
  assign n3429 = x21 & n3428 ;
  assign n3430 = ( n3424 & ~n3425 ) | ( n3424 & n3429 ) | ( ~n3425 & n3429 ) ;
  assign n3431 = ( ~x3 & x4 ) | ( ~x3 & n601 ) | ( x4 & n601 ) ;
  assign n3432 = ( x3 & x4 ) | ( x3 & ~x27 ) | ( x4 & ~x27 ) ;
  assign n3433 = n3431 & ~n3432 ;
  assign n3434 = x3 & ~x27 ;
  assign n3435 = ( x4 & x5 ) | ( x4 & n3434 ) | ( x5 & n3434 ) ;
  assign n3436 = ~x4 & n3435 ;
  assign n3437 = ~n3433 & n3436 ;
  assign n3438 = ( n918 & n3433 ) | ( n918 & n3437 ) | ( n3433 & n3437 ) ;
  assign n3439 = n3430 | n3438 ;
  assign n3440 = ~x2 & n3439 ;
  assign n3441 = n3383 | n3440 ;
  assign n3442 = ( x36 & ~n878 ) | ( x36 & n3441 ) | ( ~n878 & n3441 ) ;
  assign n3443 = n3441 & ~n3442 ;
  assign n3444 = ( x15 & n84 ) | ( x15 & n3443 ) | ( n84 & n3443 ) ;
  assign n3445 = ~x15 & n3444 ;
  assign n3446 = ( x13 & n383 ) | ( x13 & n3445 ) | ( n383 & n3445 ) ;
  assign n3447 = ~x13 & n3446 ;
  assign n3448 = ~x10 & n3447 ;
  assign n3449 = ( x9 & ~x11 ) | ( x9 & n3448 ) | ( ~x11 & n3448 ) ;
  assign n3450 = ~x9 & n3449 ;
  assign n3451 = ~x1 & n3450 ;
  assign n3452 = ( x0 & ~x8 ) | ( x0 & n3451 ) | ( ~x8 & n3451 ) ;
  assign n3453 = ~x0 & n3452 ;
  assign n3454 = n566 | n972 ;
  assign n3455 = ( x16 & x19 ) | ( x16 & x40 ) | ( x19 & x40 ) ;
  assign n3456 = ~n3454 & n3455 ;
  assign n3457 = ( x40 & n3454 ) | ( x40 & n3456 ) | ( n3454 & n3456 ) ;
  assign n3458 = x5 | n3457 ;
  assign n3459 = ~x16 & n568 ;
  assign n3460 = x5 & ~n3459 ;
  assign n3461 = n3458 & ~n3460 ;
  assign n3462 = ( x14 & x15 ) | ( x14 & n3461 ) | ( x15 & n3461 ) ;
  assign n3463 = ~x14 & n3229 ;
  assign n3464 = ( n3461 & ~n3462 ) | ( n3461 & n3463 ) | ( ~n3462 & n3463 ) ;
  assign n3465 = x13 | n3464 ;
  assign n3466 = ~x5 & n239 ;
  assign n3467 = x13 & ~n3466 ;
  assign n3468 = n3465 & ~n3467 ;
  assign n3469 = x18 & ~n3468 ;
  assign n3470 = n135 | n3289 ;
  assign n3471 = ( n135 & ~n2025 ) | ( n135 & n3470 ) | ( ~n2025 & n3470 ) ;
  assign n3472 = n135 & n1161 ;
  assign n3473 = ( n135 & n1115 ) | ( n135 & n3472 ) | ( n1115 & n3472 ) ;
  assign n3474 = x19 & n1161 ;
  assign n3475 = ( x15 & x16 ) | ( x15 & n3474 ) | ( x16 & n3474 ) ;
  assign n3476 = ~x15 & n3475 ;
  assign n3477 = ( x40 & n3473 ) | ( x40 & n3476 ) | ( n3473 & n3476 ) ;
  assign n3478 = n3471 & n3477 ;
  assign n3479 = ( x40 & ~n3471 ) | ( x40 & n3478 ) | ( ~n3471 & n3478 ) ;
  assign n3480 = ~x5 & n3479 ;
  assign n3481 = x18 | n3480 ;
  assign n3482 = ~n3469 & n3481 ;
  assign n3483 = x17 & n3482 ;
  assign n3484 = ( x13 & x14 ) | ( x13 & x40 ) | ( x14 & x40 ) ;
  assign n3485 = ( n134 & ~n322 ) | ( n134 & n878 ) | ( ~n322 & n878 ) ;
  assign n3486 = ( ~x13 & n215 ) | ( ~x13 & n1126 ) | ( n215 & n1126 ) ;
  assign n3487 = ( x17 & ~n3485 ) | ( x17 & n3486 ) | ( ~n3485 & n3486 ) ;
  assign n3488 = ( ~x14 & x18 ) | ( ~x14 & x19 ) | ( x18 & x19 ) ;
  assign n3489 = x19 & ~n3488 ;
  assign n3490 = ( x15 & x18 ) | ( x15 & n3489 ) | ( x18 & n3489 ) ;
  assign n3491 = ( ~n3488 & n3489 ) | ( ~n3488 & n3490 ) | ( n3489 & n3490 ) ;
  assign n3492 = ~x13 & n3491 ;
  assign n3493 = n2143 & ~n3289 ;
  assign n3494 = ( x13 & ~x14 ) | ( x13 & x15 ) | ( ~x14 & x15 ) ;
  assign n3495 = x13 | n3494 ;
  assign n3496 = ( ~x14 & x18 ) | ( ~x14 & n3494 ) | ( x18 & n3494 ) ;
  assign n3497 = x13 & n3496 ;
  assign n3498 = n3495 & ~n3497 ;
  assign n3499 = x15 & n66 ;
  assign n3500 = ~n3289 & n3499 ;
  assign n3501 = x19 & ~n3500 ;
  assign n3502 = ( n3498 & n3500 ) | ( n3498 & ~n3501 ) | ( n3500 & ~n3501 ) ;
  assign n3503 = x16 & ~n3502 ;
  assign n3504 = n66 & n2025 ;
  assign n3505 = x16 | n3504 ;
  assign n3506 = ~n3503 & n3505 ;
  assign n3507 = n3493 | n3506 ;
  assign n3508 = ( n3491 & ~n3492 ) | ( n3491 & n3507 ) | ( ~n3492 & n3507 ) ;
  assign n3509 = ~x17 & n3508 ;
  assign n3510 = ( n3485 & n3487 ) | ( n3485 & ~n3509 ) | ( n3487 & ~n3509 ) ;
  assign n3511 = x40 & ~n3510 ;
  assign n3512 = ( ~x13 & n3484 ) | ( ~x13 & n3511 ) | ( n3484 & n3511 ) ;
  assign n3513 = n3483 | n3512 ;
  assign n3514 = ( ~x5 & n3483 ) | ( ~x5 & n3513 ) | ( n3483 & n3513 ) ;
  assign n3515 = x12 & ~n3514 ;
  assign n3516 = ( x16 & ~n66 ) | ( x16 & n185 ) | ( ~n66 & n185 ) ;
  assign n3517 = n66 | n3516 ;
  assign n3518 = ( x14 & n2452 ) | ( x14 & ~n3517 ) | ( n2452 & ~n3517 ) ;
  assign n3519 = n3517 & n3518 ;
  assign n3520 = ~x5 & n3519 ;
  assign n3521 = x12 | n3520 ;
  assign n3522 = ~n3515 & n3521 ;
  assign n3523 = ( x0 & x3 ) | ( x0 & n3522 ) | ( x3 & n3522 ) ;
  assign n3524 = n156 & n1270 ;
  assign n3525 = n3290 & n3524 ;
  assign n3526 = ~x0 & n3525 ;
  assign n3527 = ( n3522 & ~n3523 ) | ( n3522 & n3526 ) | ( ~n3523 & n3526 ) ;
  assign n3528 = n3368 & ~n3527 ;
  assign n3529 = ( ~n848 & n3527 ) | ( ~n848 & n3528 ) | ( n3527 & n3528 ) ;
  assign n3530 = ~x9 & n3529 ;
  assign n3531 = ( x8 & ~x10 ) | ( x8 & n3530 ) | ( ~x10 & n3530 ) ;
  assign n3532 = ~x8 & n3531 ;
  assign n3533 = ~x2 & n3532 ;
  assign n3534 = ( x1 & ~x4 ) | ( x1 & n3533 ) | ( ~x4 & n3533 ) ;
  assign n3535 = ~x1 & n3534 ;
  assign n3536 = x17 & n2116 ;
  assign n3537 = ( x17 & ~n110 ) | ( x17 & n2116 ) | ( ~n110 & n2116 ) ;
  assign n3538 = ~n3536 & n3537 ;
  assign n3539 = n1017 | n3538 ;
  assign n3540 = ( n239 & n1017 ) | ( n239 & ~n3539 ) | ( n1017 & ~n3539 ) ;
  assign n3541 = x13 & n3540 ;
  assign n3542 = ( x5 & x12 ) | ( x5 & n3541 ) | ( x12 & n3541 ) ;
  assign n3543 = ~x5 & n3542 ;
  assign n3544 = ~x5 & n2679 ;
  assign n3545 = ( x3 & ~x18 ) | ( x3 & n3544 ) | ( ~x18 & n3544 ) ;
  assign n3546 = ~x3 & n3545 ;
  assign n3547 = x12 & ~x19 ;
  assign n3548 = ( x14 & n633 ) | ( x14 & n3547 ) | ( n633 & n3547 ) ;
  assign n3549 = ~x14 & n3548 ;
  assign n3550 = x3 & ~n3549 ;
  assign n3551 = x19 | n972 ;
  assign n3552 = ( x12 & x19 ) | ( x12 & ~n3551 ) | ( x19 & ~n3551 ) ;
  assign n3553 = ( x12 & ~x14 ) | ( x12 & n3552 ) | ( ~x14 & n3552 ) ;
  assign n3554 = ( n1521 & ~n3552 ) | ( n1521 & n3553 ) | ( ~n3552 & n3553 ) ;
  assign n3555 = x40 & n3554 ;
  assign n3556 = x3 | n3555 ;
  assign n3557 = ~n3550 & n3556 ;
  assign n3558 = x5 | n3557 ;
  assign n3559 = ~x14 & n2767 ;
  assign n3560 = x12 & n3559 ;
  assign n3561 = x3 & n3560 ;
  assign n3562 = x5 & ~n3561 ;
  assign n3563 = n3558 & ~n3562 ;
  assign n3564 = x2 | n3563 ;
  assign n3565 = ( x14 & n3380 ) | ( x14 & n3547 ) | ( n3380 & n3547 ) ;
  assign n3566 = ~x14 & n3565 ;
  assign n3567 = ~x3 & n3566 ;
  assign n3568 = x2 & ~n3567 ;
  assign n3569 = n3564 & ~n3568 ;
  assign n3570 = ~x15 & n3569 ;
  assign n3571 = ( x3 & n169 ) | ( x3 & n2692 ) | ( n169 & n2692 ) ;
  assign n3572 = ~x3 & n3571 ;
  assign n3573 = n3570 | n3572 ;
  assign n3574 = ( ~x2 & n3570 ) | ( ~x2 & n3573 ) | ( n3570 & n3573 ) ;
  assign n3575 = ( x16 & ~x18 ) | ( x16 & n3574 ) | ( ~x18 & n3574 ) ;
  assign n3576 = ~x3 & n2697 ;
  assign n3577 = ( x2 & ~x5 ) | ( x2 & n3576 ) | ( ~x5 & n3576 ) ;
  assign n3578 = ~x2 & n3577 ;
  assign n3579 = x18 & n3578 ;
  assign n3580 = ( n3574 & ~n3575 ) | ( n3574 & n3579 ) | ( ~n3575 & n3579 ) ;
  assign n3581 = x2 & ~n3580 ;
  assign n3582 = ( n3546 & n3580 ) | ( n3546 & ~n3581 ) | ( n3580 & ~n3581 ) ;
  assign n3583 = ( x13 & ~x17 ) | ( x13 & n3582 ) | ( ~x17 & n3582 ) ;
  assign n3584 = ~x12 & n2702 ;
  assign n3585 = n745 & n3584 ;
  assign n3586 = n1524 & ~n3585 ;
  assign n3587 = ( n396 & n3585 ) | ( n396 & n3586 ) | ( n3585 & n3586 ) ;
  assign n3588 = ~x3 & n3587 ;
  assign n3589 = ( x2 & ~x5 ) | ( x2 & n3588 ) | ( ~x5 & n3588 ) ;
  assign n3590 = ~x2 & n3589 ;
  assign n3591 = ~x13 & n3590 ;
  assign n3592 = ( n3582 & ~n3583 ) | ( n3582 & n3591 ) | ( ~n3583 & n3591 ) ;
  assign n3593 = ( x2 & x3 ) | ( x2 & ~n3592 ) | ( x3 & ~n3592 ) ;
  assign n3594 = n3543 & n3593 ;
  assign n3595 = ( n3543 & n3592 ) | ( n3543 & ~n3594 ) | ( n3592 & ~n3594 ) ;
  assign n3596 = ( x4 & x36 ) | ( x4 & n3595 ) | ( x36 & n3595 ) ;
  assign n3597 = ( x5 & x24 ) | ( x5 & n561 ) | ( x24 & n561 ) ;
  assign n3598 = ( x5 & n561 ) | ( x5 & ~n3597 ) | ( n561 & ~n3597 ) ;
  assign n3599 = ( n1823 & ~n3597 ) | ( n1823 & n3598 ) | ( ~n3597 & n3598 ) ;
  assign n3600 = ( x21 & n592 ) | ( x21 & ~n3599 ) | ( n592 & ~n3599 ) ;
  assign n3601 = n3599 & n3600 ;
  assign n3602 = x17 & n3601 ;
  assign n3603 = ( x18 & x19 ) | ( x18 & n3602 ) | ( x19 & n3602 ) ;
  assign n3604 = ~x19 & n3603 ;
  assign n3605 = ~x15 & n3604 ;
  assign n3606 = ( x14 & ~x16 ) | ( x14 & n3605 ) | ( ~x16 & n3605 ) ;
  assign n3607 = ~x14 & n3606 ;
  assign n3608 = x4 & n3607 ;
  assign n3609 = ( x12 & x13 ) | ( x12 & n3608 ) | ( x13 & n3608 ) ;
  assign n3610 = ~x13 & n3609 ;
  assign n3611 = n250 & n3610 ;
  assign n3612 = ~x36 & n3611 ;
  assign n3613 = ( n3595 & ~n3596 ) | ( n3595 & n3612 ) | ( ~n3596 & n3612 ) ;
  assign n3614 = ~x10 & n3613 ;
  assign n3615 = ( x9 & ~x11 ) | ( x9 & n3614 ) | ( ~x11 & n3614 ) ;
  assign n3616 = ~x9 & n3615 ;
  assign n3617 = ~x1 & n3616 ;
  assign n3618 = ( x0 & ~x8 ) | ( x0 & n3617 ) | ( ~x8 & n3617 ) ;
  assign n3619 = ~x0 & n3618 ;
  assign n3620 = n94 & ~n796 ;
  assign n3621 = ( n416 & n694 ) | ( n416 & n3620 ) | ( n694 & n3620 ) ;
  assign n3622 = ~n694 & n3621 ;
  assign n3623 = ( ~x15 & x16 ) | ( ~x15 & x17 ) | ( x16 & x17 ) ;
  assign n3624 = ~n524 & n3623 ;
  assign n3625 = ( x16 & x17 ) | ( x16 & ~n3624 ) | ( x17 & ~n3624 ) ;
  assign n3626 = ( x12 & n3622 ) | ( x12 & n3625 ) | ( n3622 & n3625 ) ;
  assign n3627 = x14 & ~n3626 ;
  assign n3628 = ( x14 & n3622 ) | ( x14 & ~n3627 ) | ( n3622 & ~n3627 ) ;
  assign n3629 = x12 & n127 ;
  assign n3630 = n745 & n3629 ;
  assign n3631 = ~n3628 & n3630 ;
  assign n3632 = ( n2368 & n3628 ) | ( n2368 & n3631 ) | ( n3628 & n3631 ) ;
  assign n3633 = ( x2 & ~x12 ) | ( x2 & n3466 ) | ( ~x12 & n3466 ) ;
  assign n3634 = ~x2 & n3633 ;
  assign n3635 = x5 & x20 ;
  assign n3636 = x5 | n1041 ;
  assign n3637 = x21 & n3636 ;
  assign n3638 = ( n562 & n3635 ) | ( n562 & ~n3637 ) | ( n3635 & ~n3637 ) ;
  assign n3639 = ( ~x2 & x27 ) | ( ~x2 & n3638 ) | ( x27 & n3638 ) ;
  assign n3640 = x20 | n3387 ;
  assign n3641 = x21 & ~n3640 ;
  assign n3642 = ( ~x21 & n1323 ) | ( ~x21 & n3641 ) | ( n1323 & n3641 ) ;
  assign n3643 = x40 & n3642 ;
  assign n3644 = ~x5 & n3643 ;
  assign n3645 = ( x2 & x27 ) | ( x2 & n3644 ) | ( x27 & n3644 ) ;
  assign n3646 = n3639 & n3645 ;
  assign n3647 = x21 & x40 ;
  assign n3648 = ~x5 & x20 ;
  assign n3649 = ( x2 & n3647 ) | ( x2 & n3648 ) | ( n3647 & n3648 ) ;
  assign n3650 = ~x2 & n3649 ;
  assign n3651 = ~n3646 & n3650 ;
  assign n3652 = ( n369 & n3646 ) | ( n369 & n3651 ) | ( n3646 & n3651 ) ;
  assign n3653 = x40 & ~n618 ;
  assign n3654 = ~x18 & n3653 ;
  assign n3655 = ~x5 & x16 ;
  assign n3656 = ( x2 & n3654 ) | ( x2 & n3655 ) | ( n3654 & n3655 ) ;
  assign n3657 = ~x2 & n3656 ;
  assign n3658 = ~n3652 & n3657 ;
  assign n3659 = ( n383 & n3652 ) | ( n383 & n3658 ) | ( n3652 & n3658 ) ;
  assign n3660 = ( x12 & x16 ) | ( x12 & n2677 ) | ( x16 & n2677 ) ;
  assign n3661 = ( ~n2676 & n2677 ) | ( ~n2676 & n3660 ) | ( n2677 & n3660 ) ;
  assign n3662 = ( x2 & n169 ) | ( x2 & n3661 ) | ( n169 & n3661 ) ;
  assign n3663 = ~x2 & n3662 ;
  assign n3664 = ( ~n3634 & n3659 ) | ( ~n3634 & n3663 ) | ( n3659 & n3663 ) ;
  assign n3665 = x15 & ~n3663 ;
  assign n3666 = ( n3634 & n3664 ) | ( n3634 & ~n3665 ) | ( n3664 & ~n3665 ) ;
  assign n3667 = ~x19 & n3666 ;
  assign n3668 = n546 | n635 ;
  assign n3669 = ( ~x14 & n796 ) | ( ~x14 & n1521 ) | ( n796 & n1521 ) ;
  assign n3670 = ( n1521 & n3668 ) | ( n1521 & n3669 ) | ( n3668 & n3669 ) ;
  assign n3671 = ( x19 & n487 ) | ( x19 & ~n3670 ) | ( n487 & ~n3670 ) ;
  assign n3672 = n3670 & n3671 ;
  assign n3673 = n3667 | n3672 ;
  assign n3674 = ( ~x2 & n3667 ) | ( ~x2 & n3673 ) | ( n3667 & n3673 ) ;
  assign n3675 = ( x13 & ~x17 ) | ( x13 & n3674 ) | ( ~x17 & n3674 ) ;
  assign n3676 = ( x14 & x15 ) | ( x14 & n1493 ) | ( x15 & n1493 ) ;
  assign n3677 = ~x14 & n3676 ;
  assign n3678 = ~x37 & n3677 ;
  assign n3679 = ( x19 & ~n693 ) | ( x19 & n3678 ) | ( ~n693 & n3678 ) ;
  assign n3680 = ~x19 & n3679 ;
  assign n3681 = ( ~x15 & n1521 ) | ( ~x15 & n3680 ) | ( n1521 & n3680 ) ;
  assign n3682 = n66 & ~n3681 ;
  assign n3683 = ( n66 & n3680 ) | ( n66 & ~n3682 ) | ( n3680 & ~n3682 ) ;
  assign n3684 = ( x16 & ~x40 ) | ( x16 & n3683 ) | ( ~x40 & n3683 ) ;
  assign n3685 = x40 & n1524 ;
  assign n3686 = ( n3683 & ~n3684 ) | ( n3683 & n3685 ) | ( ~n3684 & n3685 ) ;
  assign n3687 = ~x5 & n3686 ;
  assign n3688 = ( x2 & ~x17 ) | ( x2 & n3687 ) | ( ~x17 & n3687 ) ;
  assign n3689 = ~x2 & n3688 ;
  assign n3690 = ~x13 & n3689 ;
  assign n3691 = ( n3674 & ~n3675 ) | ( n3674 & n3690 ) | ( ~n3675 & n3690 ) ;
  assign n3692 = ( x2 & x5 ) | ( x2 & ~n3691 ) | ( x5 & ~n3691 ) ;
  assign n3693 = n3632 & n3692 ;
  assign n3694 = ( n3632 & n3691 ) | ( n3632 & ~n3693 ) | ( n3691 & ~n3693 ) ;
  assign n3695 = ~x4 & n3694 ;
  assign n3696 = n858 | n3695 ;
  assign n3697 = ( ~x2 & n3695 ) | ( ~x2 & n3696 ) | ( n3695 & n3696 ) ;
  assign n3698 = x3 | n3697 ;
  assign n3699 = x24 & n3385 ;
  assign n3700 = x22 & n3699 ;
  assign n3701 = ( x4 & x5 ) | ( x4 & n3700 ) | ( x5 & n3700 ) ;
  assign n3702 = ~x4 & n3701 ;
  assign n3703 = ( ~x5 & n1044 ) | ( ~x5 & n3702 ) | ( n1044 & n3702 ) ;
  assign n3704 = x4 & ~n3703 ;
  assign n3705 = ( x4 & n3702 ) | ( x4 & ~n3704 ) | ( n3702 & ~n3704 ) ;
  assign n3706 = ( x21 & x27 ) | ( x21 & ~n3705 ) | ( x27 & ~n3705 ) ;
  assign n3707 = x23 & x24 ;
  assign n3708 = ( x25 & x27 ) | ( x25 & n3707 ) | ( x27 & n3707 ) ;
  assign n3709 = ~x27 & n3708 ;
  assign n3710 = x22 & n3709 ;
  assign n3711 = ( x4 & x5 ) | ( x4 & n3710 ) | ( x5 & n3710 ) ;
  assign n3712 = ~x4 & n3711 ;
  assign n3713 = x21 & n3712 ;
  assign n3714 = ( n3705 & n3706 ) | ( n3705 & n3713 ) | ( n3706 & n3713 ) ;
  assign n3715 = ( x19 & n1691 ) | ( x19 & n3714 ) | ( n1691 & n3714 ) ;
  assign n3716 = ~x19 & n3715 ;
  assign n3717 = ( x15 & n84 ) | ( x15 & n3716 ) | ( n84 & n3716 ) ;
  assign n3718 = ~x15 & n3717 ;
  assign n3719 = ( x13 & n383 ) | ( x13 & n3718 ) | ( n383 & n3718 ) ;
  assign n3720 = ~x13 & n3719 ;
  assign n3721 = ~x2 & n3720 ;
  assign n3722 = x3 & ~n3721 ;
  assign n3723 = n3698 & ~n3722 ;
  assign n3724 = x1 | x36 ;
  assign n3725 = ( x9 & n3723 ) | ( x9 & n3724 ) | ( n3723 & n3724 ) ;
  assign n3726 = n3723 & ~n3725 ;
  assign n3727 = ( x0 & ~x9 ) | ( x0 & x11 ) | ( ~x9 & x11 ) ;
  assign n3728 = n3726 & n3727 ;
  assign n3729 = ( x9 & n3726 ) | ( x9 & ~n3728 ) | ( n3726 & ~n3728 ) ;
  assign n3730 = ( x8 & x10 ) | ( x8 & n3729 ) | ( x10 & n3729 ) ;
  assign n3731 = ( n1184 & n3729 ) | ( n1184 & ~n3730 ) | ( n3729 & ~n3730 ) ;
  assign n3732 = ( x13 & ~x14 ) | ( x13 & x18 ) | ( ~x14 & x18 ) ;
  assign n3733 = ~x14 & n3732 ;
  assign n3734 = ( x13 & ~x17 ) | ( x13 & n3732 ) | ( ~x17 & n3732 ) ;
  assign n3735 = x14 & ~n3734 ;
  assign n3736 = n3733 | n3735 ;
  assign n3737 = ( x12 & x15 ) | ( x12 & n3736 ) | ( x15 & n3736 ) ;
  assign n3738 = ( x12 & ~n95 ) | ( x12 & n190 ) | ( ~n95 & n190 ) ;
  assign n3739 = ~x12 & n3738 ;
  assign n3740 = x15 & n3739 ;
  assign n3741 = ( ~n3736 & n3737 ) | ( ~n3736 & n3740 ) | ( n3737 & n3740 ) ;
  assign n3742 = ( ~x13 & x14 ) | ( ~x13 & x18 ) | ( x14 & x18 ) ;
  assign n3743 = ( x12 & ~x14 ) | ( x12 & n3742 ) | ( ~x14 & n3742 ) ;
  assign n3744 = ( x13 & x14 ) | ( x13 & n3743 ) | ( x14 & n3743 ) ;
  assign n3745 = n3742 & ~n3744 ;
  assign n3746 = ( x12 & ~n3743 ) | ( x12 & n3745 ) | ( ~n3743 & n3745 ) ;
  assign n3747 = ( x12 & n190 ) | ( x12 & n416 ) | ( n190 & n416 ) ;
  assign n3748 = ~x12 & n3747 ;
  assign n3749 = x17 | n3748 ;
  assign n3750 = ( n3746 & n3748 ) | ( n3746 & n3749 ) | ( n3748 & n3749 ) ;
  assign n3751 = x18 & ~n84 ;
  assign n3752 = ( n878 & n2890 ) | ( n878 & ~n3751 ) | ( n2890 & ~n3751 ) ;
  assign n3753 = ( ~x18 & x19 ) | ( ~x18 & n524 ) | ( x19 & n524 ) ;
  assign n3754 = ( x15 & x16 ) | ( x15 & n3753 ) | ( x16 & n3753 ) ;
  assign n3755 = n524 & ~n3754 ;
  assign n3756 = ( n3753 & ~n3754 ) | ( n3753 & n3755 ) | ( ~n3754 & n3755 ) ;
  assign n3757 = n110 & n477 ;
  assign n3758 = x17 & ~n3757 ;
  assign n3759 = ( n3756 & n3757 ) | ( n3756 & ~n3758 ) | ( n3757 & ~n3758 ) ;
  assign n3760 = x13 & ~n3759 ;
  assign n3761 = ~n3752 & n3760 ;
  assign n3762 = x14 & n3761 ;
  assign n3763 = ( ~x18 & n42 ) | ( ~x18 & n416 ) | ( n42 & n416 ) ;
  assign n3764 = x15 & ~n3763 ;
  assign n3765 = ( x18 & ~n70 ) | ( x18 & n618 ) | ( ~n70 & n618 ) ;
  assign n3766 = x17 & ~n3765 ;
  assign n3767 = x15 | n3766 ;
  assign n3768 = ~n3764 & n3767 ;
  assign n3769 = x16 & ~n3768 ;
  assign n3770 = x15 & n1674 ;
  assign n3771 = x16 | n3770 ;
  assign n3772 = ~n3769 & n3771 ;
  assign n3773 = ~x13 & n3772 ;
  assign n3774 = x14 | n3773 ;
  assign n3775 = ~n3762 & n3774 ;
  assign n3776 = x12 & ~n3775 ;
  assign n3777 = ( x16 & ~x17 ) | ( x16 & n45 ) | ( ~x17 & n45 ) ;
  assign n3778 = ( x18 & ~x19 ) | ( x18 & n3777 ) | ( ~x19 & n3777 ) ;
  assign n3779 = ~n45 & n3778 ;
  assign n3780 = ( ~n3777 & n3778 ) | ( ~n3777 & n3779 ) | ( n3778 & n3779 ) ;
  assign n3781 = ( ~x14 & x15 ) | ( ~x14 & n3780 ) | ( x15 & n3780 ) ;
  assign n3782 = x18 & ~n94 ;
  assign n3783 = ( n878 & n2890 ) | ( n878 & ~n3782 ) | ( n2890 & ~n3782 ) ;
  assign n3784 = x14 & n3783 ;
  assign n3785 = ( n3780 & ~n3781 ) | ( n3780 & n3784 ) | ( ~n3781 & n3784 ) ;
  assign n3786 = ~x13 & n3785 ;
  assign n3787 = x12 | n3786 ;
  assign n3788 = ~n3776 & n3787 ;
  assign n3789 = ( ~n3741 & n3750 ) | ( ~n3741 & n3788 ) | ( n3750 & n3788 ) ;
  assign n3790 = n135 | n3788 ;
  assign n3791 = ( n3741 & n3789 ) | ( n3741 & n3790 ) | ( n3789 & n3790 ) ;
  assign n3792 = ( x13 & x14 ) | ( x13 & x17 ) | ( x14 & x17 ) ;
  assign n3793 = ( ~x15 & x17 ) | ( ~x15 & n3792 ) | ( x17 & n3792 ) ;
  assign n3794 = x17 & ~n3793 ;
  assign n3795 = n3793 | n3794 ;
  assign n3796 = ( ~x17 & n3794 ) | ( ~x17 & n3795 ) | ( n3794 & n3795 ) ;
  assign n3797 = ~x12 & n3796 ;
  assign n3798 = ( x12 & n190 ) | ( x12 & n570 ) | ( n190 & n570 ) ;
  assign n3799 = ~x12 & n3798 ;
  assign n3800 = ( ~x12 & x13 ) | ( ~x12 & x14 ) | ( x13 & x14 ) ;
  assign n3801 = ( x14 & x15 ) | ( x14 & ~n3800 ) | ( x15 & ~n3800 ) ;
  assign n3802 = ( x12 & ~x13 ) | ( x12 & n3801 ) | ( ~x13 & n3801 ) ;
  assign n3803 = n3800 & n3802 ;
  assign n3804 = ( ~n3801 & n3802 ) | ( ~n3801 & n3803 ) | ( n3802 & n3803 ) ;
  assign n3805 = n3799 | n3804 ;
  assign n3806 = ( n3796 & ~n3797 ) | ( n3796 & n3805 ) | ( ~n3797 & n3805 ) ;
  assign n3807 = ~n3485 & n3806 ;
  assign n3808 = ~n3791 & n3807 ;
  assign n3809 = ( n345 & n3791 ) | ( n345 & n3808 ) | ( n3791 & n3808 ) ;
  assign n3810 = n156 & n3290 ;
  assign n3811 = ( x0 & x3 ) | ( x0 & n3810 ) | ( x3 & n3810 ) ;
  assign n3812 = ~x3 & n3811 ;
  assign n3813 = ( ~n3292 & n3809 ) | ( ~n3292 & n3812 ) | ( n3809 & n3812 ) ;
  assign n3814 = x0 & ~n3812 ;
  assign n3815 = ( n3292 & n3813 ) | ( n3292 & ~n3814 ) | ( n3813 & ~n3814 ) ;
  assign n3816 = ( x11 & n391 ) | ( x11 & n3815 ) | ( n391 & n3815 ) ;
  assign n3817 = n3815 & ~n3816 ;
  assign n3818 = ~x8 & n3817 ;
  assign n3819 = ( x5 & ~x9 ) | ( x5 & n3818 ) | ( ~x9 & n3818 ) ;
  assign n3820 = ~x5 & n3819 ;
  assign n3821 = ~x2 & n3820 ;
  assign n3822 = ( x1 & ~x4 ) | ( x1 & n3821 ) | ( ~x4 & n3821 ) ;
  assign n3823 = ~x1 & n3822 ;
  assign n3824 = ( x2 & n676 ) | ( x2 & n1190 ) | ( n676 & n1190 ) ;
  assign n3825 = n1190 & ~n3824 ;
  assign n3826 = x0 & n3825 ;
  assign n3827 = ~x4 & n601 ;
  assign n3828 = ~x3 & n3827 ;
  assign n3829 = ~x1 & n3828 ;
  assign n3830 = ~x2 & n3829 ;
  assign n3831 = ( ~x1 & x3 ) | ( ~x1 & n284 ) | ( x3 & n284 ) ;
  assign n3832 = x1 | n3831 ;
  assign n3833 = ~n3830 & n3832 ;
  assign n3834 = ( n66 & n3830 ) | ( n66 & n3833 ) | ( n3830 & n3833 ) ;
  assign n3835 = x17 & n3834 ;
  assign n3836 = ( x15 & x16 ) | ( x15 & n3835 ) | ( x16 & n3835 ) ;
  assign n3837 = ~x15 & n3836 ;
  assign n3838 = x4 & n3655 ;
  assign n3839 = x1 & ~n123 ;
  assign n3840 = n3838 & n3839 ;
  assign n3841 = ( x1 & ~n135 ) | ( x1 & n230 ) | ( ~n135 & n230 ) ;
  assign n3842 = ~x3 & n3206 ;
  assign n3843 = ~x5 & n296 ;
  assign n3844 = n3842 & n3843 ;
  assign n3845 = x1 & n3844 ;
  assign n3846 = ( n135 & n3841 ) | ( n135 & n3845 ) | ( n3841 & n3845 ) ;
  assign n3847 = x4 | n123 ;
  assign n3848 = x1 & n3847 ;
  assign n3849 = x1 | n3847 ;
  assign n3850 = ~n3848 & n3849 ;
  assign n3851 = n3846 | n3850 ;
  assign n3852 = ( ~n3830 & n3840 ) | ( ~n3830 & n3851 ) | ( n3840 & n3851 ) ;
  assign n3853 = n3830 | n3852 ;
  assign n3854 = ( x18 & ~n136 ) | ( x18 & n3853 ) | ( ~n136 & n3853 ) ;
  assign n3855 = n3853 & ~n3854 ;
  assign n3856 = n3837 | n3855 ;
  assign n3857 = ~x0 & n3856 ;
  assign n3858 = n3826 | n3857 ;
  assign n3859 = ( x36 & ~n215 ) | ( x36 & n3858 ) | ( ~n215 & n3858 ) ;
  assign n3860 = n3858 & ~n3859 ;
  assign n3861 = ~x11 & n3860 ;
  assign n3862 = ( x10 & ~x12 ) | ( x10 & n3861 ) | ( ~x12 & n3861 ) ;
  assign n3863 = ~x10 & n3862 ;
  assign n3864 = ~x8 & n3863 ;
  assign n3865 = ~x9 & n3864 ;
  assign n3866 = ( x40 & n136 ) | ( x40 & n1017 ) | ( n136 & n1017 ) ;
  assign n3867 = x13 & n3866 ;
  assign n3868 = ( ~x13 & x40 ) | ( ~x13 & n3867 ) | ( x40 & n3867 ) ;
  assign n3869 = x14 & n3868 ;
  assign n3870 = ( x5 & x12 ) | ( x5 & n3869 ) | ( x12 & n3869 ) ;
  assign n3871 = ~x5 & n3870 ;
  assign n3872 = ~x3 & n3871 ;
  assign n3873 = ( x2 & ~x4 ) | ( x2 & n3872 ) | ( ~x4 & n3872 ) ;
  assign n3874 = ~x2 & n3873 ;
  assign n3875 = ( ~x15 & x18 ) | ( ~x15 & x19 ) | ( x18 & x19 ) ;
  assign n3876 = x16 | n3875 ;
  assign n3877 = ~x16 & n3875 ;
  assign n3878 = ( x18 & x19 ) | ( x18 & ~n3877 ) | ( x19 & ~n3877 ) ;
  assign n3879 = ( x15 & n3876 ) | ( x15 & ~n3878 ) | ( n3876 & ~n3878 ) ;
  assign n3880 = x17 & n3879 ;
  assign n3881 = n70 & n94 ;
  assign n3882 = x17 | n3881 ;
  assign n3883 = ~n3880 & n3882 ;
  assign n3884 = x40 & n3883 ;
  assign n3885 = ~x5 & n3884 ;
  assign n3886 = ( n79 & n87 ) | ( n79 & ~n3885 ) | ( n87 & ~n3885 ) ;
  assign n3887 = x3 & ~n87 ;
  assign n3888 = ( n3885 & n3886 ) | ( n3885 & ~n3887 ) | ( n3886 & ~n3887 ) ;
  assign n3889 = ( x0 & x13 ) | ( x0 & n3888 ) | ( x13 & n3888 ) ;
  assign n3890 = ~n83 & n85 ;
  assign n3891 = ( x0 & x3 ) | ( x0 & n3890 ) | ( x3 & n3890 ) ;
  assign n3892 = ~x3 & n3891 ;
  assign n3893 = ~x13 & n3892 ;
  assign n3894 = ( n3888 & ~n3889 ) | ( n3888 & n3893 ) | ( ~n3889 & n3893 ) ;
  assign n3895 = ( x2 & n90 ) | ( x2 & n3894 ) | ( n90 & n3894 ) ;
  assign n3896 = ~x2 & n3895 ;
  assign n3897 = ( x1 & ~x14 ) | ( x1 & n3896 ) | ( ~x14 & n3896 ) ;
  assign n3898 = ( x18 & n313 ) | ( x18 & ~n3832 ) | ( n313 & ~n3832 ) ;
  assign n3899 = n3832 & n3898 ;
  assign n3900 = n576 & n3899 ;
  assign n3901 = x5 & n3900 ;
  assign n3902 = x17 | n155 ;
  assign n3903 = n277 & ~n3902 ;
  assign n3904 = ( x3 & n477 ) | ( x3 & n2166 ) | ( n477 & n2166 ) ;
  assign n3905 = ~n3903 & n3904 ;
  assign n3906 = ( n2890 & n3903 ) | ( n2890 & n3905 ) | ( n3903 & n3905 ) ;
  assign n3907 = x12 | n3906 ;
  assign n3908 = x12 & ~n3426 ;
  assign n3909 = n3907 & ~n3908 ;
  assign n3910 = n96 & n576 ;
  assign n3911 = ( x2 & n1236 ) | ( x2 & ~n3910 ) | ( n1236 & ~n3910 ) ;
  assign n3912 = ( x2 & n1236 ) | ( x2 & ~n3909 ) | ( n1236 & ~n3909 ) ;
  assign n3913 = ( n3909 & ~n3911 ) | ( n3909 & n3912 ) | ( ~n3911 & n3912 ) ;
  assign n3914 = x5 | n3913 ;
  assign n3915 = ( ~x5 & n3901 ) | ( ~x5 & n3914 ) | ( n3901 & n3914 ) ;
  assign n3916 = ( ~x0 & x15 ) | ( ~x0 & n3915 ) | ( x15 & n3915 ) ;
  assign n3917 = x12 | x18 ;
  assign n3918 = ( x17 & n135 ) | ( x17 & n3917 ) | ( n135 & n3917 ) ;
  assign n3919 = n135 & ~n3918 ;
  assign n3920 = ( x4 & n493 ) | ( x4 & ~n3919 ) | ( n493 & ~n3919 ) ;
  assign n3921 = ( x4 & ~n58 ) | ( x4 & n493 ) | ( ~n58 & n493 ) ;
  assign n3922 = ( n58 & ~n3920 ) | ( n58 & n3921 ) | ( ~n3920 & n3921 ) ;
  assign n3923 = ( x2 & n1236 ) | ( x2 & ~n3919 ) | ( n1236 & ~n3919 ) ;
  assign n3924 = ( x2 & n1236 ) | ( x2 & ~n3922 ) | ( n1236 & ~n3922 ) ;
  assign n3925 = ( n3922 & ~n3923 ) | ( n3922 & n3924 ) | ( ~n3923 & n3924 ) ;
  assign n3926 = x5 | n3925 ;
  assign n3927 = ~x18 & n3832 ;
  assign n3928 = ( x17 & n135 ) | ( x17 & ~n3927 ) | ( n135 & ~n3927 ) ;
  assign n3929 = n135 & ~n3928 ;
  assign n3930 = ~x12 & n3929 ;
  assign n3931 = x5 & ~n3930 ;
  assign n3932 = n3926 & ~n3931 ;
  assign n3933 = ( x0 & x15 ) | ( x0 & ~n3932 ) | ( x15 & ~n3932 ) ;
  assign n3934 = n3916 & ~n3933 ;
  assign n3935 = x13 & n510 ;
  assign n3936 = ( x13 & n3934 ) | ( x13 & n3935 ) | ( n3934 & n3935 ) ;
  assign n3937 = ~x14 & n3936 ;
  assign n3938 = ( ~x1 & n3897 ) | ( ~x1 & n3937 ) | ( n3897 & n3937 ) ;
  assign n3939 = ( x0 & x1 ) | ( x0 & ~n3938 ) | ( x1 & ~n3938 ) ;
  assign n3940 = n3874 & n3939 ;
  assign n3941 = ( n3874 & n3938 ) | ( n3874 & ~n3940 ) | ( n3938 & ~n3940 ) ;
  assign n3942 = ( x11 & n391 ) | ( x11 & n3941 ) | ( n391 & n3941 ) ;
  assign n3943 = n3941 & ~n3942 ;
  assign n3944 = ~x8 & n3943 ;
  assign n3945 = ~x9 & n3944 ;
  assign n3946 = x15 & n244 ;
  assign n3947 = x14 & n3946 ;
  assign n3948 = ( x4 & n515 ) | ( x4 & n3947 ) | ( n515 & n3947 ) ;
  assign n3949 = ~x4 & n3948 ;
  assign n3950 = ( x1 & ~x17 ) | ( x1 & n3949 ) | ( ~x17 & n3949 ) ;
  assign n3951 = ~x4 & n135 ;
  assign n3952 = n601 & n3951 ;
  assign n3953 = ( x1 & ~x14 ) | ( x1 & n3952 ) | ( ~x14 & n3952 ) ;
  assign n3954 = ( x1 & x14 ) | ( x1 & ~n940 ) | ( x14 & ~n940 ) ;
  assign n3955 = n3953 & ~n3954 ;
  assign n3956 = ~x12 & n3955 ;
  assign n3957 = ( x4 & n239 ) | ( x4 & n515 ) | ( n239 & n515 ) ;
  assign n3958 = ~x4 & n3957 ;
  assign n3959 = n3956 | n3958 ;
  assign n3960 = ( ~x1 & n3956 ) | ( ~x1 & n3959 ) | ( n3956 & n3959 ) ;
  assign n3961 = ( ~x15 & x18 ) | ( ~x15 & n3960 ) | ( x18 & n3960 ) ;
  assign n3962 = x12 & x19 ;
  assign n3963 = ( x14 & x16 ) | ( x14 & ~n3962 ) | ( x16 & ~n3962 ) ;
  assign n3964 = ( ~x12 & x14 ) | ( ~x12 & n3962 ) | ( x14 & n3962 ) ;
  assign n3965 = n3963 & ~n3964 ;
  assign n3966 = ( x15 & ~n487 ) | ( x15 & n3965 ) | ( ~n487 & n3965 ) ;
  assign n3967 = n3965 & ~n3966 ;
  assign n3968 = ~x1 & n3967 ;
  assign n3969 = ~x4 & n3968 ;
  assign n3970 = ~x18 & n3969 ;
  assign n3971 = ( n3960 & ~n3961 ) | ( n3960 & n3970 ) | ( ~n3961 & n3970 ) ;
  assign n3972 = ~x17 & n3971 ;
  assign n3973 = ( ~x1 & n3950 ) | ( ~x1 & n3972 ) | ( n3950 & n3972 ) ;
  assign n3974 = ~n276 & n1276 ;
  assign n3975 = ( ~n66 & n71 ) | ( ~n66 & n3974 ) | ( n71 & n3974 ) ;
  assign n3976 = n66 & n3975 ;
  assign n3977 = x15 | n576 ;
  assign n3978 = x12 | n96 ;
  assign n3979 = ( x15 & n576 ) | ( x15 & ~n3978 ) | ( n576 & ~n3978 ) ;
  assign n3980 = n3977 & ~n3979 ;
  assign n3981 = x14 | n3980 ;
  assign n3982 = ( x15 & x17 ) | ( x15 & n296 ) | ( x17 & n296 ) ;
  assign n3983 = ~x15 & n3982 ;
  assign n3984 = x12 & n3983 ;
  assign n3985 = x14 & ~n3984 ;
  assign n3986 = n3981 & ~n3985 ;
  assign n3987 = ( ~x5 & n3976 ) | ( ~x5 & n3986 ) | ( n3976 & n3986 ) ;
  assign n3988 = x40 & ~n3987 ;
  assign n3989 = ( x40 & n3976 ) | ( x40 & ~n3988 ) | ( n3976 & ~n3988 ) ;
  assign n3990 = ( ~x1 & n3973 ) | ( ~x1 & n3989 ) | ( n3973 & n3989 ) ;
  assign n3991 = x4 | n3990 ;
  assign n3992 = ( ~x4 & n3973 ) | ( ~x4 & n3991 ) | ( n3973 & n3991 ) ;
  assign n3993 = x13 & n3992 ;
  assign n3994 = x16 & n77 ;
  assign n3995 = ( x15 & ~x19 ) | ( x15 & n3875 ) | ( ~x19 & n3875 ) ;
  assign n3996 = ( x17 & ~x19 ) | ( x17 & n3995 ) | ( ~x19 & n3995 ) ;
  assign n3997 = ( ~n477 & n3875 ) | ( ~n477 & n3996 ) | ( n3875 & n3996 ) ;
  assign n3998 = x16 & ~n73 ;
  assign n3999 = ( ~n73 & n3997 ) | ( ~n73 & n3998 ) | ( n3997 & n3998 ) ;
  assign n4000 = ~x14 & n3999 ;
  assign n4001 = ( ~n77 & n3994 ) | ( ~n77 & n4000 ) | ( n3994 & n4000 ) ;
  assign n4002 = x40 & ~n4001 ;
  assign n4003 = x5 | n4002 ;
  assign n4004 = n85 & ~n276 ;
  assign n4005 = x5 & ~n4004 ;
  assign n4006 = n4003 & ~n4005 ;
  assign n4007 = ( x13 & ~n90 ) | ( x13 & n4006 ) | ( ~n90 & n4006 ) ;
  assign n4008 = n4006 & ~n4007 ;
  assign n4009 = n3993 | n4008 ;
  assign n4010 = ( ~x1 & n3993 ) | ( ~x1 & n4009 ) | ( n3993 & n4009 ) ;
  assign n4011 = x0 | n4010 ;
  assign n4012 = ( ~x4 & x14 ) | ( ~x4 & n2161 ) | ( x14 & n2161 ) ;
  assign n4013 = ~x14 & n672 ;
  assign n4014 = ( n2161 & ~n4012 ) | ( n2161 & n4013 ) | ( ~n4012 & n4013 ) ;
  assign n4015 = ~x1 & n4014 ;
  assign n4016 = x0 & ~n4015 ;
  assign n4017 = n4011 & ~n4016 ;
  assign n4018 = x3 | n4017 ;
  assign n4019 = ~x0 & x12 ;
  assign n4020 = ~n608 & n4019 ;
  assign n4021 = n85 & n4020 ;
  assign n4022 = x0 | n4021 ;
  assign n4023 = ( n2161 & n4021 ) | ( n2161 & n4022 ) | ( n4021 & n4022 ) ;
  assign n4024 = x4 | x14 ;
  assign n4025 = ( x5 & n4023 ) | ( x5 & n4024 ) | ( n4023 & n4024 ) ;
  assign n4026 = n4023 & ~n4025 ;
  assign n4027 = ~x1 & n4026 ;
  assign n4028 = x3 & ~n4027 ;
  assign n4029 = n4018 & ~n4028 ;
  assign n4030 = ( x11 & n391 ) | ( x11 & n4029 ) | ( n391 & n4029 ) ;
  assign n4031 = n4029 & ~n4030 ;
  assign n4032 = ~x8 & n4031 ;
  assign n4033 = ( x2 & ~x9 ) | ( x2 & n4032 ) | ( ~x9 & n4032 ) ;
  assign n4034 = ~x2 & n4033 ;
  assign n4035 = x15 & ~n135 ;
  assign n4036 = ~x17 & n4035 ;
  assign n4037 = n665 & n4036 ;
  assign n4038 = x2 & n4037 ;
  assign n4039 = x15 & n51 ;
  assign n4040 = x13 & n4039 ;
  assign n4041 = x13 & n473 ;
  assign n4042 = ~x12 & n4041 ;
  assign n4043 = ( ~x15 & n332 ) | ( ~x15 & n4042 ) | ( n332 & n4042 ) ;
  assign n4044 = n154 & ~n4043 ;
  assign n4045 = ( n154 & n4042 ) | ( n154 & ~n4044 ) | ( n4042 & ~n4044 ) ;
  assign n4046 = ( x17 & x19 ) | ( x17 & n4045 ) | ( x19 & n4045 ) ;
  assign n4047 = x40 & n94 ;
  assign n4048 = ( x17 & ~n154 ) | ( x17 & n4047 ) | ( ~n154 & n4047 ) ;
  assign n4049 = n154 & n4048 ;
  assign n4050 = ~x19 & n4049 ;
  assign n4051 = ( n4045 & ~n4046 ) | ( n4045 & n4050 ) | ( ~n4046 & n4050 ) ;
  assign n4052 = ( x5 & ~x12 ) | ( x5 & n4051 ) | ( ~x12 & n4051 ) ;
  assign n4053 = n4040 & ~n4052 ;
  assign n4054 = ( n4040 & n4051 ) | ( n4040 & ~n4053 ) | ( n4051 & ~n4053 ) ;
  assign n4055 = ( x4 & n493 ) | ( x4 & ~n4037 ) | ( n493 & ~n4037 ) ;
  assign n4056 = ( x4 & n493 ) | ( x4 & ~n4054 ) | ( n493 & ~n4054 ) ;
  assign n4057 = ( n4054 & ~n4055 ) | ( n4054 & n4056 ) | ( ~n4055 & n4056 ) ;
  assign n4058 = x2 | n4057 ;
  assign n4059 = ( ~x2 & n4038 ) | ( ~x2 & n4058 ) | ( n4038 & n4058 ) ;
  assign n4060 = x15 & ~n332 ;
  assign n4061 = ( n169 & n266 ) | ( n169 & ~n4060 ) | ( n266 & ~n4060 ) ;
  assign n4062 = ( x18 & n313 ) | ( x18 & ~n4061 ) | ( n313 & ~n4061 ) ;
  assign n4063 = n4061 & n4062 ;
  assign n4064 = ( x4 & n665 ) | ( x4 & n4063 ) | ( n665 & n4063 ) ;
  assign n4065 = ~x4 & n4064 ;
  assign n4066 = ~x2 & n4065 ;
  assign n4067 = ~x3 & n4066 ;
  assign n4068 = x18 & ~n4067 ;
  assign n4069 = ( n4059 & n4067 ) | ( n4059 & ~n4068 ) | ( n4067 & ~n4068 ) ;
  assign n4070 = x0 | n4069 ;
  assign n4071 = ( x3 & x5 ) | ( x3 & ~x16 ) | ( x5 & ~x16 ) ;
  assign n4072 = ( x3 & x5 ) | ( x3 & n165 ) | ( x5 & n165 ) ;
  assign n4073 = ~n4071 & n4072 ;
  assign n4074 = ( x4 & n665 ) | ( x4 & n4073 ) | ( n665 & n4073 ) ;
  assign n4075 = ~x4 & n4074 ;
  assign n4076 = ~x2 & n4075 ;
  assign n4077 = x0 & ~n4076 ;
  assign n4078 = n4070 & ~n4077 ;
  assign n4079 = ( x1 & x14 ) | ( x1 & n4078 ) | ( x14 & n4078 ) ;
  assign n4080 = x19 & ~n1643 ;
  assign n4081 = ( x5 & x16 ) | ( x5 & ~n4080 ) | ( x16 & ~n4080 ) ;
  assign n4082 = ( n1643 & ~n4080 ) | ( n1643 & n4081 ) | ( ~n4080 & n4081 ) ;
  assign n4083 = x13 & ~n4082 ;
  assign n4084 = ( x15 & x17 ) | ( x15 & n4083 ) | ( x17 & n4083 ) ;
  assign n4085 = ~x17 & n4084 ;
  assign n4086 = ~x4 & n4085 ;
  assign n4087 = ( x3 & ~x12 ) | ( x3 & n4086 ) | ( ~x12 & n4086 ) ;
  assign n4088 = ~x3 & n4087 ;
  assign n4089 = ~x2 & n4088 ;
  assign n4090 = ( x0 & x1 ) | ( x0 & n4089 ) | ( x1 & n4089 ) ;
  assign n4091 = ~x0 & n4090 ;
  assign n4092 = ~x14 & n4091 ;
  assign n4093 = ( n4078 & ~n4079 ) | ( n4078 & n4092 ) | ( ~n4079 & n4092 ) ;
  assign n4094 = x0 | x2 ;
  assign n4095 = x1 | n4094 ;
  assign n4096 = n155 | n4095 ;
  assign n4097 = n515 & ~n4096 ;
  assign n4098 = ~n95 & n1310 ;
  assign n4099 = n1161 & n4098 ;
  assign n4100 = ( n76 & n4097 ) | ( n76 & ~n4099 ) | ( n4097 & ~n4099 ) ;
  assign n4101 = n4097 & ~n4100 ;
  assign n4102 = ~n4093 & n4101 ;
  assign n4103 = ( ~n848 & n4093 ) | ( ~n848 & n4102 ) | ( n4093 & n4102 ) ;
  assign n4104 = ~x9 & n4103 ;
  assign n4105 = ( x8 & ~x10 ) | ( x8 & n4104 ) | ( ~x10 & n4104 ) ;
  assign n4106 = ~x8 & n4105 ;
  assign n4107 = ( x19 & ~n76 ) | ( x19 & n396 ) | ( ~n76 & n396 ) ;
  assign n4108 = n76 & n4107 ;
  assign n4109 = ( x5 & n665 ) | ( x5 & n4108 ) | ( n665 & n4108 ) ;
  assign n4110 = ~x5 & n4109 ;
  assign n4111 = ( x12 & x13 ) | ( x12 & x17 ) | ( x13 & x17 ) ;
  assign n4112 = ( x13 & ~x16 ) | ( x13 & n4111 ) | ( ~x16 & n4111 ) ;
  assign n4113 = x13 & ~n4112 ;
  assign n4114 = n4112 | n4113 ;
  assign n4115 = ( ~x13 & n4113 ) | ( ~x13 & n4114 ) | ( n4113 & n4114 ) ;
  assign n4116 = x40 & n4115 ;
  assign n4117 = x15 & n4116 ;
  assign n4118 = ( x5 & ~x19 ) | ( x5 & n4117 ) | ( ~x19 & n4117 ) ;
  assign n4119 = x15 & n126 ;
  assign n4120 = n559 & n4119 ;
  assign n4121 = ( ~n558 & n559 ) | ( ~n558 & n1149 ) | ( n559 & n1149 ) ;
  assign n4122 = ( x12 & n4120 ) | ( x12 & n4121 ) | ( n4120 & n4121 ) ;
  assign n4123 = ( x5 & x19 ) | ( x5 & ~n4122 ) | ( x19 & ~n4122 ) ;
  assign n4124 = n4118 & ~n4123 ;
  assign n4125 = ( x13 & n487 ) | ( x13 & ~n3980 ) | ( n487 & ~n3980 ) ;
  assign n4126 = n3980 & n4125 ;
  assign n4127 = ( ~n4110 & n4124 ) | ( ~n4110 & n4126 ) | ( n4124 & n4126 ) ;
  assign n4128 = x18 & ~n4126 ;
  assign n4129 = ( n4110 & n4127 ) | ( n4110 & ~n4128 ) | ( n4127 & ~n4128 ) ;
  assign n4130 = ~x14 & n4129 ;
  assign n4131 = ( ~x15 & x40 ) | ( ~x15 & n126 ) | ( x40 & n126 ) ;
  assign n4132 = ( x16 & ~x18 ) | ( x16 & x19 ) | ( ~x18 & x19 ) ;
  assign n4133 = ( ~x17 & x19 ) | ( ~x17 & n4132 ) | ( x19 & n4132 ) ;
  assign n4134 = x19 & ~n4133 ;
  assign n4135 = n4133 | n4134 ;
  assign n4136 = ( ~x19 & n4134 ) | ( ~x19 & n4135 ) | ( n4134 & n4135 ) ;
  assign n4137 = ( x15 & x40 ) | ( x15 & n4136 ) | ( x40 & n4136 ) ;
  assign n4138 = n4131 & n4137 ;
  assign n4139 = ( x13 & n2684 ) | ( x13 & ~n4138 ) | ( n2684 & ~n4138 ) ;
  assign n4140 = n4138 & n4139 ;
  assign n4141 = n4130 | n4140 ;
  assign n4142 = ( ~x5 & n4130 ) | ( ~x5 & n4141 ) | ( n4130 & n4141 ) ;
  assign n4143 = ( x0 & x1 ) | ( x0 & n4142 ) | ( x1 & n4142 ) ;
  assign n4144 = x5 & n1237 ;
  assign n4145 = ( x1 & ~n1755 ) | ( x1 & n4144 ) | ( ~n1755 & n4144 ) ;
  assign n4146 = n1755 & n4145 ;
  assign n4147 = ~x0 & n4146 ;
  assign n4148 = ( n4142 & ~n4143 ) | ( n4142 & n4147 ) | ( ~n4143 & n4147 ) ;
  assign n4149 = x0 & x5 ;
  assign n4150 = ( x1 & n665 ) | ( x1 & n4149 ) | ( n665 & n4149 ) ;
  assign n4151 = ~x1 & n4150 ;
  assign n4152 = n96 & n4151 ;
  assign n4153 = ( x14 & n110 ) | ( x14 & n4152 ) | ( n110 & n4152 ) ;
  assign n4154 = ~x14 & n4153 ;
  assign n4155 = ~n4148 & n4154 ;
  assign n4156 = ( ~n848 & n4148 ) | ( ~n848 & n4155 ) | ( n4148 & n4155 ) ;
  assign n4157 = ~x9 & n4156 ;
  assign n4158 = ( x8 & ~x10 ) | ( x8 & n4157 ) | ( ~x10 & n4157 ) ;
  assign n4159 = ~x8 & n4158 ;
  assign n4160 = ~x3 & n4159 ;
  assign n4161 = ( x2 & ~x4 ) | ( x2 & n4160 ) | ( ~x4 & n4160 ) ;
  assign n4162 = ~x2 & n4161 ;
  assign n4163 = n90 & n1311 ;
  assign n4164 = ( n159 & n1117 ) | ( n159 & ~n4163 ) | ( n1117 & ~n4163 ) ;
  assign n4165 = n1117 & ~n4164 ;
  assign n4166 = ( x15 & ~x17 ) | ( x15 & x18 ) | ( ~x17 & x18 ) ;
  assign n4167 = ( ~x16 & x18 ) | ( ~x16 & n4166 ) | ( x18 & n4166 ) ;
  assign n4168 = x18 & ~n4167 ;
  assign n4169 = n4167 | n4168 ;
  assign n4170 = ( ~x18 & n4168 ) | ( ~x18 & n4169 ) | ( n4168 & n4169 ) ;
  assign n4171 = ( ~x4 & x19 ) | ( ~x4 & n4170 ) | ( x19 & n4170 ) ;
  assign n4172 = ( x4 & x19 ) | ( x4 & n484 ) | ( x19 & n484 ) ;
  assign n4173 = n4171 & n4172 ;
  assign n4174 = ( ~x4 & n110 ) | ( ~x4 & n4173 ) | ( n110 & n4173 ) ;
  assign n4175 = n4098 & ~n4174 ;
  assign n4176 = ( n4098 & n4173 ) | ( n4098 & ~n4175 ) | ( n4173 & ~n4175 ) ;
  assign n4177 = x12 | n4176 ;
  assign n4178 = ( x15 & x40 ) | ( x15 & n477 ) | ( x40 & n477 ) ;
  assign n4179 = ~n1938 & n4178 ;
  assign n4180 = ( x40 & n1938 ) | ( x40 & n4179 ) | ( n1938 & n4179 ) ;
  assign n4181 = ~x4 & n4180 ;
  assign n4182 = x12 & ~n4181 ;
  assign n4183 = n4177 & ~n4182 ;
  assign n4184 = ( ~x13 & x14 ) | ( ~x13 & n4183 ) | ( x14 & n4183 ) ;
  assign n4185 = ( ~x15 & x17 ) | ( ~x15 & x40 ) | ( x17 & x40 ) ;
  assign n4186 = ( ~x15 & x17 ) | ( ~x15 & x19 ) | ( x17 & x19 ) ;
  assign n4187 = n4185 & ~n4186 ;
  assign n4188 = ~x16 & n4187 ;
  assign n4189 = ( x13 & ~x18 ) | ( x13 & n4188 ) | ( ~x18 & n4188 ) ;
  assign n4190 = ~x13 & n4189 ;
  assign n4191 = n90 & n4190 ;
  assign n4192 = ~x14 & n4191 ;
  assign n4193 = ( n4183 & ~n4184 ) | ( n4183 & n4192 ) | ( ~n4184 & n4192 ) ;
  assign n4194 = n635 & n1035 ;
  assign n4195 = ( n43 & n1237 ) | ( n43 & n4194 ) | ( n1237 & n4194 ) ;
  assign n4196 = ~n43 & n4195 ;
  assign n4197 = ( ~n4165 & n4193 ) | ( ~n4165 & n4196 ) | ( n4193 & n4196 ) ;
  assign n4198 = x5 & ~n4196 ;
  assign n4199 = ( n4165 & n4197 ) | ( n4165 & ~n4198 ) | ( n4197 & ~n4198 ) ;
  assign n4200 = ( x11 & n391 ) | ( x11 & n4199 ) | ( n391 & n4199 ) ;
  assign n4201 = n4199 & ~n4200 ;
  assign n4202 = ~x8 & n4201 ;
  assign n4203 = ( x3 & ~x9 ) | ( x3 & n4202 ) | ( ~x9 & n4202 ) ;
  assign n4204 = ~x3 & n4203 ;
  assign n4205 = ~x1 & n4204 ;
  assign n4206 = ( x0 & ~x2 ) | ( x0 & n4205 ) | ( ~x2 & n4205 ) ;
  assign n4207 = ~x0 & n4206 ;
  assign n4208 = ( x14 & x17 ) | ( x14 & ~n952 ) | ( x17 & ~n952 ) ;
  assign n4209 = x16 & n4208 ;
  assign n4210 = ( x14 & ~x16 ) | ( x14 & n4209 ) | ( ~x16 & n4209 ) ;
  assign n4211 = ( x15 & n196 ) | ( x15 & n4210 ) | ( n196 & n4210 ) ;
  assign n4212 = ~n4210 & n4211 ;
  assign n4213 = x13 & n4212 ;
  assign n4214 = ( x11 & x12 ) | ( x11 & n4213 ) | ( x12 & n4213 ) ;
  assign n4215 = ~x11 & n4214 ;
  assign n4216 = ~x9 & n4215 ;
  assign n4217 = ( x8 & ~x10 ) | ( x8 & n4216 ) | ( ~x10 & n4216 ) ;
  assign n4218 = ~x8 & n4217 ;
  assign n4219 = ~x4 & n4218 ;
  assign n4220 = ( x3 & ~x5 ) | ( x3 & n4219 ) | ( ~x5 & n4219 ) ;
  assign n4221 = ~x3 & n4220 ;
  assign n4222 = ~x1 & n4221 ;
  assign n4223 = ( x0 & ~x2 ) | ( x0 & n4222 ) | ( ~x2 & n4222 ) ;
  assign n4224 = ~x0 & n4223 ;
  assign n4225 = ( x15 & n76 ) | ( x15 & n477 ) | ( n76 & n477 ) ;
  assign n4226 = x40 & n4225 ;
  assign n4227 = x12 & n4226 ;
  assign n4228 = ( x4 & ~x5 ) | ( x4 & n4227 ) | ( ~x5 & n4227 ) ;
  assign n4229 = x19 & n4170 ;
  assign n4230 = ~x12 & n4229 ;
  assign n4231 = ( x4 & x5 ) | ( x4 & ~n4230 ) | ( x5 & ~n4230 ) ;
  assign n4232 = n4228 & ~n4231 ;
  assign n4233 = n1035 & n2418 ;
  assign n4234 = ~n42 & n4233 ;
  assign n4235 = n126 & n4234 ;
  assign n4236 = ~n4232 & n4235 ;
  assign n4237 = x14 | x36 ;
  assign n4238 = ( n4232 & n4236 ) | ( n4232 & ~n4237 ) | ( n4236 & ~n4237 ) ;
  assign n4239 = ~x11 & x13 ;
  assign n4240 = ( x10 & n4238 ) | ( x10 & n4239 ) | ( n4238 & n4239 ) ;
  assign n4241 = ~x10 & n4240 ;
  assign n4242 = ~x8 & n4241 ;
  assign n4243 = ( x3 & ~x9 ) | ( x3 & n4242 ) | ( ~x9 & n4242 ) ;
  assign n4244 = ~x3 & n4243 ;
  assign n4245 = ~x1 & n4244 ;
  assign n4246 = ( x0 & ~x2 ) | ( x0 & n4245 ) | ( ~x2 & n4245 ) ;
  assign n4247 = ~x0 & n4246 ;
  assign n4248 = ( n43 & ~n796 ) | ( n43 & n4194 ) | ( ~n796 & n4194 ) ;
  assign n4249 = ~n43 & n4248 ;
  assign n4250 = ~x17 & n277 ;
  assign n4251 = x16 & n4250 ;
  assign n4252 = ( x4 & x19 ) | ( x4 & n4251 ) | ( x19 & n4251 ) ;
  assign n4253 = n4171 & n4252 ;
  assign n4254 = ( ~x4 & n94 ) | ( ~x4 & n4253 ) | ( n94 & n4253 ) ;
  assign n4255 = n4098 & ~n4254 ;
  assign n4256 = ( n4098 & n4253 ) | ( n4098 & ~n4255 ) | ( n4253 & ~n4255 ) ;
  assign n4257 = x12 | n4256 ;
  assign n4258 = ( x40 & n1221 ) | ( x40 & n1938 ) | ( n1221 & n1938 ) ;
  assign n4259 = ~x4 & n4258 ;
  assign n4260 = x12 & ~n4259 ;
  assign n4261 = n4257 & ~n4260 ;
  assign n4262 = ( x5 & x14 ) | ( x5 & n4261 ) | ( x14 & n4261 ) ;
  assign n4263 = n90 & n3185 ;
  assign n4264 = ~x5 & n4263 ;
  assign n4265 = ( n4261 & ~n4262 ) | ( n4261 & n4264 ) | ( ~n4262 & n4264 ) ;
  assign n4266 = n156 & n1035 ;
  assign n4267 = n3290 & n4266 ;
  assign n4268 = ( ~n4249 & n4265 ) | ( ~n4249 & n4267 ) | ( n4265 & n4267 ) ;
  assign n4269 = x13 | n4267 ;
  assign n4270 = ( n4249 & n4268 ) | ( n4249 & n4269 ) | ( n4268 & n4269 ) ;
  assign n4271 = ( x11 & n391 ) | ( x11 & n4270 ) | ( n391 & n4270 ) ;
  assign n4272 = n4270 & ~n4271 ;
  assign n4273 = ~x8 & n4272 ;
  assign n4274 = ( x3 & ~x9 ) | ( x3 & n4273 ) | ( ~x9 & n4273 ) ;
  assign n4275 = ~x3 & n4274 ;
  assign n4276 = ~x1 & n4275 ;
  assign n4277 = ( x0 & ~x2 ) | ( x0 & n4276 ) | ( ~x2 & n4276 ) ;
  assign n4278 = ~x0 & n4277 ;
  assign n4279 = x40 & ~n135 ;
  assign n4280 = ~x17 & n4279 ;
  assign n4281 = x15 & n4280 ;
  assign n4282 = ( x12 & x13 ) | ( x12 & n4281 ) | ( x13 & n4281 ) ;
  assign n4283 = ~x12 & n4282 ;
  assign n4284 = x5 | n4283 ;
  assign n4285 = n153 & n1553 ;
  assign n4286 = x5 & ~n4285 ;
  assign n4287 = n4284 & ~n4286 ;
  assign n4288 = ( x18 & n4237 ) | ( x18 & n4287 ) | ( n4237 & n4287 ) ;
  assign n4289 = n4287 & ~n4288 ;
  assign n4290 = ~x10 & n4289 ;
  assign n4291 = ( x9 & ~x11 ) | ( x9 & n4290 ) | ( ~x11 & n4290 ) ;
  assign n4292 = ~x9 & n4291 ;
  assign n4293 = ~x4 & n4292 ;
  assign n4294 = ( x3 & ~x8 ) | ( x3 & n4293 ) | ( ~x8 & n4293 ) ;
  assign n4295 = ~x3 & n4294 ;
  assign n4296 = ~x1 & n4295 ;
  assign n4297 = ( x0 & ~x2 ) | ( x0 & n4296 ) | ( ~x2 & n4296 ) ;
  assign n4298 = ~x0 & n4297 ;
  assign n4299 = ( x40 & n126 ) | ( x40 & n714 ) | ( n126 & n714 ) ;
  assign n4300 = x13 & n4299 ;
  assign n4301 = ( x15 & x36 ) | ( x15 & n4300 ) | ( x36 & n4300 ) ;
  assign n4302 = ~x36 & n4301 ;
  assign n4303 = ( x10 & n198 ) | ( x10 & n4302 ) | ( n198 & n4302 ) ;
  assign n4304 = ~x10 & n4303 ;
  assign n4305 = ~x8 & n4304 ;
  assign n4306 = ( x5 & ~x9 ) | ( x5 & n4305 ) | ( ~x9 & n4305 ) ;
  assign n4307 = ~x5 & n4306 ;
  assign n4308 = ~x3 & n4307 ;
  assign n4309 = ( x2 & ~x4 ) | ( x2 & n4308 ) | ( ~x4 & n4308 ) ;
  assign n4310 = ~x2 & n4309 ;
  assign n4311 = ~x0 & n4310 ;
  assign n4312 = ~x1 & n4311 ;
  assign n4313 = x3 | n2310 ;
  assign n4314 = ( ~x2 & x4 ) | ( ~x2 & n4313 ) | ( x4 & n4313 ) ;
  assign n4315 = x2 | n4314 ;
  assign n4316 = x5 & ~x9 ;
  assign n4317 = ( x8 & ~n4315 ) | ( x8 & n4316 ) | ( ~n4315 & n4316 ) ;
  assign n4318 = ~x8 & n4317 ;
  assign n4319 = ~x11 & n4318 ;
  assign n4320 = ( x10 & ~x12 ) | ( x10 & n4319 ) | ( ~x12 & n4319 ) ;
  assign n4321 = ~x10 & n4320 ;
  assign n4322 = ( x14 & n192 ) | ( x14 & n4321 ) | ( n192 & n4321 ) ;
  assign n4323 = ~x14 & n4322 ;
  assign n4324 = x16 & n4323 ;
  assign n4325 = ( x17 & x18 ) | ( x17 & n4324 ) | ( x18 & n4324 ) ;
  assign n4326 = ~x18 & n4325 ;
  assign n4327 = ~x19 & n4326 ;
  assign n4328 = ~x36 & n4327 ;
  assign n4329 = ~x8 & n2836 ;
  assign n4330 = ( x5 & ~x9 ) | ( x5 & n4329 ) | ( ~x9 & n4329 ) ;
  assign n4331 = ~x5 & n4330 ;
  assign n4332 = ~x3 & n4331 ;
  assign n4333 = ( x2 & ~x4 ) | ( x2 & n4332 ) | ( ~x4 & n4332 ) ;
  assign n4334 = ~x2 & n4333 ;
  assign n4335 = ~x0 & n4334 ;
  assign n4336 = ~x1 & n4335 ;
  assign n4337 = n1242 & n1270 ;
  assign n4338 = n665 & n4337 ;
  assign n4339 = ( x5 & ~x12 ) | ( x5 & x15 ) | ( ~x12 & x15 ) ;
  assign n4340 = ( x5 & ~x14 ) | ( x5 & n4339 ) | ( ~x14 & n4339 ) ;
  assign n4341 = x5 & ~n4340 ;
  assign n4342 = n4340 | n4341 ;
  assign n4343 = ( ~x5 & n4341 ) | ( ~x5 & n4342 ) | ( n4341 & n4342 ) ;
  assign n4344 = ( x16 & n416 ) | ( x16 & ~n4343 ) | ( n416 & ~n4343 ) ;
  assign n4345 = n4343 & n4344 ;
  assign n4346 = ~x17 & n745 ;
  assign n4347 = x5 & x13 ;
  assign n4348 = x5 & ~n4347 ;
  assign n4349 = n4346 & n4348 ;
  assign n4350 = x15 & x17 ;
  assign n4351 = ~x14 & n4350 ;
  assign n4352 = ( ~n4347 & n4348 ) | ( ~n4347 & n4351 ) | ( n4348 & n4351 ) ;
  assign n4353 = ( x13 & n4349 ) | ( x13 & n4352 ) | ( n4349 & n4352 ) ;
  assign n4354 = x12 | n4353 ;
  assign n4355 = n1115 | n1161 ;
  assign n4356 = ( n570 & n1115 ) | ( n570 & n4355 ) | ( n1115 & n4355 ) ;
  assign n4357 = x5 & n4356 ;
  assign n4358 = x12 & ~n4357 ;
  assign n4359 = n4354 & ~n4358 ;
  assign n4360 = x14 & n558 ;
  assign n4361 = ( x5 & ~n4350 ) | ( x5 & n4360 ) | ( ~n4350 & n4360 ) ;
  assign n4362 = n4350 & n4361 ;
  assign n4363 = x5 & ~x14 ;
  assign n4364 = ( ~x5 & n1090 ) | ( ~x5 & n4363 ) | ( n1090 & n4363 ) ;
  assign n4365 = ( ~n185 & n1090 ) | ( ~n185 & n4364 ) | ( n1090 & n4364 ) ;
  assign n4366 = ( x12 & ~n4362 ) | ( x12 & n4365 ) | ( ~n4362 & n4365 ) ;
  assign n4367 = ~x13 & n4366 ;
  assign n4368 = ( x13 & ~n4362 ) | ( x13 & n4367 ) | ( ~n4362 & n4367 ) ;
  assign n4369 = ~x16 & n4368 ;
  assign n4370 = ( ~n4359 & n4368 ) | ( ~n4359 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4371 = ~x13 & n4370 ;
  assign n4372 = ( ~n4345 & n4370 ) | ( ~n4345 & n4371 ) | ( n4370 & n4371 ) ;
  assign n4373 = ( x3 & ~n4338 ) | ( x3 & n4372 ) | ( ~n4338 & n4372 ) ;
  assign n4374 = x40 & n4373 ;
  assign n4375 = ( x40 & n4338 ) | ( x40 & ~n4374 ) | ( n4338 & ~n4374 ) ;
  assign n4376 = ( x5 & n85 ) | ( x5 & n1117 ) | ( n85 & n1117 ) ;
  assign n4377 = ~x5 & n4376 ;
  assign n4378 = n190 & ~n1867 ;
  assign n4379 = n43 | n76 ;
  assign n4380 = n4378 & ~n4379 ;
  assign n4381 = ( n1130 & ~n4377 ) | ( n1130 & n4380 ) | ( ~n4377 & n4380 ) ;
  assign n4382 = x12 | n4380 ;
  assign n4383 = ( n4377 & n4381 ) | ( n4377 & n4382 ) | ( n4381 & n4382 ) ;
  assign n4384 = ( ~x3 & n4375 ) | ( ~x3 & n4383 ) | ( n4375 & n4383 ) ;
  assign n4385 = x40 & ~n4384 ;
  assign n4386 = ( x40 & n4375 ) | ( x40 & ~n4385 ) | ( n4375 & ~n4385 ) ;
  assign n4387 = x8 | n4386 ;
  assign n4388 = x8 & n2349 ;
  assign n4389 = n4387 & ~n4388 ;
  assign n4390 = x11 | n4389 ;
  assign n4391 = x8 & ~n2349 ;
  assign n4392 = x11 & ~n4391 ;
  assign n4393 = n4390 & ~n4392 ;
  assign n4394 = ( x10 & x36 ) | ( x10 & n4393 ) | ( x36 & n4393 ) ;
  assign n4395 = ~x5 & x10 ;
  assign n4396 = ( x3 & x8 ) | ( x3 & n4395 ) | ( x8 & n4395 ) ;
  assign n4397 = ~x3 & n4396 ;
  assign n4398 = ~x36 & n4397 ;
  assign n4399 = ( n4393 & ~n4394 ) | ( n4393 & n4398 ) | ( ~n4394 & n4398 ) ;
  assign n4400 = ~x4 & n4399 ;
  assign n4401 = ( x2 & ~x9 ) | ( x2 & n4400 ) | ( ~x9 & n4400 ) ;
  assign n4402 = ~x2 & n4401 ;
  assign n4403 = ~x0 & n4402 ;
  assign n4404 = ~x1 & n4403 ;
  assign n4405 = x15 & ~x39 ;
  assign n4406 = ( x17 & x18 ) | ( x17 & n4405 ) | ( x18 & n4405 ) ;
  assign n4407 = ~x17 & n4406 ;
  assign n4408 = n559 & n4407 ;
  assign n4409 = x17 | x39 ;
  assign n4410 = x15 & n4409 ;
  assign n4411 = ( n313 & n1304 ) | ( n313 & ~n4410 ) | ( n1304 & ~n4410 ) ;
  assign n4412 = ~x18 & n4411 ;
  assign n4413 = ( ~n558 & n559 ) | ( ~n558 & n4412 ) | ( n559 & n4412 ) ;
  assign n4414 = ( x12 & n4408 ) | ( x12 & n4413 ) | ( n4408 & n4413 ) ;
  assign n4415 = ( x37 & n2826 ) | ( x37 & ~n4414 ) | ( n2826 & ~n4414 ) ;
  assign n4416 = n4414 & n4415 ;
  assign n4417 = ~x14 & n4416 ;
  assign n4418 = ( x11 & ~x16 ) | ( x11 & n4417 ) | ( ~x16 & n4417 ) ;
  assign n4419 = ~x11 & n4418 ;
  assign n4420 = ( x10 & ~x36 ) | ( x10 & n4419 ) | ( ~x36 & n4419 ) ;
  assign n4421 = x8 & ~x36 ;
  assign n4422 = ( ~x10 & n4420 ) | ( ~x10 & n4421 ) | ( n4420 & n4421 ) ;
  assign n4423 = ~x5 & n4422 ;
  assign n4424 = ( x4 & ~x9 ) | ( x4 & n4423 ) | ( ~x9 & n4423 ) ;
  assign n4425 = ~x4 & n4424 ;
  assign n4426 = ~x2 & n4425 ;
  assign n4427 = ( x1 & ~x3 ) | ( x1 & n4426 ) | ( ~x3 & n4426 ) ;
  assign n4428 = ~x1 & n4427 ;
  assign n4429 = ~x0 & n4428 ;
  assign n4430 = x8 | n4315 ;
  assign n4431 = ( ~x5 & x9 ) | ( ~x5 & n4430 ) | ( x9 & n4430 ) ;
  assign n4432 = x5 | n4431 ;
  assign n4433 = x11 | n4432 ;
  assign n4434 = ( ~x10 & x12 ) | ( ~x10 & n4433 ) | ( x12 & n4433 ) ;
  assign n4435 = x10 | n4434 ;
  assign n4436 = ( x14 & n1822 ) | ( x14 & ~n4435 ) | ( n1822 & ~n4435 ) ;
  assign n4437 = ~x14 & n4436 ;
  assign n4438 = ( x16 & n416 ) | ( x16 & n4437 ) | ( n416 & n4437 ) ;
  assign n4439 = ~x16 & n4438 ;
  assign n4440 = x19 & ~x37 ;
  assign n4441 = ( x36 & n4439 ) | ( x36 & n4440 ) | ( n4439 & n4440 ) ;
  assign n4442 = ~x36 & n4441 ;
  assign n4443 = ~x39 & x40 ;
  assign n4444 = ( x38 & n4442 ) | ( x38 & n4443 ) | ( n4442 & n4443 ) ;
  assign n4445 = ~x38 & n4444 ;
  assign n4446 = ( ~x13 & x16 ) | ( ~x13 & n96 ) | ( x16 & n96 ) ;
  assign n4447 = ( ~x16 & n190 ) | ( ~x16 & n4446 ) | ( n190 & n4446 ) ;
  assign n4448 = x17 & ~n135 ;
  assign n4449 = ~x14 & n4448 ;
  assign n4450 = ( x13 & ~x18 ) | ( x13 & n4449 ) | ( ~x18 & n4449 ) ;
  assign n4451 = ( x14 & x16 ) | ( x14 & ~x17 ) | ( x16 & ~x17 ) ;
  assign n4452 = ( x14 & ~x19 ) | ( x14 & n4451 ) | ( ~x19 & n4451 ) ;
  assign n4453 = x14 & ~n4452 ;
  assign n4454 = n4452 | n4453 ;
  assign n4455 = ( ~x14 & n4453 ) | ( ~x14 & n4454 ) | ( n4453 & n4454 ) ;
  assign n4456 = ( x13 & x18 ) | ( x13 & ~n4455 ) | ( x18 & ~n4455 ) ;
  assign n4457 = n4450 & ~n4456 ;
  assign n4458 = x14 & ~n2553 ;
  assign n4459 = ( n1025 & n2553 ) | ( n1025 & n4458 ) | ( n2553 & n4458 ) ;
  assign n4460 = ( ~n4447 & n4457 ) | ( ~n4447 & n4459 ) | ( n4457 & n4459 ) ;
  assign n4461 = x15 & ~n4459 ;
  assign n4462 = ( n4447 & n4460 ) | ( n4447 & ~n4461 ) | ( n4460 & ~n4461 ) ;
  assign n4463 = x14 & n209 ;
  assign n4464 = x13 & n4463 ;
  assign n4465 = x16 & n477 ;
  assign n4466 = ( x13 & ~n276 ) | ( x13 & n4465 ) | ( ~n276 & n4465 ) ;
  assign n4467 = ~x13 & n4466 ;
  assign n4468 = ( x12 & n4464 ) | ( x12 & n4467 ) | ( n4464 & n4467 ) ;
  assign n4469 = ~n4462 & n4468 ;
  assign n4470 = ( x12 & n4462 ) | ( x12 & n4469 ) | ( n4462 & n4469 ) ;
  assign n4471 = n84 & n304 ;
  assign n4472 = ( ~n70 & n665 ) | ( ~n70 & n4471 ) | ( n665 & n4471 ) ;
  assign n4473 = n70 & n4472 ;
  assign n4474 = ~n4470 & n4473 ;
  assign n4475 = ( n345 & n4470 ) | ( n345 & n4474 ) | ( n4470 & n4474 ) ;
  assign n4476 = ( ~n3292 & n3812 ) | ( ~n3292 & n4475 ) | ( n3812 & n4475 ) ;
  assign n4477 = ( n3292 & ~n3814 ) | ( n3292 & n4476 ) | ( ~n3814 & n4476 ) ;
  assign n4478 = ( x11 & n391 ) | ( x11 & n4477 ) | ( n391 & n4477 ) ;
  assign n4479 = n4477 & ~n4478 ;
  assign n4480 = ~x8 & n4479 ;
  assign n4481 = ( x5 & ~x9 ) | ( x5 & n4480 ) | ( ~x9 & n4480 ) ;
  assign n4482 = ~x5 & n4481 ;
  assign n4483 = ~x2 & n4482 ;
  assign n4484 = ( x1 & ~x4 ) | ( x1 & n4483 ) | ( ~x4 & n4483 ) ;
  assign n4485 = ~x1 & n4484 ;
  assign n4486 = ( x4 & ~n601 ) | ( x4 & n3642 ) | ( ~n601 & n3642 ) ;
  assign n4487 = x24 & x40 ;
  assign n4488 = ( ~x23 & x26 ) | ( ~x23 & n4487 ) | ( x26 & n4487 ) ;
  assign n4489 = x23 & n4488 ;
  assign n4490 = ~x20 & n4489 ;
  assign n4491 = ( x5 & n1818 ) | ( x5 & n4490 ) | ( n1818 & n4490 ) ;
  assign n4492 = ~x5 & n4491 ;
  assign n4493 = ~x4 & n4492 ;
  assign n4494 = ( n3642 & ~n4486 ) | ( n3642 & n4493 ) | ( ~n4486 & n4493 ) ;
  assign n4495 = ( x2 & x27 ) | ( x2 & n4494 ) | ( x27 & n4494 ) ;
  assign n4496 = ( x2 & x4 ) | ( x2 & ~x20 ) | ( x4 & ~x20 ) ;
  assign n4497 = ( x2 & x4 ) | ( x2 & ~x21 ) | ( x4 & ~x21 ) ;
  assign n4498 = ~n4496 & n4497 ;
  assign n4499 = ( ~x2 & n564 ) | ( ~x2 & n4498 ) | ( n564 & n4498 ) ;
  assign n4500 = x4 & ~n4499 ;
  assign n4501 = ( x4 & n4498 ) | ( x4 & ~n4500 ) | ( n4498 & ~n4500 ) ;
  assign n4502 = x27 & n4501 ;
  assign n4503 = ( ~x2 & n4495 ) | ( ~x2 & n4502 ) | ( n4495 & n4502 ) ;
  assign n4504 = ( x27 & n566 ) | ( x27 & ~n601 ) | ( n566 & ~n601 ) ;
  assign n4505 = ( x22 & ~x23 ) | ( x22 & x40 ) | ( ~x23 & x40 ) ;
  assign n4506 = ( x23 & n4487 ) | ( x23 & n4505 ) | ( n4487 & n4505 ) ;
  assign n4507 = ( x5 & n562 ) | ( x5 & n4506 ) | ( n562 & n4506 ) ;
  assign n4508 = ~x5 & n4507 ;
  assign n4509 = ~x27 & n4508 ;
  assign n4510 = ( n566 & ~n4504 ) | ( n566 & n4509 ) | ( ~n4504 & n4509 ) ;
  assign n4511 = ( ~x5 & n3647 ) | ( ~x5 & n4510 ) | ( n3647 & n4510 ) ;
  assign n4512 = x20 & ~n4511 ;
  assign n4513 = ( x20 & n4510 ) | ( x20 & ~n4512 ) | ( n4510 & ~n4512 ) ;
  assign n4514 = ( ~x2 & n4503 ) | ( ~x2 & n4513 ) | ( n4503 & n4513 ) ;
  assign n4515 = x4 | n4514 ;
  assign n4516 = ( ~x4 & n4503 ) | ( ~x4 & n4515 ) | ( n4503 & n4515 ) ;
  assign n4517 = ( ~x18 & x19 ) | ( ~x18 & n4516 ) | ( x19 & n4516 ) ;
  assign n4518 = ~x4 & n1416 ;
  assign n4519 = ( x2 & ~x5 ) | ( x2 & n4518 ) | ( ~x5 & n4518 ) ;
  assign n4520 = ~x2 & n4519 ;
  assign n4521 = x18 & n4520 ;
  assign n4522 = ( n4516 & ~n4517 ) | ( n4516 & n4521 ) | ( ~n4517 & n4521 ) ;
  assign n4523 = ( ~x3 & x16 ) | ( ~x3 & n4522 ) | ( x16 & n4522 ) ;
  assign n4524 = ~n129 & n797 ;
  assign n4525 = ( x2 & n1416 ) | ( x2 & n4524 ) | ( n1416 & n4524 ) ;
  assign n4526 = ~x2 & n4525 ;
  assign n4527 = ~x3 & n4526 ;
  assign n4528 = ( ~x16 & n4523 ) | ( ~x16 & n4527 ) | ( n4523 & n4527 ) ;
  assign n4529 = ~x16 & n250 ;
  assign n4530 = ( x4 & x5 ) | ( x4 & n4529 ) | ( x5 & n4529 ) ;
  assign n4531 = ~x4 & n4530 ;
  assign n4532 = ( n878 & n4528 ) | ( n878 & n4531 ) | ( n4528 & n4531 ) ;
  assign n4533 = n1061 & ~n4532 ;
  assign n4534 = ( n1061 & n4528 ) | ( n1061 & ~n4533 ) | ( n4528 & ~n4533 ) ;
  assign n4535 = ( x36 & ~n570 ) | ( x36 & n4534 ) | ( ~n570 & n4534 ) ;
  assign n4536 = n4534 & ~n4535 ;
  assign n4537 = ( x13 & n383 ) | ( x13 & n4536 ) | ( n383 & n4536 ) ;
  assign n4538 = ~x13 & n4537 ;
  assign n4539 = ~x10 & n4538 ;
  assign n4540 = ( x9 & ~x11 ) | ( x9 & n4539 ) | ( ~x11 & n4539 ) ;
  assign n4541 = ~x9 & n4540 ;
  assign n4542 = ~x1 & n4541 ;
  assign n4543 = ( x0 & ~x8 ) | ( x0 & n4542 ) | ( ~x8 & n4542 ) ;
  assign n4544 = ~x0 & n4543 ;
  assign n4545 = ( x5 & x24 ) | ( x5 & ~x27 ) | ( x24 & ~x27 ) ;
  assign n4546 = x5 & x24 ;
  assign n4547 = ( x3 & x27 ) | ( x3 & ~n4546 ) | ( x27 & ~n4546 ) ;
  assign n4548 = n4545 & n4547 ;
  assign n4549 = ( x2 & ~x4 ) | ( x2 & n4548 ) | ( ~x4 & n4548 ) ;
  assign n4550 = x2 & ~x5 ;
  assign n4551 = ( x3 & n1742 ) | ( x3 & n4550 ) | ( n1742 & n4550 ) ;
  assign n4552 = ~x3 & n4551 ;
  assign n4553 = ~x4 & n4552 ;
  assign n4554 = ( ~x2 & n4549 ) | ( ~x2 & n4553 ) | ( n4549 & n4553 ) ;
  assign n4555 = x3 & n3206 ;
  assign n4556 = ( n1742 & n4554 ) | ( n1742 & n4555 ) | ( n4554 & n4555 ) ;
  assign n4557 = x5 & ~n4556 ;
  assign n4558 = ( x5 & n4554 ) | ( x5 & ~n4557 ) | ( n4554 & ~n4557 ) ;
  assign n4559 = x4 & ~n1044 ;
  assign n4560 = x4 | n3700 ;
  assign n4561 = ~n4559 & n4560 ;
  assign n4562 = ( x4 & x23 ) | ( x4 & n3235 ) | ( x23 & n3235 ) ;
  assign n4563 = ~x4 & n4562 ;
  assign n4564 = x27 | n4563 ;
  assign n4565 = ( n4561 & n4563 ) | ( n4561 & n4564 ) | ( n4563 & n4564 ) ;
  assign n4566 = x5 | n4565 ;
  assign n4567 = ~x4 & n1366 ;
  assign n4568 = x5 & ~n4567 ;
  assign n4569 = n4566 & ~n4568 ;
  assign n4570 = x3 & n4569 ;
  assign n4571 = ~x2 & n4570 ;
  assign n4572 = n561 & ~n4571 ;
  assign n4573 = ( n4558 & n4571 ) | ( n4558 & ~n4572 ) | ( n4571 & ~n4572 ) ;
  assign n4574 = ( x18 & n562 ) | ( x18 & ~n4573 ) | ( n562 & ~n4573 ) ;
  assign n4575 = n4573 & n4574 ;
  assign n4576 = ~x5 & n277 ;
  assign n4577 = ( x2 & ~n155 ) | ( x2 & n4576 ) | ( ~n155 & n4576 ) ;
  assign n4578 = ~x2 & n4577 ;
  assign n4579 = ~n4575 & n4578 ;
  assign n4580 = x19 | x36 ;
  assign n4581 = ( n4575 & n4579 ) | ( n4575 & ~n4580 ) | ( n4579 & ~n4580 ) ;
  assign n4582 = ( x15 & n84 ) | ( x15 & n4581 ) | ( n84 & n4581 ) ;
  assign n4583 = ~x15 & n4582 ;
  assign n4584 = ( x13 & n383 ) | ( x13 & n4583 ) | ( n383 & n4583 ) ;
  assign n4585 = ~x13 & n4584 ;
  assign n4586 = ~x10 & n4585 ;
  assign n4587 = ( x9 & ~x11 ) | ( x9 & n4586 ) | ( ~x11 & n4586 ) ;
  assign n4588 = ~x9 & n4587 ;
  assign n4589 = ~x1 & n4588 ;
  assign n4590 = ( x0 & ~x8 ) | ( x0 & n4589 ) | ( ~x8 & n4589 ) ;
  assign n4591 = ~x0 & n4590 ;
  assign n4592 = ~x14 & n954 ;
  assign n4593 = ~x15 & n4592 ;
  assign n4594 = ( x15 & ~n304 ) | ( x15 & n4593 ) | ( ~n304 & n4593 ) ;
  assign n4595 = ( x13 & ~n487 ) | ( x13 & n4594 ) | ( ~n487 & n4594 ) ;
  assign n4596 = n4594 & ~n4595 ;
  assign n4597 = ( ~x0 & x4 ) | ( ~x0 & n4596 ) | ( x4 & n4596 ) ;
  assign n4598 = ( x14 & n570 ) | ( x14 & n2687 ) | ( n570 & n2687 ) ;
  assign n4599 = ~x14 & n4598 ;
  assign n4600 = ( x13 & x40 ) | ( x13 & n4599 ) | ( x40 & n4599 ) ;
  assign n4601 = x14 | x19 ;
  assign n4602 = x17 & n4601 ;
  assign n4603 = ( n1161 & n2869 ) | ( n1161 & ~n4602 ) | ( n2869 & ~n4602 ) ;
  assign n4604 = x15 & n4603 ;
  assign n4605 = x40 & n4604 ;
  assign n4606 = ( ~x13 & n4600 ) | ( ~x13 & n4605 ) | ( n4600 & n4605 ) ;
  assign n4607 = x5 | n4606 ;
  assign n4608 = ( x14 & n570 ) | ( x14 & n870 ) | ( n570 & n870 ) ;
  assign n4609 = ~x14 & n4608 ;
  assign n4610 = ~x13 & n4609 ;
  assign n4611 = x5 & ~n4610 ;
  assign n4612 = n4607 & ~n4611 ;
  assign n4613 = x4 | n4612 ;
  assign n4614 = ( x14 & n568 ) | ( x14 & n570 ) | ( n568 & n570 ) ;
  assign n4615 = ~x14 & n4614 ;
  assign n4616 = ~x13 & n4615 ;
  assign n4617 = x4 & ~n4616 ;
  assign n4618 = n4613 & ~n4617 ;
  assign n4619 = ( x16 & ~x18 ) | ( x16 & n4618 ) | ( ~x18 & n4618 ) ;
  assign n4620 = n129 | n3289 ;
  assign n4621 = ( n1417 & ~n4350 ) | ( n1417 & n4620 ) | ( ~n4350 & n4620 ) ;
  assign n4622 = n1417 & ~n4621 ;
  assign n4623 = ~x16 & n4622 ;
  assign n4624 = ( n4618 & ~n4619 ) | ( n4618 & n4623 ) | ( ~n4619 & n4623 ) ;
  assign n4625 = ~x0 & n4624 ;
  assign n4626 = ( ~x4 & n4597 ) | ( ~x4 & n4625 ) | ( n4597 & n4625 ) ;
  assign n4627 = x0 & ~x5 ;
  assign n4628 = ( x4 & ~n3289 ) | ( x4 & n4627 ) | ( ~n3289 & n4627 ) ;
  assign n4629 = ~x4 & n4628 ;
  assign n4630 = n4626 | n4629 ;
  assign n4631 = ( n156 & n4626 ) | ( n156 & n4630 ) | ( n4626 & n4630 ) ;
  assign n4632 = ( x36 & ~n198 ) | ( x36 & n4631 ) | ( ~n198 & n4631 ) ;
  assign n4633 = n4631 & ~n4632 ;
  assign n4634 = ~x9 & n4633 ;
  assign n4635 = ( x8 & ~x10 ) | ( x8 & n4634 ) | ( ~x10 & n4634 ) ;
  assign n4636 = ~x8 & n4635 ;
  assign n4637 = ~x2 & n4636 ;
  assign n4638 = ( x1 & ~x3 ) | ( x1 & n4637 ) | ( ~x3 & n4637 ) ;
  assign n4639 = ~x1 & n4638 ;
  assign n4640 = x14 | x16 ;
  assign n4641 = ( x16 & x17 ) | ( x16 & n51 ) | ( x17 & n51 ) ;
  assign n4642 = ( x14 & x16 ) | ( x14 & n4641 ) | ( x16 & n4641 ) ;
  assign n4643 = ( n4640 & n4641 ) | ( n4640 & ~n4642 ) | ( n4641 & ~n4642 ) ;
  assign n4644 = ( x15 & n196 ) | ( x15 & n4643 ) | ( n196 & n4643 ) ;
  assign n4645 = ~n4643 & n4644 ;
  assign n4646 = x13 & n4645 ;
  assign n4647 = ( x11 & x12 ) | ( x11 & n4646 ) | ( x12 & n4646 ) ;
  assign n4648 = ~x11 & n4647 ;
  assign n4649 = ~x9 & n4648 ;
  assign n4650 = ( x8 & ~x10 ) | ( x8 & n4649 ) | ( ~x10 & n4649 ) ;
  assign n4651 = ~x8 & n4650 ;
  assign n4652 = ~x4 & n4651 ;
  assign n4653 = ( x3 & ~x5 ) | ( x3 & n4652 ) | ( ~x5 & n4652 ) ;
  assign n4654 = ~x3 & n4653 ;
  assign n4655 = ~x1 & n4654 ;
  assign n4656 = ( x0 & ~x2 ) | ( x0 & n4655 ) | ( ~x2 & n4655 ) ;
  assign n4657 = ~x0 & n4656 ;
  assign n4658 = ( ~x5 & x19 ) | ( ~x5 & n1121 ) | ( x19 & n1121 ) ;
  assign n4659 = x14 & n4119 ;
  assign n4660 = x13 & n4659 ;
  assign n4661 = ~x38 & n418 ;
  assign n4662 = x37 & n4661 ;
  assign n4663 = ( ~n76 & n4660 ) | ( ~n76 & n4662 ) | ( n4660 & n4662 ) ;
  assign n4664 = n3289 | n4663 ;
  assign n4665 = ( ~n3289 & n4660 ) | ( ~n3289 & n4664 ) | ( n4660 & n4664 ) ;
  assign n4666 = ( x5 & x19 ) | ( x5 & n4665 ) | ( x19 & n4665 ) ;
  assign n4667 = n4658 & n4666 ;
  assign n4668 = x14 & ~x16 ;
  assign n4669 = x14 & ~n890 ;
  assign n4670 = ( n635 & n4668 ) | ( n635 & ~n4669 ) | ( n4668 & ~n4669 ) ;
  assign n4671 = ( ~x5 & n4667 ) | ( ~x5 & n4670 ) | ( n4667 & n4670 ) ;
  assign n4672 = x13 & ~n4671 ;
  assign n4673 = ( x13 & n4667 ) | ( x13 & ~n4672 ) | ( n4667 & ~n4672 ) ;
  assign n4674 = ( x12 & x40 ) | ( x12 & ~n4673 ) | ( x40 & ~n4673 ) ;
  assign n4675 = x40 & n4380 ;
  assign n4676 = ( n4673 & n4674 ) | ( n4673 & n4675 ) | ( n4674 & n4675 ) ;
  assign n4677 = ( x3 & ~x36 ) | ( x3 & n4676 ) | ( ~x36 & n4676 ) ;
  assign n4678 = ~x36 & n4375 ;
  assign n4679 = ( ~x3 & n4677 ) | ( ~x3 & n4678 ) | ( n4677 & n4678 ) ;
  assign n4680 = ~x10 & n4679 ;
  assign n4681 = ( x9 & ~x11 ) | ( x9 & n4680 ) | ( ~x11 & n4680 ) ;
  assign n4682 = ~x9 & n4681 ;
  assign n4683 = ~x4 & n4682 ;
  assign n4684 = ( x2 & ~x8 ) | ( x2 & n4683 ) | ( ~x8 & n4683 ) ;
  assign n4685 = ~x2 & n4684 ;
  assign n4686 = ~x0 & n4685 ;
  assign n4687 = ~x1 & n4686 ;
  assign n4688 = ~n159 & n2745 ;
  assign n4689 = n66 & n4688 ;
  assign n4690 = ( x19 & ~n731 ) | ( x19 & n2745 ) | ( ~n731 & n2745 ) ;
  assign n4691 = ( x18 & ~n153 ) | ( x18 & n1334 ) | ( ~n153 & n1334 ) ;
  assign n4692 = n1334 & ~n4691 ;
  assign n4693 = ~x19 & n4692 ;
  assign n4694 = ( n2745 & ~n4690 ) | ( n2745 & n4693 ) | ( ~n4690 & n4693 ) ;
  assign n4695 = x39 & n418 ;
  assign n4696 = ( x19 & ~n1734 ) | ( x19 & n4695 ) | ( ~n1734 & n4695 ) ;
  assign n4697 = n1734 & n4696 ;
  assign n4698 = ( ~n4689 & n4694 ) | ( ~n4689 & n4697 ) | ( n4694 & n4697 ) ;
  assign n4699 = n693 | n4697 ;
  assign n4700 = ( n4689 & n4698 ) | ( n4689 & n4699 ) | ( n4698 & n4699 ) ;
  assign n4701 = ( x14 & ~x36 ) | ( x14 & n4700 ) | ( ~x36 & n4700 ) ;
  assign n4702 = x36 | x40 ;
  assign n4703 = ( x14 & ~n4701 ) | ( x14 & n4702 ) | ( ~n4701 & n4702 ) ;
  assign n4704 = x4 | n4703 ;
  assign n4705 = ( ~x3 & x5 ) | ( ~x3 & n4704 ) | ( x5 & n4704 ) ;
  assign n4706 = x3 | n4705 ;
  assign n4707 = x1 | n4706 ;
  assign n4708 = ( ~x0 & x2 ) | ( ~x0 & n4707 ) | ( x2 & n4707 ) ;
  assign n4709 = x0 | n4708 ;
  assign n4710 = ~x36 & n4709 ;
  assign n4711 = x9 & x10 ;
  assign n4712 = ( x10 & n2823 ) | ( x10 & ~n4711 ) | ( n2823 & ~n4711 ) ;
  assign n4713 = ( n4710 & ~n4711 ) | ( n4710 & n4712 ) | ( ~n4711 & n4712 ) ;
  assign n4714 = x11 | n4713 ;
  assign n4715 = x8 | n4714 ;
  assign y0 = n184 ;
  assign y1 = 1'b0 ;
  assign y2 = n208 ;
  assign y3 = n229 ;
  assign y4 = n395 ;
  assign y5 = n468 ;
  assign y6 = n544 ;
  assign y7 = n687 ;
  assign y8 = n729 ;
  assign y9 = n759 ;
  assign y10 = n784 ;
  assign y11 = n856 ;
  assign y12 = n868 ;
  assign y13 = n916 ;
  assign y14 = n1102 ;
  assign y15 = n1187 ;
  assign y16 = ~n1435 ;
  assign y17 = n1471 ;
  assign y18 = n1520 ;
  assign y19 = n1598 ;
  assign y20 = n1789 ;
  assign y21 = n1806 ;
  assign y22 = ~n2013 ;
  assign y23 = n2038 ;
  assign y24 = ~n2319 ;
  assign y25 = n2448 ;
  assign y26 = n2597 ;
  assign y27 = ~n2822 ;
  assign y28 = n2845 ;
  assign y29 = ~n2941 ;
  assign y30 = n2957 ;
  assign y31 = 1'b0 ;
  assign y32 = 1'b0 ;
  assign y33 = n2966 ;
  assign y34 = ~n2986 ;
  assign y35 = n2990 ;
  assign y36 = n3009 ;
  assign y37 = ~n3067 ;
  assign y38 = ~n3098 ;
  assign y39 = 1'b0 ;
  assign y40 = n3118 ;
  assign y41 = n3216 ;
  assign y42 = n3288 ;
  assign y43 = n3376 ;
  assign y44 = n3453 ;
  assign y45 = n3535 ;
  assign y46 = n3619 ;
  assign y47 = n3731 ;
  assign y48 = n3823 ;
  assign y49 = n3865 ;
  assign y50 = n3945 ;
  assign y51 = n4034 ;
  assign y52 = n4106 ;
  assign y53 = n4162 ;
  assign y54 = n4207 ;
  assign y55 = n4224 ;
  assign y56 = n4247 ;
  assign y57 = n4278 ;
  assign y58 = n4298 ;
  assign y59 = n4312 ;
  assign y60 = n4328 ;
  assign y61 = n4336 ;
  assign y62 = n4404 ;
  assign y63 = n4429 ;
  assign y64 = n4445 ;
  assign y65 = n4485 ;
  assign y66 = n4544 ;
  assign y67 = n4591 ;
  assign y68 = n4639 ;
  assign y69 = n4657 ;
  assign y70 = n4687 ;
  assign y71 = n1114 ;
  assign y72 = ~n4715 ;
endmodule
