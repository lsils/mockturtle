module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246;
  assign n65 = x32 ^ x0;
  assign n67 = x33 ^ x1;
  assign n66 = x0 & x32;
  assign n68 = n67 ^ n66;
  assign n69 = n66 ^ x33;
  assign n70 = n67 & ~n69;
  assign n71 = n70 ^ x1;
  assign n72 = n71 ^ x2;
  assign n73 = n72 ^ x34;
  assign n74 = x34 ^ x2;
  assign n75 = n71 ^ x34;
  assign n76 = n74 & ~n75;
  assign n77 = n76 ^ x2;
  assign n78 = n77 ^ x3;
  assign n79 = n78 ^ x35;
  assign n80 = x35 ^ x3;
  assign n81 = n77 ^ x35;
  assign n82 = n80 & ~n81;
  assign n83 = n82 ^ x3;
  assign n84 = n83 ^ x4;
  assign n85 = n84 ^ x36;
  assign n86 = x36 ^ x4;
  assign n87 = n83 ^ x36;
  assign n88 = n86 & ~n87;
  assign n89 = n88 ^ x4;
  assign n90 = n89 ^ x5;
  assign n91 = n90 ^ x37;
  assign n92 = x37 ^ x5;
  assign n93 = n89 ^ x37;
  assign n94 = n92 & ~n93;
  assign n95 = n94 ^ x5;
  assign n96 = n95 ^ x6;
  assign n97 = n96 ^ x38;
  assign n98 = x38 ^ x6;
  assign n99 = n95 ^ x38;
  assign n100 = n98 & ~n99;
  assign n101 = n100 ^ x6;
  assign n102 = n101 ^ x7;
  assign n103 = n102 ^ x39;
  assign n104 = x39 ^ x7;
  assign n105 = n101 ^ x39;
  assign n106 = n104 & ~n105;
  assign n107 = n106 ^ x7;
  assign n108 = n107 ^ x8;
  assign n109 = n108 ^ x40;
  assign n110 = x40 ^ x8;
  assign n111 = n107 ^ x40;
  assign n112 = n110 & ~n111;
  assign n113 = n112 ^ x8;
  assign n114 = n113 ^ x9;
  assign n115 = n114 ^ x41;
  assign n116 = x41 ^ x9;
  assign n117 = n113 ^ x41;
  assign n118 = n116 & ~n117;
  assign n119 = n118 ^ x9;
  assign n120 = n119 ^ x10;
  assign n121 = n120 ^ x42;
  assign n122 = x42 ^ x10;
  assign n123 = n119 ^ x42;
  assign n124 = n122 & ~n123;
  assign n125 = n124 ^ x10;
  assign n126 = n125 ^ x11;
  assign n127 = n126 ^ x43;
  assign n128 = x43 ^ x11;
  assign n129 = n125 ^ x43;
  assign n130 = n128 & ~n129;
  assign n131 = n130 ^ x11;
  assign n132 = n131 ^ x12;
  assign n133 = n132 ^ x44;
  assign n134 = x44 ^ x12;
  assign n135 = n131 ^ x44;
  assign n136 = n134 & ~n135;
  assign n137 = n136 ^ x12;
  assign n138 = n137 ^ x13;
  assign n139 = n138 ^ x45;
  assign n140 = x45 ^ x13;
  assign n141 = n137 ^ x45;
  assign n142 = n140 & ~n141;
  assign n143 = n142 ^ x13;
  assign n144 = n143 ^ x14;
  assign n145 = n144 ^ x46;
  assign n146 = x46 ^ x14;
  assign n147 = n143 ^ x46;
  assign n148 = n146 & ~n147;
  assign n149 = n148 ^ x14;
  assign n150 = n149 ^ x15;
  assign n151 = n150 ^ x47;
  assign n152 = x47 ^ x15;
  assign n153 = n149 ^ x47;
  assign n154 = n152 & ~n153;
  assign n155 = n154 ^ x15;
  assign n156 = n155 ^ x48;
  assign n157 = n156 ^ x16;
  assign n158 = x48 ^ x16;
  assign n159 = ~n156 & n158;
  assign n160 = n159 ^ x16;
  assign n161 = n160 ^ x17;
  assign n162 = n161 ^ x49;
  assign n163 = x49 ^ x17;
  assign n164 = n160 ^ x49;
  assign n165 = n163 & ~n164;
  assign n166 = n165 ^ x17;
  assign n167 = n166 ^ x18;
  assign n168 = n167 ^ x50;
  assign n169 = x50 ^ x18;
  assign n170 = n166 ^ x50;
  assign n171 = n169 & ~n170;
  assign n172 = n171 ^ x18;
  assign n173 = n172 ^ x19;
  assign n174 = n173 ^ x51;
  assign n175 = x51 ^ x19;
  assign n176 = n172 ^ x51;
  assign n177 = n175 & ~n176;
  assign n178 = n177 ^ x19;
  assign n179 = n178 ^ x20;
  assign n180 = n179 ^ x52;
  assign n181 = x52 ^ x20;
  assign n182 = n178 ^ x52;
  assign n183 = n181 & ~n182;
  assign n184 = n183 ^ x20;
  assign n185 = n184 ^ x53;
  assign n186 = n185 ^ x21;
  assign n187 = x53 ^ x21;
  assign n188 = ~n185 & n187;
  assign n189 = n188 ^ x21;
  assign n190 = n189 ^ x22;
  assign n191 = n190 ^ x54;
  assign n192 = x54 ^ x22;
  assign n193 = n189 ^ x54;
  assign n194 = n192 & ~n193;
  assign n195 = n194 ^ x22;
  assign n196 = n195 ^ x23;
  assign n197 = n196 ^ x55;
  assign n198 = x55 ^ x23;
  assign n199 = n195 ^ x55;
  assign n200 = n198 & ~n199;
  assign n201 = n200 ^ x23;
  assign n202 = n201 ^ x24;
  assign n203 = n202 ^ x56;
  assign n204 = x56 ^ x24;
  assign n205 = n201 ^ x56;
  assign n206 = n204 & ~n205;
  assign n207 = n206 ^ x24;
  assign n208 = n207 ^ x25;
  assign n209 = n208 ^ x57;
  assign n210 = x57 ^ x25;
  assign n211 = n207 ^ x57;
  assign n212 = n210 & ~n211;
  assign n213 = n212 ^ x25;
  assign n214 = n213 ^ x26;
  assign n215 = n214 ^ x58;
  assign n216 = x58 ^ x26;
  assign n217 = n213 ^ x58;
  assign n218 = n216 & ~n217;
  assign n219 = n218 ^ x26;
  assign n220 = n219 ^ x59;
  assign n221 = n220 ^ x27;
  assign n222 = x59 ^ x27;
  assign n223 = ~n220 & n222;
  assign n224 = n223 ^ x27;
  assign n225 = n224 ^ x28;
  assign n226 = n225 ^ x60;
  assign n227 = x60 ^ x28;
  assign n228 = n224 ^ x60;
  assign n229 = n227 & ~n228;
  assign n230 = n229 ^ x28;
  assign n231 = n230 ^ x61;
  assign n232 = n231 ^ x29;
  assign n233 = x61 ^ x29;
  assign n234 = ~n231 & n233;
  assign n235 = n234 ^ x29;
  assign n236 = n235 ^ x30;
  assign n237 = n236 ^ x62;
  assign n242 = x63 ^ x31;
  assign n238 = x62 ^ x30;
  assign n239 = n235 ^ x62;
  assign n240 = n238 & ~n239;
  assign n241 = n240 ^ x30;
  assign n243 = n242 ^ n241;
  assign n244 = n241 ^ x63;
  assign n245 = n242 & ~n244;
  assign n246 = n245 ^ x31;
  assign y0 = n65;
  assign y1 = n68;
  assign y2 = n73;
  assign y3 = n79;
  assign y4 = n85;
  assign y5 = n91;
  assign y6 = n97;
  assign y7 = n103;
  assign y8 = n109;
  assign y9 = n115;
  assign y10 = n121;
  assign y11 = n127;
  assign y12 = n133;
  assign y13 = n139;
  assign y14 = n145;
  assign y15 = n151;
  assign y16 = n157;
  assign y17 = n162;
  assign y18 = n168;
  assign y19 = n174;
  assign y20 = n180;
  assign y21 = n186;
  assign y22 = n191;
  assign y23 = n197;
  assign y24 = n203;
  assign y25 = n209;
  assign y26 = n215;
  assign y27 = n221;
  assign y28 = n226;
  assign y29 = n232;
  assign y30 = n237;
  assign y31 = n243;
  assign y32 = n246;
endmodule
