module top( G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 , G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 );
  input G1 , G10 , G100 , G101 , G102 , G103 , G104 , G105 , G106 , G107 , G108 , G109 , G11 , G110 , G111 , G112 , G113 , G114 , G115 , G116 , G117 , G118 , G119 , G12 , G120 , G121 , G122 , G123 , G124 , G125 , G126 , G127 , G128 , G129 , G13 , G130 , G131 , G132 , G133 , G134 , G135 , G136 , G137 , G138 , G139 , G14 , G140 , G141 , G142 , G143 , G144 , G145 , G146 , G147 , G148 , G149 , G15 , G150 , G151 , G152 , G153 , G154 , G155 , G156 , G157 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G42 , G43 , G44 , G45 , G46 , G47 , G48 , G49 , G5 , G50 , G51 , G52 , G53 , G54 , G55 , G56 , G57 , G58 , G59 , G6 , G60 , G61 , G62 , G63 , G64 , G65 , G66 , G67 , G68 , G69 , G7 , G70 , G71 , G72 , G73 , G74 , G75 , G76 , G77 , G78 , G79 , G8 , G80 , G81 , G82 , G83 , G84 , G85 , G86 , G87 , G88 , G89 , G9 , G90 , G91 , G92 , G93 , G94 , G95 , G96 , G97 , G98 , G99 ;
  output G2531 , G2532 , G2533 , G2534 , G2535 , G2536 , G2537 , G2538 , G2539 , G2540 , G2541 , G2542 , G2543 , G2544 , G2545 , G2546 , G2547 , G2548 , G2549 , G2550 , G2551 , G2552 , G2553 , G2554 , G2555 , G2556 , G2557 , G2558 , G2559 , G2560 , G2561 , G2562 , G2563 , G2564 , G2565 , G2566 , G2567 , G2568 , G2569 , G2570 , G2571 , G2572 , G2573 , G2574 , G2575 , G2576 , G2577 , G2578 , G2579 , G2580 , G2581 , G2582 , G2583 , G2584 , G2585 , G2586 , G2587 , G2588 , G2589 , G2590 , G2591 , G2592 , G2593 , G2594 ;
  wire n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 ;
  assign n158 = G141 | G142 ;
  assign n159 = G139 | G140 ;
  assign n160 = n158 | n159 ;
  assign n161 = G121 | G2 ;
  assign n162 = G11 | n161 ;
  assign n163 = G115 & ~G74 ;
  assign n164 = G121 | G7 ;
  assign n165 = G119 | n164 ;
  assign n166 = G147 | n164 ;
  assign n167 = G53 & ~G96 ;
  assign n168 = G43 | G86 ;
  assign n169 = n167 & ~n168 ;
  assign n170 = ~G106 & G32 ;
  assign n171 = G64 | G76 ;
  assign n172 = n170 & ~n171 ;
  assign n173 = n169 | n172 ;
  assign n174 = G147 & ~n172 ;
  assign n175 = G119 & ~n169 ;
  assign n176 = n174 | n175 ;
  assign n177 = G145 | G146 ;
  assign n178 = G109 & ~n177 ;
  assign n179 = G79 & ~n177 ;
  assign n180 = n178 | n179 ;
  assign n181 = G89 & ~n177 ;
  assign n182 = G99 & ~n177 ;
  assign n183 = n181 | n182 ;
  assign n184 = n180 | n183 ;
  assign n185 = G108 | n177 ;
  assign n186 = G98 & ~n177 ;
  assign n187 = n185 & ~n186 ;
  assign n188 = G88 & ~n177 ;
  assign n189 = G78 & ~n177 ;
  assign n190 = n188 | n189 ;
  assign n191 = n187 & ~n190 ;
  assign n192 = G80 | n177 ;
  assign n193 = G90 & ~n177 ;
  assign n194 = n192 & ~n193 ;
  assign n195 = G100 & ~n177 ;
  assign n196 = G110 & ~n177 ;
  assign n197 = n195 | n196 ;
  assign n198 = n194 & ~n197 ;
  assign n199 = G117 & ~G36 ;
  assign n200 = G117 & ~G68 ;
  assign n201 = G120 | n200 ;
  assign n202 = n199 & ~n201 ;
  assign n203 = G117 | G120 ;
  assign n204 = G46 & ~n203 ;
  assign n205 = G57 & ~n203 ;
  assign n206 = n204 | n205 ;
  assign n207 = n202 & ~n206 ;
  assign n208 = G117 & ~G37 ;
  assign n209 = G117 & ~G69 ;
  assign n210 = G120 | n209 ;
  assign n211 = n208 & ~n210 ;
  assign n212 = G47 & ~n203 ;
  assign n213 = G58 & ~n203 ;
  assign n214 = n212 | n213 ;
  assign n215 = n211 & ~n214 ;
  assign n216 = G117 & ~G38 ;
  assign n217 = G117 & ~G70 ;
  assign n218 = G120 | n217 ;
  assign n219 = n216 & ~n218 ;
  assign n220 = G48 & ~n203 ;
  assign n221 = G59 & ~n203 ;
  assign n222 = n220 | n221 ;
  assign n223 = n219 & ~n222 ;
  assign n224 = G117 & ~G31 ;
  assign n225 = G117 & ~G63 ;
  assign n226 = G120 | n225 ;
  assign n227 = n224 & ~n226 ;
  assign n228 = G42 & ~n203 ;
  assign n229 = G52 & ~n203 ;
  assign n230 = n228 | n229 ;
  assign n231 = n227 & ~n230 ;
  assign n232 = G122 | n231 ;
  assign n233 = G116 | G121 ;
  assign n234 = n176 | n233 ;
  assign n235 = G28 | n234 ;
  assign n236 = G1 & ~G3 ;
  assign n237 = n234 | n236 ;
  assign n238 = G117 | G39 ;
  assign n239 = G117 & ~G71 ;
  assign n240 = G120 | n239 ;
  assign n241 = n238 & ~n240 ;
  assign n242 = G49 & ~n203 ;
  assign n243 = G60 & ~n203 ;
  assign n244 = n242 | n243 ;
  assign n245 = n241 | n244 ;
  assign n246 = G56 & ~n203 ;
  assign n247 = G117 | G35 ;
  assign n248 = G117 & ~G67 ;
  assign n249 = G120 | n248 ;
  assign n250 = n247 & ~n249 ;
  assign n251 = n246 & ~n250 ;
  assign n252 = G117 & ~G34 ;
  assign n253 = G117 & ~G66 ;
  assign n254 = G120 | n253 ;
  assign n255 = n252 & ~n254 ;
  assign n256 = G45 & ~n203 ;
  assign n257 = G55 & ~n203 ;
  assign n258 = n256 | n257 ;
  assign n259 = n255 & ~n258 ;
  assign n260 = G117 & ~G33 ;
  assign n261 = G117 & ~G65 ;
  assign n262 = G120 | n261 ;
  assign n263 = n260 & ~n262 ;
  assign n264 = G44 & ~n203 ;
  assign n265 = G54 & ~n203 ;
  assign n266 = n264 | n265 ;
  assign n267 = n263 & ~n266 ;
  assign n268 = G117 & ~G40 ;
  assign n269 = G117 & ~G72 ;
  assign n270 = G120 | n269 ;
  assign n271 = n268 & ~n270 ;
  assign n272 = G50 & ~n203 ;
  assign n273 = G61 & ~n203 ;
  assign n274 = n272 | n273 ;
  assign n275 = n271 & ~n274 ;
  assign n276 = G123 | n275 ;
  assign n277 = G123 & ~n223 ;
  assign n278 = n276 & ~n277 ;
  assign n279 = G123 | n245 ;
  assign n280 = ~G123 & n215 ;
  assign n281 = n279 & ~n280 ;
  assign n282 = G118 & ~G122 ;
  assign n283 = n275 | n282 ;
  assign n284 = G123 & ~n231 ;
  assign n285 = G118 | G123 ;
  assign n286 = n275 & ~n285 ;
  assign n287 = n284 | n286 ;
  assign n288 = G77 & ~n177 ;
  assign n289 = G97 & ~n177 ;
  assign n290 = n288 & ~n289 ;
  assign n291 = G107 & ~n177 ;
  assign n292 = G87 & ~n177 ;
  assign n293 = n291 | n292 ;
  assign n294 = n290 & ~n293 ;
  assign n295 = G143 | n294 ;
  assign n296 = G143 & ~n294 ;
  assign n297 = n295 & ~n296 ;
  assign n298 = G144 | n297 ;
  assign n299 = ~G19 & G23 ;
  assign n300 = G75 & ~n177 ;
  assign n301 = G85 & ~n177 ;
  assign n302 = n300 & ~n301 ;
  assign n303 = G95 & ~n177 ;
  assign n304 = G105 & ~n177 ;
  assign n305 = n303 | n304 ;
  assign n306 = n302 & ~n305 ;
  assign n307 = G23 & ~n306 ;
  assign n308 = n299 & ~n307 ;
  assign n309 = G135 & ~n308 ;
  assign n310 = G12 & ~G13 ;
  assign n311 = G12 & ~n231 ;
  assign n312 = n310 & ~n311 ;
  assign n313 = G125 & ~n312 ;
  assign n314 = G12 & ~G15 ;
  assign n315 = ~G12 & n215 ;
  assign n316 = n314 & ~n315 ;
  assign n317 = G130 & ~n316 ;
  assign n318 = n313 | n317 ;
  assign n319 = n309 | n318 ;
  assign n320 = G12 & ~G5 ;
  assign n321 = G12 & ~n223 ;
  assign n322 = n320 & ~n321 ;
  assign n323 = G129 & ~n322 ;
  assign n324 = ~G21 & G23 ;
  assign n325 = G23 & ~n198 ;
  assign n326 = n324 & ~n325 ;
  assign n327 = G140 & ~n326 ;
  assign n328 = n323 | n327 ;
  assign n329 = G23 & ~G27 ;
  assign n330 = G23 & ~n191 ;
  assign n331 = n329 & ~n330 ;
  assign n332 = G142 & ~n331 ;
  assign n333 = n309 | n332 ;
  assign n334 = n328 | n333 ;
  assign n335 = G12 & ~G14 ;
  assign n336 = ~G12 & n245 ;
  assign n337 = n335 & ~n336 ;
  assign n338 = G128 & ~n337 ;
  assign n339 = G12 & ~G4 ;
  assign n340 = G12 & ~n275 ;
  assign n341 = n339 & ~n340 ;
  assign n342 = G126 & ~n341 ;
  assign n343 = n338 | n342 ;
  assign n344 = G23 & ~G26 ;
  assign n345 = G23 & ~n184 ;
  assign n346 = n344 & ~n345 ;
  assign n347 = G141 & ~n346 ;
  assign n348 = n327 | n347 ;
  assign n349 = n343 | n348 ;
  assign n350 = n334 | n349 ;
  assign n351 = n319 | n350 ;
  assign n352 = G23 & ~G24 ;
  assign n353 = G93 & ~n177 ;
  assign n354 = G103 & ~n177 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = G113 & ~n177 ;
  assign n357 = G83 & ~n177 ;
  assign n358 = n356 | n357 ;
  assign n359 = n355 & ~n358 ;
  assign n360 = G23 & ~n359 ;
  assign n361 = n352 & ~n360 ;
  assign n362 = G136 | n361 ;
  assign n363 = G136 & ~n361 ;
  assign n364 = n362 & ~n363 ;
  assign n365 = G12 & ~G16 ;
  assign n366 = G12 & ~n207 ;
  assign n367 = n365 & ~n366 ;
  assign n368 = G131 | n367 ;
  assign n369 = G131 & ~n367 ;
  assign n370 = n368 & ~n369 ;
  assign n371 = ~G20 & G23 ;
  assign n372 = G82 & ~n177 ;
  assign n373 = G102 & ~n177 ;
  assign n374 = n372 & ~n373 ;
  assign n375 = G112 & ~n177 ;
  assign n376 = G92 & ~n177 ;
  assign n377 = n375 | n376 ;
  assign n378 = n374 & ~n377 ;
  assign n379 = G23 & ~n378 ;
  assign n380 = n371 & ~n379 ;
  assign n381 = G138 | n380 ;
  assign n382 = G138 & ~n380 ;
  assign n383 = n381 & ~n382 ;
  assign n384 = n370 | n383 ;
  assign n385 = n364 | n384 ;
  assign n386 = G23 & ~G25 ;
  assign n387 = G81 & ~n177 ;
  assign n388 = G101 & ~n177 ;
  assign n389 = n387 & ~n388 ;
  assign n390 = G111 & ~n177 ;
  assign n391 = G91 & ~n177 ;
  assign n392 = n390 | n391 ;
  assign n393 = n389 & ~n392 ;
  assign n394 = G23 & ~n393 ;
  assign n395 = n386 & ~n394 ;
  assign n396 = G139 & ~n395 ;
  assign n397 = n317 | n396 ;
  assign n398 = G12 & ~G18 ;
  assign n399 = G12 & ~n267 ;
  assign n400 = n398 & ~n399 ;
  assign n401 = G134 & ~n400 ;
  assign n402 = n342 | n401 ;
  assign n403 = n397 | n402 ;
  assign n404 = G12 & ~G6 ;
  assign n405 = G12 & ~n259 ;
  assign n406 = n404 & ~n405 ;
  assign n407 = G133 & ~n406 ;
  assign n408 = G23 & ~n294 ;
  assign n409 = ~G22 & G23 ;
  assign n410 = G9 | n409 ;
  assign n411 = n408 | n410 ;
  assign n412 = n407 | n411 ;
  assign n413 = n332 | n407 ;
  assign n414 = n412 | n413 ;
  assign n415 = n403 | n414 ;
  assign n416 = n323 | n347 ;
  assign n417 = n313 | n338 ;
  assign n418 = n416 | n417 ;
  assign n419 = n396 | n401 ;
  assign n420 = G12 & ~G17 ;
  assign n421 = G12 & ~n251 ;
  assign n422 = n420 & ~n421 ;
  assign n423 = G132 & ~n422 ;
  assign n424 = n419 | n423 ;
  assign n425 = n418 | n424 ;
  assign n426 = n415 | n425 ;
  assign n427 = n385 | n426 ;
  assign n428 = n351 | n427 ;
  assign n429 = G117 & ~G41 ;
  assign n430 = G117 & ~G73 ;
  assign n431 = G120 | n430 ;
  assign n432 = n429 & ~n431 ;
  assign n433 = G51 & ~n203 ;
  assign n434 = G62 & ~n203 ;
  assign n435 = n433 | n434 ;
  assign n436 = n432 & ~n435 ;
  assign n437 = G122 & ~n436 ;
  assign n438 = G122 | n437 ;
  assign n439 = n191 | n294 ;
  assign n440 = n191 & ~n294 ;
  assign n441 = n439 & ~n440 ;
  assign n442 = n184 | n441 ;
  assign n443 = ~n184 & n441 ;
  assign n444 = n442 & ~n443 ;
  assign n445 = G29 | n444 ;
  assign n446 = G123 & ~n436 ;
  assign n447 = G123 | n446 ;
  assign n448 = G127 | n198 ;
  assign n449 = G30 | n184 ;
  assign n450 = n448 | n449 ;
  assign n451 = ~G8 & n450 ;
  assign n452 = ~G133 & n451 ;
  assign n453 = G8 | n450 ;
  assign n454 = n259 | n453 ;
  assign n455 = ~G132 & n451 ;
  assign n456 = G129 & n450 ;
  assign n457 = G140 & ~n450 ;
  assign n458 = n456 & ~n457 ;
  assign n459 = n223 & ~n458 ;
  assign n460 = ~G128 & n450 ;
  assign n461 = G139 & ~n450 ;
  assign n462 = n460 | n461 ;
  assign n463 = ~n245 & n462 ;
  assign n464 = ~G126 & n450 ;
  assign n465 = G138 & ~n450 ;
  assign n466 = n464 | n465 ;
  assign n467 = n275 | n466 ;
  assign n468 = ~G125 & n450 ;
  assign n469 = G136 & ~n450 ;
  assign n470 = n468 | n469 ;
  assign n471 = ~n231 & n470 ;
  assign n472 = n467 & n471 ;
  assign n473 = n275 & n466 ;
  assign n474 = n245 & n462 ;
  assign n475 = n473 | n474 ;
  assign n476 = n472 | n475 ;
  assign n477 = ~n463 & n476 ;
  assign n478 = n459 | n477 ;
  assign n479 = G8 & ~n215 ;
  assign n480 = G130 & n451 ;
  assign n481 = G141 & ~n453 ;
  assign n482 = n480 & ~n481 ;
  assign n483 = n479 & ~n482 ;
  assign n484 = n459 | n483 ;
  assign n485 = n478 & ~n484 ;
  assign n486 = G8 & ~n207 ;
  assign n487 = G131 & n451 ;
  assign n488 = G142 & ~n453 ;
  assign n489 = n487 & ~n488 ;
  assign n490 = n486 & ~n489 ;
  assign n491 = n483 | n490 ;
  assign n492 = n485 | n491 ;
  assign n493 = n251 & ~n453 ;
  assign n494 = n490 | n493 ;
  assign n495 = n492 & ~n494 ;
  assign n496 = n455 | n495 ;
  assign n497 = n454 & n496 ;
  assign n498 = n452 | n497 ;
  assign n499 = n448 & ~n449 ;
  assign n500 = G136 | n359 ;
  assign n501 = n499 & ~n500 ;
  assign n502 = G138 | n378 ;
  assign n503 = n499 & ~n502 ;
  assign n504 = n501 & ~n503 ;
  assign n505 = G135 | n306 ;
  assign n506 = G134 & ~n267 ;
  assign n507 = n505 & ~n506 ;
  assign n508 = n499 & ~n507 ;
  assign n509 = n503 | n508 ;
  assign n510 = G135 & ~n306 ;
  assign n511 = n500 & ~n510 ;
  assign n512 = n499 & ~n511 ;
  assign n513 = G134 | n267 ;
  assign n514 = n499 & ~n513 ;
  assign n515 = n512 | n514 ;
  assign n516 = n509 | n515 ;
  assign n517 = n504 & ~n516 ;
  assign n518 = n498 & n517 ;
  assign n519 = n505 & ~n514 ;
  assign n520 = n512 & ~n519 ;
  assign n521 = n504 & ~n520 ;
  assign n522 = n503 | n521 ;
  assign n523 = n518 | n522 ;
  assign n524 = G10 & ~n176 ;
  assign n525 = n445 & n524 ;
  assign G2531 = G115 ;
  assign G2532 = G115 ;
  assign G2533 = G115 ;
  assign G2534 = G124 ;
  assign G2535 = G124 ;
  assign G2536 = G137 ;
  assign G2537 = G137 ;
  assign G2538 = G137 ;
  assign G2539 = G32 ;
  assign G2540 = G106 ;
  assign G2541 = G64 ;
  assign G2542 = G76 ;
  assign G2543 = G53 ;
  assign G2544 = G96 ;
  assign G2545 = G43 ;
  assign G2546 = G86 ;
  assign G2547 = n160 ;
  assign G2548 = n162 ;
  assign G2549 = G115 ;
  assign G2550 = n163 ;
  assign G2551 = n164 ;
  assign G2552 = n165 ;
  assign G2553 = n166 ;
  assign G2554 = n173 ;
  assign G2555 = n173 ;
  assign G2556 = n176 ;
  assign G2557 = n184 ;
  assign G2558 = n191 ;
  assign G2559 = n198 ;
  assign G2560 = n207 ;
  assign G2561 = n215 ;
  assign G2562 = n223 ;
  assign G2563 = n232 ;
  assign G2564 = n235 ;
  assign G2565 = n237 ;
  assign G2566 = n245 ;
  assign G2567 = n223 ;
  assign G2568 = n215 ;
  assign G2569 = n207 ;
  assign G2570 = n251 ;
  assign G2571 = n259 ;
  assign G2572 = n267 ;
  assign G2573 = n278 ;
  assign G2574 = n278 ;
  assign G2575 = n281 ;
  assign G2576 = n281 ;
  assign G2577 = n283 ;
  assign G2578 = n287 ;
  assign G2579 = n287 ;
  assign G2580 = n298 ;
  assign G2581 = ~G10 ;
  assign G2582 = 1'b0 ;
  assign G2583 = 1'b0 ;
  assign G2584 = n428 ;
  assign G2585 = n428 ;
  assign G2586 = n438 ;
  assign G2587 = ~n445 ;
  assign G2588 = n447 ;
  assign G2589 = n447 ;
  assign G2590 = 1'b0 ;
  assign G2591 = ~n523 ;
  assign G2592 = 1'b0 ;
  assign G2593 = ~n525 ;
  assign G2594 = ~n525 ;
endmodule
