module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 ;
  assign n67 = ~x9 & x11 ;
  assign n68 = x10 | n67 ;
  assign n32 = ~x12 & x13 ;
  assign n69 = x8 & x11 ;
  assign n70 = x9 & n69 ;
  assign n71 = x10 & ~n70 ;
  assign n72 = x9 | x10 ;
  assign n73 = ( ~x10 & n71 ) | ( ~x10 & n72 ) | ( n71 & n72 ) ;
  assign n86 = x3 & x5 ;
  assign n88 = ( x2 & n73 ) | ( x2 & n86 ) | ( n73 & n86 ) ;
  assign n87 = x4 & ~x5 ;
  assign n89 = ( ~x2 & n73 ) | ( ~x2 & n87 ) | ( n73 & n87 ) ;
  assign n90 = n88 & n89 ;
  assign n77 = x2 & ~x5 ;
  assign n78 = ( x2 & x4 ) | ( x2 & x5 ) | ( x4 & x5 ) ;
  assign n79 = ( x6 & n77 ) | ( x6 & n78 ) | ( n77 & n78 ) ;
  assign n83 = ( x3 & ~n73 ) | ( x3 & n79 ) | ( ~n73 & n79 ) ;
  assign n80 = x3 | x6 ;
  assign n81 = ~x4 & x5 ;
  assign n82 = ( x3 & ~n80 ) | ( x3 & n81 ) | ( ~n80 & n81 ) ;
  assign n84 = n73 & n82 ;
  assign n85 = ( n79 & ~n83 ) | ( n79 & n84 ) | ( ~n83 & n84 ) ;
  assign n91 = n85 & ~n90 ;
  assign n92 = ( n32 & n90 ) | ( n32 & n91 ) | ( n90 & n91 ) ;
  assign n122 = ( x1 & x7 ) | ( x1 & ~n92 ) | ( x7 & ~n92 ) ;
  assign n93 = ~x8 & x11 ;
  assign n94 = x9 | x11 ;
  assign n95 = ( ~x11 & n93 ) | ( ~x11 & n94 ) | ( n93 & n94 ) ;
  assign n96 = ( x8 & x10 ) | ( x8 & ~x11 ) | ( x10 & ~x11 ) ;
  assign n97 = x9 & ~n96 ;
  assign n98 = ( ~x8 & x9 ) | ( ~x8 & x11 ) | ( x9 & x11 ) ;
  assign n99 = x10 & ~n98 ;
  assign n100 = ( ~x7 & x8 ) | ( ~x7 & n99 ) | ( x8 & n99 ) ;
  assign n101 = x11 & ~n100 ;
  assign n102 = ( x11 & n99 ) | ( x11 & ~n101 ) | ( n99 & ~n101 ) ;
  assign n103 = n97 | n102 ;
  assign n104 = x7 | n103 ;
  assign n105 = ( n95 & n103 ) | ( n95 & n104 ) | ( n103 & n104 ) ;
  assign n106 = x7 & ~x11 ;
  assign n107 = x10 & n106 ;
  assign n108 = x6 | n107 ;
  assign n109 = ( n105 & n107 ) | ( n105 & n108 ) | ( n107 & n108 ) ;
  assign n115 = x0 | x4 ;
  assign n110 = x3 | x5 ;
  assign n116 = ( x0 & ~x4 ) | ( x0 & n110 ) | ( ~x4 & n110 ) ;
  assign n15 = x3 & ~x4 ;
  assign n111 = x2 | x5 ;
  assign n112 = x3 | x4 ;
  assign n113 = ( ~x3 & n15 ) | ( ~x3 & n112 ) | ( n15 & n112 ) ;
  assign n114 = ( n15 & n111 ) | ( n15 & n113 ) | ( n111 & n113 ) ;
  assign n117 = x0 & n114 ;
  assign n118 = ( n115 & ~n116 ) | ( n115 & n117 ) | ( ~n116 & n117 ) ;
  assign n119 = x12 & n118 ;
  assign n120 = ( x13 & n109 ) | ( x13 & ~n119 ) | ( n109 & ~n119 ) ;
  assign n121 = n109 & ~n120 ;
  assign n123 = x1 & n121 ;
  assign n124 = ( n92 & n122 ) | ( n92 & n123 ) | ( n122 & n123 ) ;
  assign n16 = ( x3 & x5 ) | ( x3 & n15 ) | ( x5 & n15 ) ;
  assign n17 = ( ~x3 & x5 ) | ( ~x3 & n15 ) | ( x5 & n15 ) ;
  assign n18 = ( x3 & ~n16 ) | ( x3 & n17 ) | ( ~n16 & n17 ) ;
  assign n74 = ~x13 & n18 ;
  assign n75 = ( x12 & n73 ) | ( x12 & ~n74 ) | ( n73 & ~n74 ) ;
  assign n76 = n73 & ~n75 ;
  assign n125 = ( x2 & n76 ) | ( x2 & n124 ) | ( n76 & n124 ) ;
  assign n126 = x7 & ~n125 ;
  assign n127 = ( x7 & n124 ) | ( x7 & ~n126 ) | ( n124 & ~n126 ) ;
  assign n19 = x8 & ~x12 ;
  assign n20 = ( x13 & n18 ) | ( x13 & ~n19 ) | ( n18 & ~n19 ) ;
  assign n21 = n18 & ~n20 ;
  assign n22 = ( ~x3 & x4 ) | ( ~x3 & x6 ) | ( x4 & x6 ) ;
  assign n23 = ~x4 & n22 ;
  assign n24 = ( ~x5 & n22 ) | ( ~x5 & n23 ) | ( n22 & n23 ) ;
  assign n25 = x3 & ~n15 ;
  assign n26 = x2 & n25 ;
  assign n27 = ( x4 & n15 ) | ( x4 & ~n26 ) | ( n15 & ~n26 ) ;
  assign n28 = ( x6 & n15 ) | ( x6 & n27 ) | ( n15 & n27 ) ;
  assign n29 = x5 & n28 ;
  assign n30 = x2 | n29 ;
  assign n31 = ( n24 & n29 ) | ( n24 & n30 ) | ( n29 & n30 ) ;
  assign n33 = ( x8 & ~n31 ) | ( x8 & n32 ) | ( ~n31 & n32 ) ;
  assign n34 = n31 & n33 ;
  assign n61 = ( x1 & x7 ) | ( x1 & n34 ) | ( x7 & n34 ) ;
  assign n37 = x0 & x3 ;
  assign n38 = x7 & ~x13 ;
  assign n39 = ( x12 & n37 ) | ( x12 & n38 ) | ( n37 & n38 ) ;
  assign n40 = ~n37 & n39 ;
  assign n35 = x8 & n32 ;
  assign n36 = x5 | x7 ;
  assign n41 = ( n35 & ~n36 ) | ( n35 & n40 ) | ( ~n36 & n40 ) ;
  assign n42 = x2 & ~n41 ;
  assign n43 = ( x2 & n40 ) | ( x2 & ~n42 ) | ( n40 & ~n42 ) ;
  assign n58 = ( ~x4 & x6 ) | ( ~x4 & n43 ) | ( x6 & n43 ) ;
  assign n44 = x12 & n38 ;
  assign n45 = ~x4 & n44 ;
  assign n46 = x0 & n45 ;
  assign n47 = ( x5 & ~x7 ) | ( x5 & n46 ) | ( ~x7 & n46 ) ;
  assign n48 = n35 & ~n47 ;
  assign n49 = ( n35 & n46 ) | ( n35 & ~n48 ) | ( n46 & ~n48 ) ;
  assign n50 = ~x2 & n49 ;
  assign n51 = n45 | n50 ;
  assign n52 = ( x0 & n50 ) | ( x0 & n51 ) | ( n50 & n51 ) ;
  assign n53 = ~x7 & n35 ;
  assign n54 = ( x4 & x5 ) | ( x4 & n53 ) | ( x5 & n53 ) ;
  assign n55 = ~x4 & n54 ;
  assign n56 = x3 | n55 ;
  assign n57 = ( n52 & n55 ) | ( n52 & n56 ) | ( n55 & n56 ) ;
  assign n59 = ~x6 & n57 ;
  assign n60 = ( n43 & ~n58 ) | ( n43 & n59 ) | ( ~n58 & n59 ) ;
  assign n62 = x1 & n60 ;
  assign n63 = ( ~x7 & n61 ) | ( ~x7 & n62 ) | ( n61 & n62 ) ;
  assign n64 = ( x2 & ~x7 ) | ( x2 & n63 ) | ( ~x7 & n63 ) ;
  assign n65 = n21 & ~n64 ;
  assign n66 = ( n21 & n63 ) | ( n21 & ~n65 ) | ( n63 & ~n65 ) ;
  assign n128 = n66 | n127 ;
  assign n129 = ( n68 & n127 ) | ( n68 & n128 ) | ( n127 & n128 ) ;
  assign n130 = x3 & x4 ;
  assign n131 = n81 & ~n130 ;
  assign n132 = x12 & ~x13 ;
  assign n133 = ( n130 & n131 ) | ( n130 & n132 ) | ( n131 & n132 ) ;
  assign n134 = ~x6 & x7 ;
  assign n135 = ( x1 & n133 ) | ( x1 & n134 ) | ( n133 & n134 ) ;
  assign n136 = ~x1 & n135 ;
  assign n152 = ( x0 & x2 ) | ( x0 & ~n136 ) | ( x2 & ~n136 ) ;
  assign n141 = x1 | x5 ;
  assign n139 = x4 | x6 ;
  assign n142 = ( x1 & ~x5 ) | ( x1 & n139 ) | ( ~x5 & n139 ) ;
  assign n137 = x4 | x5 ;
  assign n138 = ( ~x4 & n87 ) | ( ~x4 & n137 ) | ( n87 & n137 ) ;
  assign n140 = ( n80 & n87 ) | ( n80 & n138 ) | ( n87 & n138 ) ;
  assign n143 = x1 & n140 ;
  assign n144 = ( n141 & ~n142 ) | ( n141 & n143 ) | ( ~n142 & n143 ) ;
  assign n145 = x13 & ~n144 ;
  assign n146 = x3 & n138 ;
  assign n147 = x13 | n146 ;
  assign n148 = ~n145 & n147 ;
  assign n149 = ~x7 & x8 ;
  assign n150 = ( x12 & n148 ) | ( x12 & ~n149 ) | ( n148 & ~n149 ) ;
  assign n151 = n148 & ~n150 ;
  assign n153 = x2 & n151 ;
  assign n154 = ( n136 & n152 ) | ( n136 & n153 ) | ( n152 & n153 ) ;
  assign n156 = ~x2 & x5 ;
  assign n159 = ~x1 & x2 ;
  assign n160 = ( x4 & ~n156 ) | ( x4 & n159 ) | ( ~n156 & n159 ) ;
  assign n161 = x0 & ~n160 ;
  assign n158 = x1 & x4 ;
  assign n162 = x0 | n158 ;
  assign n163 = ( ~x0 & n161 ) | ( ~x0 & n162 ) | ( n161 & n162 ) ;
  assign n164 = ~x6 & x12 ;
  assign n165 = ( x7 & ~n163 ) | ( x7 & n164 ) | ( ~n163 & n164 ) ;
  assign n166 = n163 & n165 ;
  assign n155 = ~x12 & n149 ;
  assign n157 = n155 & n156 ;
  assign n167 = n157 & ~n166 ;
  assign n168 = x3 & ~x13 ;
  assign n169 = ( n166 & n167 ) | ( n166 & n168 ) | ( n167 & n168 ) ;
  assign n170 = ( ~x1 & x2 ) | ( ~x1 & x4 ) | ( x2 & x4 ) ;
  assign n171 = x4 & x5 ;
  assign n172 = ( x2 & x4 ) | ( x2 & n171 ) | ( x4 & n171 ) ;
  assign n173 = ( n158 & n170 ) | ( n158 & ~n172 ) | ( n170 & ~n172 ) ;
  assign n174 = n81 & n159 ;
  assign n175 = x3 | n174 ;
  assign n176 = ( ~n173 & n174 ) | ( ~n173 & n175 ) | ( n174 & n175 ) ;
  assign n177 = x0 & ~n176 ;
  assign n178 = x1 & n130 ;
  assign n179 = x0 | n178 ;
  assign n180 = ~n177 & n179 ;
  assign n191 = x6 & n95 ;
  assign n192 = x10 | n191 ;
  assign n193 = ( ~x11 & n191 ) | ( ~x11 & n192 ) | ( n191 & n192 ) ;
  assign n194 = n180 & n193 ;
  assign n195 = x12 & ~n194 ;
  assign n187 = ( x2 & x4 ) | ( x2 & ~n73 ) | ( x4 & ~n73 ) ;
  assign n188 = ~x5 & n187 ;
  assign n189 = ( ~x5 & n73 ) | ( ~x5 & n187 ) | ( n73 & n187 ) ;
  assign n190 = ( n73 & n188 ) | ( n73 & ~n189 ) | ( n188 & ~n189 ) ;
  assign n196 = x3 & n190 ;
  assign n197 = x12 | n196 ;
  assign n198 = ~n195 & n197 ;
  assign n199 = ~x13 & n198 ;
  assign n184 = x13 & n144 ;
  assign n185 = ( x12 & n73 ) | ( x12 & ~n184 ) | ( n73 & ~n184 ) ;
  assign n186 = n73 & ~n185 ;
  assign n200 = n186 | n199 ;
  assign n201 = ( x2 & n199 ) | ( x2 & n200 ) | ( n199 & n200 ) ;
  assign n202 = x7 & n201 ;
  assign n181 = x12 & n103 ;
  assign n182 = ( x13 & n180 ) | ( x13 & ~n181 ) | ( n180 & ~n181 ) ;
  assign n183 = n180 & ~n182 ;
  assign n203 = n183 | n202 ;
  assign n204 = ( x6 & n202 ) | ( x6 & n203 ) | ( n202 & n203 ) ;
  assign n205 = ( ~n154 & n169 ) | ( ~n154 & n204 ) | ( n169 & n204 ) ;
  assign n206 = n68 | n204 ;
  assign n207 = ( n154 & n205 ) | ( n154 & n206 ) | ( n205 & n206 ) ;
  assign n233 = x3 & ~n158 ;
  assign n234 = x0 & n233 ;
  assign n230 = x0 & ~x2 ;
  assign n231 = x1 & ~x3 ;
  assign n232 = ( ~x0 & n230 ) | ( ~x0 & n231 ) | ( n230 & n231 ) ;
  assign n235 = n193 & n232 ;
  assign n236 = ( n193 & n234 ) | ( n193 & n235 ) | ( n234 & n235 ) ;
  assign n213 = x2 | x3 ;
  assign n238 = x2 & ~x3 ;
  assign n241 = ( ~x2 & n213 ) | ( ~x2 & n238 ) | ( n213 & n238 ) ;
  assign n242 = n73 & n241 ;
  assign n243 = x12 | n242 ;
  assign n237 = x0 | x1 ;
  assign n239 = x0 & ~n238 ;
  assign n240 = n237 & ~n239 ;
  assign n244 = n193 & n240 ;
  assign n245 = x12 & ~n244 ;
  assign n246 = n243 & ~n245 ;
  assign n247 = x4 & n246 ;
  assign n248 = x12 | n247 ;
  assign n249 = ( n236 & n247 ) | ( n236 & n248 ) | ( n247 & n248 ) ;
  assign n250 = ~x13 & n249 ;
  assign n223 = x1 | x2 ;
  assign n224 = ~x2 & x3 ;
  assign n225 = x1 & n224 ;
  assign n226 = ( ~x1 & n223 ) | ( ~x1 & n225 ) | ( n223 & n225 ) ;
  assign n227 = x13 & n226 ;
  assign n228 = ( x12 & n73 ) | ( x12 & ~n227 ) | ( n73 & ~n227 ) ;
  assign n229 = n73 & ~n228 ;
  assign n251 = n229 | n250 ;
  assign n252 = ( x4 & n250 ) | ( x4 & n251 ) | ( n250 & n251 ) ;
  assign n253 = x7 & n252 ;
  assign n208 = ( x1 & ~x3 ) | ( x1 & x4 ) | ( ~x3 & x4 ) ;
  assign n209 = x3 & ~n208 ;
  assign n210 = ~x3 & x4 ;
  assign n211 = ( x2 & n209 ) | ( x2 & n210 ) | ( n209 & n210 ) ;
  assign n212 = n209 | n211 ;
  assign n214 = x0 & ~n213 ;
  assign n215 = ~x0 & n15 ;
  assign n216 = ( x0 & ~n214 ) | ( x0 & n215 ) | ( ~n214 & n215 ) ;
  assign n217 = x1 & ~n216 ;
  assign n218 = x0 | n217 ;
  assign n219 = ( n212 & n217 ) | ( n212 & n218 ) | ( n217 & n218 ) ;
  assign n220 = x12 & n219 ;
  assign n221 = ( x13 & n103 ) | ( x13 & ~n220 ) | ( n103 & ~n220 ) ;
  assign n222 = n103 & ~n221 ;
  assign n254 = n222 | n253 ;
  assign n255 = ( x6 & n253 ) | ( x6 & n254 ) | ( n253 & n254 ) ;
  assign n288 = ~x5 & n255 ;
  assign n262 = x4 & ~x13 ;
  assign n263 = ( x2 & x5 ) | ( x2 & n262 ) | ( x5 & n262 ) ;
  assign n264 = ~x5 & n263 ;
  assign n256 = ~x3 & x6 ;
  assign n257 = ( x5 & n224 ) | ( x5 & ~n256 ) | ( n224 & ~n256 ) ;
  assign n258 = ~x5 & x6 ;
  assign n259 = n224 & n258 ;
  assign n260 = x4 | n259 ;
  assign n261 = ( ~n257 & n259 ) | ( ~n257 & n260 ) | ( n259 & n260 ) ;
  assign n265 = ( x1 & n261 ) | ( x1 & n264 ) | ( n261 & n264 ) ;
  assign n266 = x13 & ~n265 ;
  assign n267 = ( x13 & n264 ) | ( x13 & ~n266 ) | ( n264 & ~n266 ) ;
  assign n268 = x7 & n73 ;
  assign n269 = ( x12 & n267 ) | ( x12 & ~n268 ) | ( n267 & ~n268 ) ;
  assign n270 = n267 & ~n269 ;
  assign n271 = ( x8 & n32 ) | ( x8 & ~n226 ) | ( n32 & ~n226 ) ;
  assign n272 = n226 & n271 ;
  assign n273 = ( x12 & ~n149 ) | ( x12 & n241 ) | ( ~n149 & n241 ) ;
  assign n274 = n241 & ~n273 ;
  assign n277 = ( ~x4 & x13 ) | ( ~x4 & n274 ) | ( x13 & n274 ) ;
  assign n275 = ( x7 & n164 ) | ( x7 & ~n219 ) | ( n164 & ~n219 ) ;
  assign n276 = n219 & n275 ;
  assign n278 = ~x13 & n276 ;
  assign n279 = ( n274 & ~n277 ) | ( n274 & n278 ) | ( ~n277 & n278 ) ;
  assign n280 = ( x4 & ~x7 ) | ( x4 & n279 ) | ( ~x7 & n279 ) ;
  assign n281 = n272 & ~n280 ;
  assign n282 = ( n272 & n279 ) | ( n272 & ~n281 ) | ( n279 & ~n281 ) ;
  assign n285 = ( x5 & n68 ) | ( x5 & ~n282 ) | ( n68 & ~n282 ) ;
  assign n283 = ( x12 & ~n149 ) | ( x12 & n267 ) | ( ~n149 & n267 ) ;
  assign n284 = n267 & ~n283 ;
  assign n286 = n68 & n284 ;
  assign n287 = ( n282 & n285 ) | ( n282 & n286 ) | ( n285 & n286 ) ;
  assign n289 = n270 | n287 ;
  assign n290 = ( n255 & ~n288 ) | ( n255 & n289 ) | ( ~n288 & n289 ) ;
  assign n291 = ( x4 & x5 ) | ( x4 & ~x13 ) | ( x5 & ~x13 ) ;
  assign n292 = ( x3 & x4 ) | ( x3 & x13 ) | ( x4 & x13 ) ;
  assign n293 = n291 & ~n292 ;
  assign n294 = ( ~x5 & n291 ) | ( ~x5 & n293 ) | ( n291 & n293 ) ;
  assign n295 = x2 & ~x4 ;
  assign n296 = ( x2 & x5 ) | ( x2 & n295 ) | ( x5 & n295 ) ;
  assign n297 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n298 = ( ~x3 & x4 ) | ( ~x3 & n295 ) | ( x4 & n295 ) ;
  assign n299 = n297 | n298 ;
  assign n300 = ( n295 & ~n296 ) | ( n295 & n299 ) | ( ~n296 & n299 ) ;
  assign n301 = x13 & n300 ;
  assign n302 = x1 & n301 ;
  assign n303 = x2 | n302 ;
  assign n304 = ( n294 & n302 ) | ( n294 & n303 ) | ( n302 & n303 ) ;
  assign n305 = ( x12 & ~n268 ) | ( x12 & n304 ) | ( ~n268 & n304 ) ;
  assign n306 = n304 & ~n305 ;
  assign n384 = ~x6 & n306 ;
  assign n307 = ( x1 & x2 ) | ( x1 & x5 ) | ( x2 & x5 ) ;
  assign n308 = x5 & n15 ;
  assign n309 = ( ~x1 & n307 ) | ( ~x1 & n308 ) | ( n307 & n308 ) ;
  assign n310 = ( ~x2 & x3 ) | ( ~x2 & x5 ) | ( x3 & x5 ) ;
  assign n311 = x4 & ~n310 ;
  assign n312 = ( ~x0 & x2 ) | ( ~x0 & x5 ) | ( x2 & x5 ) ;
  assign n313 = ( x0 & x3 ) | ( x0 & x5 ) | ( x3 & x5 ) ;
  assign n314 = ~n312 & n313 ;
  assign n315 = ( ~x0 & x3 ) | ( ~x0 & x5 ) | ( x3 & x5 ) ;
  assign n316 = ~x0 & x4 ;
  assign n317 = ( ~x3 & n315 ) | ( ~x3 & n316 ) | ( n315 & n316 ) ;
  assign n318 = ( x1 & n314 ) | ( x1 & n317 ) | ( n314 & n317 ) ;
  assign n319 = ~n87 & n318 ;
  assign n320 = ( x1 & n87 ) | ( x1 & n319 ) | ( n87 & n319 ) ;
  assign n321 = ( ~n309 & n311 ) | ( ~n309 & n320 ) | ( n311 & n320 ) ;
  assign n322 = x0 | n320 ;
  assign n323 = ( n309 & n321 ) | ( n309 & n322 ) | ( n321 & n322 ) ;
  assign n324 = ( ~x7 & x10 ) | ( ~x7 & x11 ) | ( x10 & x11 ) ;
  assign n325 = ( x7 & ~x9 ) | ( x7 & n324 ) | ( ~x9 & n324 ) ;
  assign n326 = ( x7 & x10 ) | ( x7 & ~n325 ) | ( x10 & ~n325 ) ;
  assign n327 = n324 | n326 ;
  assign n328 = ~x9 & n327 ;
  assign n329 = ( ~n325 & n327 ) | ( ~n325 & n328 ) | ( n327 & n328 ) ;
  assign n330 = x12 & n329 ;
  assign n331 = ( x13 & n323 ) | ( x13 & ~n330 ) | ( n323 & ~n330 ) ;
  assign n332 = n323 & ~n331 ;
  assign n350 = ( x6 & x8 ) | ( x6 & ~n332 ) | ( x8 & ~n332 ) ;
  assign n333 = x6 & ~x12 ;
  assign n334 = ( x7 & n301 ) | ( x7 & n333 ) | ( n301 & n333 ) ;
  assign n335 = ~x7 & n334 ;
  assign n347 = ( x1 & n68 ) | ( x1 & ~n335 ) | ( n68 & ~n335 ) ;
  assign n336 = ( x4 & x5 ) | ( x4 & ~x12 ) | ( x5 & ~x12 ) ;
  assign n337 = ( x3 & x4 ) | ( x3 & x12 ) | ( x4 & x12 ) ;
  assign n338 = n336 & ~n337 ;
  assign n339 = ( ~x5 & n336 ) | ( ~x5 & n338 ) | ( n336 & n338 ) ;
  assign n340 = ~x7 & n339 ;
  assign n341 = x6 & n340 ;
  assign n344 = ( ~x2 & x13 ) | ( ~x2 & n341 ) | ( x13 & n341 ) ;
  assign n342 = ( x7 & n164 ) | ( x7 & ~n323 ) | ( n164 & ~n323 ) ;
  assign n343 = n323 & n342 ;
  assign n345 = ~x13 & n343 ;
  assign n346 = ( n341 & ~n344 ) | ( n341 & n345 ) | ( ~n344 & n345 ) ;
  assign n348 = n68 & n346 ;
  assign n349 = ( n335 & n347 ) | ( n335 & n348 ) | ( n347 & n348 ) ;
  assign n351 = x8 & n349 ;
  assign n352 = ( n332 & n350 ) | ( n332 & n351 ) | ( n350 & n351 ) ;
  assign n353 = x2 & ~x13 ;
  assign n354 = x2 & ~n353 ;
  assign n355 = ~x1 & n354 ;
  assign n356 = ( x3 & ~n353 ) | ( x3 & n354 ) | ( ~n353 & n354 ) ;
  assign n357 = ( ~x13 & n355 ) | ( ~x13 & n356 ) | ( n355 & n356 ) ;
  assign n358 = x7 & n357 ;
  assign n359 = ( x12 & n73 ) | ( x12 & ~n358 ) | ( n73 & ~n358 ) ;
  assign n360 = n73 & ~n359 ;
  assign n381 = ( ~x6 & n87 ) | ( ~x6 & n360 ) | ( n87 & n360 ) ;
  assign n363 = x6 & ~x7 ;
  assign n364 = x7 & x12 ;
  assign n365 = x0 & ~x6 ;
  assign n366 = x12 & ~n365 ;
  assign n367 = ( n363 & n364 ) | ( n363 & ~n366 ) | ( n364 & ~n366 ) ;
  assign n368 = ( x13 & ~n224 ) | ( x13 & n367 ) | ( ~n224 & n367 ) ;
  assign n369 = n367 & ~n368 ;
  assign n361 = ~x1 & x6 ;
  assign n362 = x2 & n361 ;
  assign n370 = ( ~x7 & n362 ) | ( ~x7 & n369 ) | ( n362 & n369 ) ;
  assign n371 = n32 & ~n370 ;
  assign n372 = ( n32 & n369 ) | ( n32 & ~n371 ) | ( n369 & ~n371 ) ;
  assign n378 = ( x8 & n68 ) | ( x8 & ~n372 ) | ( n68 & ~n372 ) ;
  assign n373 = x6 & ~x13 ;
  assign n374 = ( x12 & ~n329 ) | ( x12 & n373 ) | ( ~n329 & n373 ) ;
  assign n375 = n329 & n374 ;
  assign n376 = ( x2 & n37 ) | ( x2 & n375 ) | ( n37 & n375 ) ;
  assign n377 = ~x2 & n376 ;
  assign n379 = x8 & n377 ;
  assign n380 = ( n372 & n378 ) | ( n372 & n379 ) | ( n378 & n379 ) ;
  assign n382 = ~n87 & n380 ;
  assign n383 = ( n360 & ~n381 ) | ( n360 & n382 ) | ( ~n381 & n382 ) ;
  assign n385 = n352 | n383 ;
  assign n386 = ( n306 & ~n384 ) | ( n306 & n385 ) | ( ~n384 & n385 ) ;
  assign n387 = x5 & x13 ;
  assign n388 = x5 & ~n387 ;
  assign n389 = x2 & n388 ;
  assign n390 = ( n158 & ~n387 ) | ( n158 & n388 ) | ( ~n387 & n388 ) ;
  assign n391 = ( x13 & n389 ) | ( x13 & n390 ) | ( n389 & n390 ) ;
  assign n392 = ~x13 & n224 ;
  assign n393 = ( x1 & ~n22 ) | ( x1 & n392 ) | ( ~n22 & n392 ) ;
  assign n394 = x13 & ~n393 ;
  assign n395 = ( x13 & n392 ) | ( x13 & ~n394 ) | ( n392 & ~n394 ) ;
  assign n396 = ( x1 & x6 ) | ( x1 & ~x13 ) | ( x6 & ~x13 ) ;
  assign n397 = ( x4 & x6 ) | ( x4 & x13 ) | ( x6 & x13 ) ;
  assign n398 = n396 & n397 ;
  assign n399 = x5 & ~x13 ;
  assign n400 = x1 & ~x6 ;
  assign n401 = x13 & ~n400 ;
  assign n402 = n399 | n401 ;
  assign n403 = x4 & ~n402 ;
  assign n404 = x5 | n403 ;
  assign n405 = ( ~n398 & n403 ) | ( ~n398 & n404 ) | ( n403 & n404 ) ;
  assign n406 = x2 & n405 ;
  assign n407 = x5 | n406 ;
  assign n408 = ( n395 & n406 ) | ( n395 & n407 ) | ( n406 & n407 ) ;
  assign n409 = x3 & ~n408 ;
  assign n410 = ( n391 & n408 ) | ( n391 & ~n409 ) | ( n408 & ~n409 ) ;
  assign n411 = x8 & ~x9 ;
  assign n412 = ( x8 & x10 ) | ( x8 & n411 ) | ( x10 & n411 ) ;
  assign n413 = ( ~x8 & x10 ) | ( ~x8 & n411 ) | ( x10 & n411 ) ;
  assign n414 = ( x8 & ~n412 ) | ( x8 & n413 ) | ( ~n412 & n413 ) ;
  assign n415 = n410 & n414 ;
  assign n416 = x4 | n224 ;
  assign n417 = ( ~n86 & n224 ) | ( ~n86 & n416 ) | ( n224 & n416 ) ;
  assign n418 = ( x1 & ~x2 ) | ( x1 & x3 ) | ( ~x2 & x3 ) ;
  assign n419 = ( x1 & x2 ) | ( x1 & ~x4 ) | ( x2 & ~x4 ) ;
  assign n420 = ~n418 & n419 ;
  assign n421 = x1 | n420 ;
  assign n422 = ( n417 & n420 ) | ( n417 & n421 ) | ( n420 & n421 ) ;
  assign n423 = x13 & n414 ;
  assign n424 = ( x12 & n422 ) | ( x12 & ~n423 ) | ( n422 & ~n423 ) ;
  assign n425 = n422 & ~n424 ;
  assign n478 = ( x6 & x7 ) | ( x6 & ~n425 ) | ( x7 & ~n425 ) ;
  assign n426 = x2 & x5 ;
  assign n427 = x1 & ~n311 ;
  assign n428 = ( n311 & n426 ) | ( n311 & ~n427 ) | ( n426 & ~n427 ) ;
  assign n433 = x9 & ~x11 ;
  assign n434 = ~x7 & x9 ;
  assign n435 = ( ~x8 & x9 ) | ( ~x8 & n434 ) | ( x9 & n434 ) ;
  assign n436 = ( n98 & n433 ) | ( n98 & ~n435 ) | ( n433 & ~n435 ) ;
  assign n437 = ( ~x0 & n428 ) | ( ~x0 & n436 ) | ( n428 & n436 ) ;
  assign n429 = x5 & ~n230 ;
  assign n430 = n137 & ~n429 ;
  assign n431 = x1 & n430 ;
  assign n432 = ( x1 & n317 ) | ( x1 & n431 ) | ( n317 & n431 ) ;
  assign n438 = n432 & ~n436 ;
  assign n439 = ( n428 & ~n437 ) | ( n428 & n438 ) | ( ~n437 & n438 ) ;
  assign n443 = x12 & ~n436 ;
  assign n444 = x5 & n443 ;
  assign n451 = ( ~x0 & x2 ) | ( ~x0 & n444 ) | ( x2 & n444 ) ;
  assign n448 = ( ~x0 & x4 ) | ( ~x0 & n443 ) | ( x4 & n443 ) ;
  assign n445 = x8 & x9 ;
  assign n446 = x7 & ~n445 ;
  assign n447 = ~x12 & n446 ;
  assign n449 = ~x4 & n447 ;
  assign n450 = ( n443 & ~n448 ) | ( n443 & n449 ) | ( ~n448 & n449 ) ;
  assign n452 = ~x2 & n450 ;
  assign n453 = ( n444 & ~n451 ) | ( n444 & n452 ) | ( ~n451 & n452 ) ;
  assign n440 = ( x1 & x5 ) | ( x1 & ~n436 ) | ( x5 & ~n436 ) ;
  assign n441 = ( x4 & x5 ) | ( x4 & n436 ) | ( x5 & n436 ) ;
  assign n442 = n440 & ~n441 ;
  assign n454 = ( x0 & n442 ) | ( x0 & n453 ) | ( n442 & n453 ) ;
  assign n455 = x12 & ~n454 ;
  assign n456 = ( x12 & n453 ) | ( x12 & ~n455 ) | ( n453 & ~n455 ) ;
  assign n457 = x3 & n456 ;
  assign n458 = x12 | n457 ;
  assign n459 = ( n439 & n457 ) | ( n439 & n458 ) | ( n457 & n458 ) ;
  assign n475 = ( ~x10 & x13 ) | ( ~x10 & n459 ) | ( x13 & n459 ) ;
  assign n461 = ( x2 & x4 ) | ( x2 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n462 = x3 & ~n461 ;
  assign n463 = ( n320 & n428 ) | ( n320 & ~n462 ) | ( n428 & ~n462 ) ;
  assign n464 = ( n322 & n462 ) | ( n322 & n463 ) | ( n462 & n463 ) ;
  assign n465 = ( x8 & n67 ) | ( x8 & n464 ) | ( n67 & n464 ) ;
  assign n460 = x9 & ~x10 ;
  assign n466 = n460 & n464 ;
  assign n467 = ( ~x8 & n465 ) | ( ~x8 & n466 ) | ( n465 & n466 ) ;
  assign n472 = ( x7 & x12 ) | ( x7 & ~n467 ) | ( x12 & ~n467 ) ;
  assign n468 = ~x2 & n15 ;
  assign n469 = ~x12 & n445 ;
  assign n470 = ( x10 & n468 ) | ( x10 & n469 ) | ( n468 & n469 ) ;
  assign n471 = ~x10 & n470 ;
  assign n473 = x7 & n471 ;
  assign n474 = ( n467 & n472 ) | ( n467 & n473 ) | ( n472 & n473 ) ;
  assign n476 = ~x13 & n474 ;
  assign n477 = ( n459 & ~n475 ) | ( n459 & n476 ) | ( ~n475 & n476 ) ;
  assign n479 = x6 & n477 ;
  assign n480 = ( n425 & n478 ) | ( n425 & n479 ) | ( n478 & n479 ) ;
  assign n481 = ( x7 & ~x12 ) | ( x7 & n480 ) | ( ~x12 & n480 ) ;
  assign n482 = n415 & ~n481 ;
  assign n483 = ( n415 & n480 ) | ( n415 & ~n482 ) | ( n480 & ~n482 ) ;
  assign n495 = ~x4 & x6 ;
  assign n496 = x5 | n495 ;
  assign n525 = ( x12 & ~n357 ) | ( x12 & n496 ) | ( ~n357 & n496 ) ;
  assign n501 = ( ~x2 & x3 ) | ( ~x2 & x6 ) | ( x3 & x6 ) ;
  assign n502 = ( x2 & x4 ) | ( x2 & x6 ) | ( x4 & x6 ) ;
  assign n503 = ~n501 & n502 ;
  assign n497 = ( x3 & x5 ) | ( x3 & ~x6 ) | ( x5 & ~x6 ) ;
  assign n498 = x4 & ~n497 ;
  assign n499 = ~x2 & x6 ;
  assign n500 = x3 & n499 ;
  assign n504 = ( x13 & n498 ) | ( x13 & n500 ) | ( n498 & n500 ) ;
  assign n505 = ~n503 & n504 ;
  assign n506 = ( x13 & n503 ) | ( x13 & n505 ) | ( n503 & n505 ) ;
  assign n522 = ~x1 & n506 ;
  assign n513 = x2 | x13 ;
  assign n514 = x1 & x3 ;
  assign n515 = x13 & ~n514 ;
  assign n516 = n513 & ~n515 ;
  assign n517 = ~x6 & n516 ;
  assign n518 = ( ~x4 & n516 ) | ( ~x4 & n517 ) | ( n516 & n517 ) ;
  assign n507 = ( ~x2 & x6 ) | ( ~x2 & x13 ) | ( x6 & x13 ) ;
  assign n508 = ( x2 & ~x3 ) | ( x2 & x13 ) | ( ~x3 & x13 ) ;
  assign n509 = ~n507 & n508 ;
  assign n510 = ~x6 & x13 ;
  assign n511 = ( x1 & x4 ) | ( x1 & n510 ) | ( x4 & n510 ) ;
  assign n512 = ~x4 & n511 ;
  assign n519 = ( x5 & n509 ) | ( x5 & n512 ) | ( n509 & n512 ) ;
  assign n520 = ~n518 & n519 ;
  assign n521 = ( x5 & n518 ) | ( x5 & n520 ) | ( n518 & n520 ) ;
  assign n523 = n264 | n521 ;
  assign n524 = ( n506 & ~n522 ) | ( n506 & n523 ) | ( ~n522 & n523 ) ;
  assign n526 = ~x12 & n524 ;
  assign n527 = ( n496 & ~n525 ) | ( n496 & n526 ) | ( ~n525 & n526 ) ;
  assign n539 = x9 & x10 ;
  assign n540 = x9 & ~n539 ;
  assign n541 = n527 & n540 ;
  assign n528 = ~x4 & n224 ;
  assign n529 = ~x12 & n528 ;
  assign n530 = x12 & n464 ;
  assign n531 = x13 & n422 ;
  assign n532 = ~x12 & n531 ;
  assign n533 = ( ~n529 & n530 ) | ( ~n529 & n532 ) | ( n530 & n532 ) ;
  assign n534 = x13 & ~n532 ;
  assign n535 = ( n529 & n533 ) | ( n529 & ~n534 ) | ( n533 & ~n534 ) ;
  assign n536 = ~x12 & n410 ;
  assign n537 = x6 | n536 ;
  assign n538 = ( n535 & n536 ) | ( n535 & n537 ) | ( n536 & n537 ) ;
  assign n542 = ( n538 & ~n539 ) | ( n538 & n540 ) | ( ~n539 & n540 ) ;
  assign n543 = ( x10 & n541 ) | ( x10 & n542 ) | ( n541 & n542 ) ;
  assign n544 = x7 & ~n543 ;
  assign n545 = x10 & n527 ;
  assign n546 = x7 | n545 ;
  assign n547 = ~n544 & n546 ;
  assign n548 = x8 & n547 ;
  assign n488 = x6 | x10 ;
  assign n489 = ( x6 & ~x10 ) | ( x6 & n94 ) | ( ~x10 & n94 ) ;
  assign n484 = x8 | x11 ;
  assign n485 = ( x8 & x10 ) | ( x8 & ~n484 ) | ( x10 & ~n484 ) ;
  assign n486 = ( ~x9 & x10 ) | ( ~x9 & n485 ) | ( x10 & n485 ) ;
  assign n487 = ( n460 & ~n485 ) | ( n460 & n486 ) | ( ~n485 & n486 ) ;
  assign n490 = x6 & n487 ;
  assign n491 = ( n488 & ~n489 ) | ( n488 & n490 ) | ( ~n489 & n490 ) ;
  assign n492 = x12 & n491 ;
  assign n493 = ( x13 & n464 ) | ( x13 & ~n492 ) | ( n464 & ~n492 ) ;
  assign n494 = n464 & ~n493 ;
  assign n549 = n494 | n548 ;
  assign n550 = ( x7 & n548 ) | ( x7 & n549 ) | ( n548 & n549 ) ;
  assign n551 = ~x13 & n530 ;
  assign n552 = ( x10 & n69 ) | ( x10 & n551 ) | ( n69 & n551 ) ;
  assign n553 = ~x10 & n552 ;
  assign n572 = ( x7 & x10 ) | ( x7 & n538 ) | ( x10 & n538 ) ;
  assign n573 = ~x10 & n572 ;
  assign n574 = ( ~x7 & x8 ) | ( ~x7 & n573 ) | ( x8 & n573 ) ;
  assign n575 = ( n572 & n573 ) | ( n572 & n574 ) | ( n573 & n574 ) ;
  assign n554 = x10 & x11 ;
  assign n555 = ( ~x10 & n530 ) | ( ~x10 & n554 ) | ( n530 & n554 ) ;
  assign n556 = x7 & n468 ;
  assign n557 = ( x10 & x12 ) | ( x10 & n556 ) | ( x12 & n556 ) ;
  assign n558 = ~x12 & n557 ;
  assign n559 = x10 & n532 ;
  assign n560 = x7 & n559 ;
  assign n561 = ( ~n555 & n558 ) | ( ~n555 & n560 ) | ( n558 & n560 ) ;
  assign n562 = x13 & ~n560 ;
  assign n563 = ( n555 & n561 ) | ( n555 & ~n562 ) | ( n561 & ~n562 ) ;
  assign n566 = ( ~x6 & x8 ) | ( ~x6 & n563 ) | ( x8 & n563 ) ;
  assign n564 = x10 & n536 ;
  assign n565 = x7 & n564 ;
  assign n567 = ~x8 & n565 ;
  assign n568 = ( n563 & ~n566 ) | ( n563 & n567 ) | ( ~n566 & n567 ) ;
  assign n569 = x10 & n551 ;
  assign n570 = ( x6 & x7 ) | ( x6 & n569 ) | ( x7 & n569 ) ;
  assign n571 = ~x6 & n570 ;
  assign n576 = ( x9 & n568 ) | ( x9 & n571 ) | ( n568 & n571 ) ;
  assign n577 = ~n575 & n576 ;
  assign n578 = ( x9 & n575 ) | ( x9 & n577 ) | ( n575 & n577 ) ;
  assign n579 = ( x6 & ~x7 ) | ( x6 & n578 ) | ( ~x7 & n578 ) ;
  assign n580 = n553 & ~n579 ;
  assign n581 = ( n553 & n578 ) | ( n553 & ~n580 ) | ( n578 & ~n580 ) ;
  assign n599 = ( x6 & x9 ) | ( x6 & n530 ) | ( x9 & n530 ) ;
  assign n596 = x9 & n468 ;
  assign n597 = ( x10 & x12 ) | ( x10 & n596 ) | ( x12 & n596 ) ;
  assign n598 = ~x12 & n597 ;
  assign n600 = x6 & n598 ;
  assign n601 = ( ~x9 & n599 ) | ( ~x9 & n600 ) | ( n599 & n600 ) ;
  assign n593 = ( x2 & ~x12 ) | ( x2 & n86 ) | ( ~x12 & n86 ) ;
  assign n582 = x3 & x6 ;
  assign n583 = x4 & n582 ;
  assign n584 = x5 & ~n583 ;
  assign n585 = ( ~x5 & n137 ) | ( ~x5 & n584 ) | ( n137 & n584 ) ;
  assign n594 = ( x2 & x12 ) | ( x2 & ~n585 ) | ( x12 & ~n585 ) ;
  assign n595 = n593 & ~n594 ;
  assign n602 = ( x9 & n595 ) | ( x9 & n601 ) | ( n595 & n601 ) ;
  assign n603 = x10 & ~n602 ;
  assign n604 = ( x10 & n601 ) | ( x10 & ~n603 ) | ( n601 & ~n603 ) ;
  assign n605 = ~x8 & n604 ;
  assign n587 = x2 & ~n585 ;
  assign n586 = x3 & n496 ;
  assign n588 = ~x2 & n586 ;
  assign n589 = ( x2 & ~n587 ) | ( x2 & n588 ) | ( ~n587 & n588 ) ;
  assign n590 = ( x9 & x10 ) | ( x9 & ~n589 ) | ( x10 & ~n589 ) ;
  assign n591 = x9 & ~n590 ;
  assign n592 = ( x10 & ~n590 ) | ( x10 & n591 ) | ( ~n590 & n591 ) ;
  assign n606 = n592 | n605 ;
  assign n607 = ( ~x12 & n605 ) | ( ~x12 & n606 ) | ( n605 & n606 ) ;
  assign n628 = ~x7 & n607 ;
  assign n608 = ( x7 & ~x9 ) | ( x7 & x10 ) | ( ~x9 & x10 ) ;
  assign n609 = x9 & ~n608 ;
  assign n610 = ~x9 & x10 ;
  assign n611 = ( x8 & n609 ) | ( x8 & n610 ) | ( n609 & n610 ) ;
  assign n612 = n609 | n611 ;
  assign n613 = x12 & n612 ;
  assign n614 = ( x6 & ~n464 ) | ( x6 & n613 ) | ( ~n464 & n613 ) ;
  assign n615 = n464 & n614 ;
  assign n616 = ( ~x2 & x3 ) | ( ~x2 & x4 ) | ( x3 & x4 ) ;
  assign n617 = n78 & ~n616 ;
  assign n618 = ( ~x5 & n78 ) | ( ~x5 & n617 ) | ( n78 & n617 ) ;
  assign n619 = ~n588 & n618 ;
  assign n620 = ( n19 & n588 ) | ( n19 & n619 ) | ( n588 & n619 ) ;
  assign n625 = ( x7 & ~n460 ) | ( x7 & n620 ) | ( ~n460 & n620 ) ;
  assign n622 = ( x6 & ~x7 ) | ( x6 & n530 ) | ( ~x7 & n530 ) ;
  assign n621 = n155 & n426 ;
  assign n623 = ~x6 & n621 ;
  assign n624 = ( n530 & ~n622 ) | ( n530 & n623 ) | ( ~n622 & n623 ) ;
  assign n626 = ~n460 & n624 ;
  assign n627 = ( ~x7 & n625 ) | ( ~x7 & n626 ) | ( n625 & n626 ) ;
  assign n629 = n615 | n627 ;
  assign n630 = ( n607 & ~n628 ) | ( n607 & n629 ) | ( ~n628 & n629 ) ;
  assign n652 = ( ~x11 & x13 ) | ( ~x11 & n630 ) | ( x13 & n630 ) ;
  assign n631 = ( ~x1 & x3 ) | ( ~x1 & x6 ) | ( x3 & x6 ) ;
  assign n632 = ( x1 & x4 ) | ( x1 & x6 ) | ( x4 & x6 ) ;
  assign n633 = ~n631 & n632 ;
  assign n634 = x5 & ~x6 ;
  assign n635 = ( ~x4 & x5 ) | ( ~x4 & x6 ) | ( x5 & x6 ) ;
  assign n636 = x1 & x6 ;
  assign n637 = ( n634 & n635 ) | ( n634 & ~n636 ) | ( n635 & ~n636 ) ;
  assign n638 = x5 & ~n22 ;
  assign n639 = ( x1 & n498 ) | ( x1 & n500 ) | ( n498 & n500 ) ;
  assign n640 = ~n638 & n639 ;
  assign n641 = ( x1 & n638 ) | ( x1 & n640 ) | ( n638 & n640 ) ;
  assign n642 = ( ~n633 & n637 ) | ( ~n633 & n641 ) | ( n637 & n641 ) ;
  assign n643 = x2 | n641 ;
  assign n644 = ( n633 & n642 ) | ( n633 & n643 ) | ( n642 & n643 ) ;
  assign n645 = ( x7 & x9 ) | ( x7 & x10 ) | ( x9 & x10 ) ;
  assign n646 = ( ~x7 & x8 ) | ( ~x7 & x10 ) | ( x8 & x10 ) ;
  assign n647 = x9 & n646 ;
  assign n648 = ( n149 & n645 ) | ( n149 & ~n647 ) | ( n645 & ~n647 ) ;
  assign n649 = x13 & n648 ;
  assign n650 = ( x12 & n644 ) | ( x12 & ~n649 ) | ( n644 & ~n649 ) ;
  assign n651 = n644 & ~n650 ;
  assign n653 = x11 & n651 ;
  assign n654 = ( n630 & ~n652 ) | ( n630 & n653 ) | ( ~n652 & n653 ) ;
  assign n688 = ( x7 & x8 ) | ( x7 & x10 ) | ( x8 & x10 ) ;
  assign n689 = ( ~x9 & x10 ) | ( ~x9 & n688 ) | ( x10 & n688 ) ;
  assign n690 = x10 & ~n689 ;
  assign n691 = n689 | n690 ;
  assign n692 = ( ~x10 & n690 ) | ( ~x10 & n691 ) | ( n690 & n691 ) ;
  assign n693 = ( x12 & ~n156 ) | ( x12 & n692 ) | ( ~n156 & n692 ) ;
  assign n694 = n692 & ~n693 ;
  assign n681 = ( x7 & ~x8 ) | ( x7 & x9 ) | ( ~x8 & x9 ) ;
  assign n682 = ( x8 & x10 ) | ( x8 & ~n681 ) | ( x10 & ~n681 ) ;
  assign n683 = n681 & ~n682 ;
  assign n684 = n149 | n683 ;
  assign n695 = x0 & x12 ;
  assign n696 = ( x2 & ~n684 ) | ( x2 & n695 ) | ( ~n684 & n695 ) ;
  assign n697 = n684 & n696 ;
  assign n698 = ( x0 & x1 ) | ( x0 & n684 ) | ( x1 & n684 ) ;
  assign n699 = ( x0 & x5 ) | ( x0 & ~n684 ) | ( x5 & ~n684 ) ;
  assign n700 = n698 & ~n699 ;
  assign n701 = x12 & n700 ;
  assign n702 = x2 & n701 ;
  assign n703 = ( ~n694 & n697 ) | ( ~n694 & n702 ) | ( n697 & n702 ) ;
  assign n704 = x3 & ~n702 ;
  assign n705 = ( n694 & n703 ) | ( n694 & ~n704 ) | ( n703 & ~n704 ) ;
  assign n706 = x4 & n705 ;
  assign n678 = x1 | n15 ;
  assign n679 = x0 & x5 ;
  assign n680 = ( n15 & ~n678 ) | ( n15 & n679 ) | ( ~n678 & n679 ) ;
  assign n674 = ( x0 & ~x1 ) | ( x0 & x5 ) | ( ~x1 & x5 ) ;
  assign n675 = ( x3 & x5 ) | ( x3 & ~n674 ) | ( x5 & ~n674 ) ;
  assign n676 = ( ~x0 & x3 ) | ( ~x0 & n674 ) | ( x3 & n674 ) ;
  assign n677 = n675 & ~n676 ;
  assign n685 = n677 & ~n680 ;
  assign n686 = x12 & n684 ;
  assign n687 = ( n680 & n685 ) | ( n680 & n686 ) | ( n685 & n686 ) ;
  assign n707 = n687 | n706 ;
  assign n708 = ( x2 & n706 ) | ( x2 & n707 ) | ( n706 & n707 ) ;
  assign n709 = x11 & n708 ;
  assign n656 = ( x7 & x9 ) | ( x7 & x11 ) | ( x9 & x11 ) ;
  assign n655 = x8 | x10 ;
  assign n657 = x9 & ~n655 ;
  assign n658 = ( ~x11 & n656 ) | ( ~x11 & n657 ) | ( n656 & n657 ) ;
  assign n671 = n99 & ~n658 ;
  assign n659 = x4 & ~n86 ;
  assign n660 = ~x1 & x5 ;
  assign n661 = ( ~x4 & n86 ) | ( ~x4 & n660 ) | ( n86 & n660 ) ;
  assign n662 = n659 | n661 ;
  assign n663 = ( x0 & ~x3 ) | ( x0 & x5 ) | ( ~x3 & x5 ) ;
  assign n664 = x0 & n663 ;
  assign n665 = ( x0 & x4 ) | ( x0 & ~n663 ) | ( x4 & ~n663 ) ;
  assign n666 = n663 | n665 ;
  assign n667 = ~n664 & n666 ;
  assign n668 = x1 & n667 ;
  assign n669 = x0 | n668 ;
  assign n670 = ( n662 & n668 ) | ( n662 & n669 ) | ( n668 & n669 ) ;
  assign n672 = x12 & n670 ;
  assign n673 = ( n658 & n671 ) | ( n658 & n672 ) | ( n671 & n672 ) ;
  assign n710 = n673 | n709 ;
  assign n711 = ( x2 & n709 ) | ( x2 & n710 ) | ( n709 & n710 ) ;
  assign n733 = ( ~x6 & x13 ) | ( ~x6 & n711 ) | ( x13 & n711 ) ;
  assign n715 = n36 | n213 ;
  assign n716 = x11 | n655 ;
  assign n717 = x12 | n716 ;
  assign n727 = ( x6 & ~n715 ) | ( x6 & n717 ) | ( ~n715 & n717 ) ;
  assign n723 = ( x2 & ~n68 ) | ( x2 & n672 ) | ( ~n68 & n672 ) ;
  assign n724 = n68 & n723 ;
  assign n718 = ~x5 & x8 ;
  assign n719 = ~n213 & n718 ;
  assign n720 = n539 & n719 ;
  assign n721 = ( x11 & x12 ) | ( x11 & n720 ) | ( x12 & n720 ) ;
  assign n722 = ~x12 & n721 ;
  assign n725 = x7 & n722 ;
  assign n726 = ( x7 & n724 ) | ( x7 & n725 ) | ( n724 & n725 ) ;
  assign n728 = ~x6 & n726 ;
  assign n729 = ( n715 & n727 ) | ( n715 & ~n728 ) | ( n727 & ~n728 ) ;
  assign n712 = ~x11 & x12 ;
  assign n713 = ( x10 & ~n670 ) | ( x10 & n712 ) | ( ~n670 & n712 ) ;
  assign n714 = n670 & n713 ;
  assign n730 = ( x2 & n714 ) | ( x2 & ~n729 ) | ( n714 & ~n729 ) ;
  assign n731 = x7 & ~n730 ;
  assign n732 = ( ~x7 & n729 ) | ( ~x7 & n731 ) | ( n729 & n731 ) ;
  assign n734 = x13 | n732 ;
  assign n735 = ( ~n711 & n733 ) | ( ~n711 & n734 ) | ( n733 & n734 ) ;
  assign n736 = x4 & x7 ;
  assign n737 = ( x5 & n213 ) | ( x5 & n736 ) | ( n213 & n736 ) ;
  assign n738 = ~n213 & n737 ;
  assign n739 = ~x10 & x11 ;
  assign n740 = ~x12 & n739 ;
  assign n741 = ~x9 & n740 ;
  assign n742 = x8 & n741 ;
  assign n752 = ( x13 & n738 ) | ( x13 & ~n742 ) | ( n738 & ~n742 ) ;
  assign n743 = ( x3 & n156 ) | ( x3 & ~n159 ) | ( n156 & ~n159 ) ;
  assign n744 = ~x3 & x5 ;
  assign n745 = ( x1 & x2 ) | ( x1 & n744 ) | ( x2 & n744 ) ;
  assign n746 = ~x2 & n745 ;
  assign n747 = x4 | n746 ;
  assign n748 = ( ~n743 & n746 ) | ( ~n743 & n747 ) | ( n746 & n747 ) ;
  assign n749 = x12 & n748 ;
  assign n750 = ( x0 & ~n105 ) | ( x0 & n749 ) | ( ~n105 & n749 ) ;
  assign n751 = n105 & n750 ;
  assign n753 = ~x13 & n751 ;
  assign n754 = ( n738 & ~n752 ) | ( n738 & n753 ) | ( ~n752 & n753 ) ;
  assign n755 = x1 | x4 ;
  assign n756 = x4 & ~n156 ;
  assign n757 = n755 & ~n756 ;
  assign n758 = x12 & n757 ;
  assign n759 = ( x13 & n105 ) | ( x13 & ~n758 ) | ( n105 & ~n758 ) ;
  assign n760 = n105 & ~n759 ;
  assign n798 = ( x0 & x3 ) | ( x0 & ~n760 ) | ( x3 & ~n760 ) ;
  assign n763 = x7 & ~n73 ;
  assign n764 = x8 & n68 ;
  assign n765 = x7 | n764 ;
  assign n766 = ~n763 & n765 ;
  assign n767 = x4 | n766 ;
  assign n761 = ~x8 & x9 ;
  assign n762 = n554 & n761 ;
  assign n768 = ~n36 & n762 ;
  assign n769 = x4 & ~n768 ;
  assign n770 = n767 & ~n769 ;
  assign n773 = x10 | x11 ;
  assign n774 = ~x4 & x11 ;
  assign n775 = ( x5 & n692 ) | ( x5 & ~n774 ) | ( n692 & ~n774 ) ;
  assign n776 = n692 & ~n775 ;
  assign n771 = x4 & ~x7 ;
  assign n772 = x5 & n771 ;
  assign n777 = ( n761 & n772 ) | ( n761 & n776 ) | ( n772 & n776 ) ;
  assign n778 = n773 | n777 ;
  assign n779 = ( ~n773 & n776 ) | ( ~n773 & n778 ) | ( n776 & n778 ) ;
  assign n780 = x1 & x13 ;
  assign n781 = ( x13 & n779 ) | ( x13 & ~n780 ) | ( n779 & ~n780 ) ;
  assign n782 = ( x13 & n770 ) | ( x13 & ~n780 ) | ( n770 & ~n780 ) ;
  assign n783 = ( n770 & n781 ) | ( n770 & ~n782 ) | ( n781 & ~n782 ) ;
  assign n795 = ( ~x2 & x12 ) | ( ~x2 & n783 ) | ( x12 & n783 ) ;
  assign n784 = x10 & n761 ;
  assign n785 = ( x11 & x13 ) | ( x11 & n784 ) | ( x13 & n784 ) ;
  assign n786 = ~x13 & n785 ;
  assign n789 = x2 | n87 ;
  assign n790 = x13 & n766 ;
  assign n791 = ( n87 & ~n789 ) | ( n87 & n790 ) | ( ~n789 & n790 ) ;
  assign n792 = x1 & n791 ;
  assign n787 = ~x2 & x4 ;
  assign n788 = ~n36 & n787 ;
  assign n793 = n788 | n792 ;
  assign n794 = ( n786 & n792 ) | ( n786 & n793 ) | ( n792 & n793 ) ;
  assign n796 = ~x12 & n794 ;
  assign n797 = ( n783 & ~n795 ) | ( n783 & n796 ) | ( ~n795 & n796 ) ;
  assign n799 = x3 & n797 ;
  assign n800 = ( n760 & n798 ) | ( n760 & n799 ) | ( n798 & n799 ) ;
  assign n806 = ( x0 & ~n68 ) | ( x0 & n749 ) | ( ~n68 & n749 ) ;
  assign n807 = n68 & n806 ;
  assign n803 = x10 & n445 ;
  assign n804 = ( x11 & x12 ) | ( x11 & n803 ) | ( x12 & n803 ) ;
  assign n805 = ~x12 & n804 ;
  assign n808 = ( ~n213 & n805 ) | ( ~n213 & n807 ) | ( n805 & n807 ) ;
  assign n809 = n137 | n808 ;
  assign n810 = ( ~n137 & n807 ) | ( ~n137 & n809 ) | ( n807 & n809 ) ;
  assign n817 = ( x6 & ~x7 ) | ( x6 & n810 ) | ( ~x7 & n810 ) ;
  assign n811 = x7 | x8 ;
  assign n812 = x11 | n811 ;
  assign n813 = ( ~x10 & x12 ) | ( ~x10 & n812 ) | ( x12 & n812 ) ;
  assign n814 = x10 | n813 ;
  assign n815 = n137 | n814 ;
  assign n816 = n213 | n815 ;
  assign n818 = x6 | n816 ;
  assign n819 = ( ~n810 & n817 ) | ( ~n810 & n818 ) | ( n817 & n818 ) ;
  assign n801 = ( x10 & n712 ) | ( x10 & ~n748 ) | ( n712 & ~n748 ) ;
  assign n802 = n748 & n801 ;
  assign n820 = ( x0 & n802 ) | ( x0 & ~n819 ) | ( n802 & ~n819 ) ;
  assign n821 = x7 & ~n820 ;
  assign n822 = ( ~x7 & n819 ) | ( ~x7 & n821 ) | ( n819 & n821 ) ;
  assign n839 = x0 & ~x13 ;
  assign n840 = ( x12 & ~n757 ) | ( x12 & n839 ) | ( ~n757 & n839 ) ;
  assign n841 = n757 & n840 ;
  assign n824 = x4 & ~x6 ;
  assign n825 = x1 & ~n824 ;
  assign n826 = n141 & ~n825 ;
  assign n827 = x2 & n826 ;
  assign n823 = ( ~x4 & x5 ) | ( ~x4 & n634 ) | ( x5 & n634 ) ;
  assign n828 = n823 | n827 ;
  assign n829 = ( x1 & n827 ) | ( x1 & n828 ) | ( n827 & n828 ) ;
  assign n830 = x13 & n829 ;
  assign n831 = ~x12 & n830 ;
  assign n842 = x13 & ~n445 ;
  assign n843 = ( x12 & n829 ) | ( x12 & ~n842 ) | ( n829 & ~n842 ) ;
  assign n844 = n829 & ~n843 ;
  assign n845 = ( n831 & ~n841 ) | ( n831 & n844 ) | ( ~n841 & n844 ) ;
  assign n846 = x11 & ~n844 ;
  assign n847 = ( n841 & n845 ) | ( n841 & ~n846 ) | ( n845 & ~n846 ) ;
  assign n848 = x10 & ~n847 ;
  assign n849 = x9 & n831 ;
  assign n850 = x10 | n849 ;
  assign n851 = ~n848 & n850 ;
  assign n852 = x7 & n851 ;
  assign n832 = ( x12 & n38 ) | ( x12 & ~n757 ) | ( n38 & ~n757 ) ;
  assign n833 = n757 & n832 ;
  assign n834 = ~x6 & n833 ;
  assign n835 = x0 & n834 ;
  assign n836 = ( ~x7 & n831 ) | ( ~x7 & n835 ) | ( n831 & n835 ) ;
  assign n837 = x8 & ~n836 ;
  assign n838 = ( x8 & n835 ) | ( x8 & ~n837 ) | ( n835 & ~n837 ) ;
  assign n853 = n838 | n852 ;
  assign n854 = ( n68 & n852 ) | ( n68 & n853 ) | ( n852 & n853 ) ;
  assign n855 = x3 & n854 ;
  assign n856 = x13 & ~n855 ;
  assign n857 = ( n822 & ~n855 ) | ( n822 & n856 ) | ( ~n855 & n856 ) ;
  assign n858 = ( n754 & ~n800 ) | ( n754 & n857 ) | ( ~n800 & n857 ) ;
  assign n859 = ~x6 & n857 ;
  assign n860 = ( ~n754 & n858 ) | ( ~n754 & n859 ) | ( n858 & n859 ) ;
  assign n861 = x11 | x13 ;
  assign n862 = x12 | n861 ;
  assign n863 = x8 | n72 ;
  assign n864 = n862 | n863 ;
  assign n900 = ~x9 & n32 ;
  assign n901 = n258 & n900 ;
  assign n897 = ( x6 & x9 ) | ( x6 & ~x12 ) | ( x9 & ~x12 ) ;
  assign n898 = ( x6 & x9 ) | ( x6 & ~x13 ) | ( x9 & ~x13 ) ;
  assign n899 = ~n897 & n898 ;
  assign n902 = ( ~x0 & n899 ) | ( ~x0 & n901 ) | ( n899 & n901 ) ;
  assign n903 = x5 & ~n902 ;
  assign n904 = ( x5 & n901 ) | ( x5 & ~n903 ) | ( n901 & ~n903 ) ;
  assign n905 = x7 & ~x10 ;
  assign n906 = ( x8 & ~n904 ) | ( x8 & n905 ) | ( ~n904 & n905 ) ;
  assign n907 = n904 & n906 ;
  assign n896 = n258 & ~n811 ;
  assign n908 = ( n32 & n896 ) | ( n32 & n907 ) | ( n896 & n907 ) ;
  assign n909 = n539 & ~n908 ;
  assign n910 = ( n539 & n907 ) | ( n539 & ~n909 ) | ( n907 & ~n909 ) ;
  assign n911 = x1 & n910 ;
  assign n894 = ( x13 & ~n333 ) | ( x13 & n692 ) | ( ~n333 & n692 ) ;
  assign n895 = n692 & ~n894 ;
  assign n912 = n895 | n911 ;
  assign n913 = ( ~x5 & n911 ) | ( ~x5 & n912 ) | ( n911 & n912 ) ;
  assign n914 = x4 | n913 ;
  assign n879 = x7 & ~x9 ;
  assign n880 = x7 | x9 ;
  assign n881 = ( ~x7 & n879 ) | ( ~x7 & n880 ) | ( n879 & n880 ) ;
  assign n888 = ~x10 & x13 ;
  assign n889 = ( x12 & n881 ) | ( x12 & ~n888 ) | ( n881 & ~n888 ) ;
  assign n890 = n881 & ~n889 ;
  assign n891 = x8 & n890 ;
  assign n892 = ( x5 & x6 ) | ( x5 & n891 ) | ( x6 & n891 ) ;
  assign n893 = ~x5 & n892 ;
  assign n915 = ~x1 & n893 ;
  assign n916 = x4 & ~n915 ;
  assign n917 = n914 & ~n916 ;
  assign n918 = x2 & ~n917 ;
  assign n882 = x10 | x13 ;
  assign n883 = ( x12 & n881 ) | ( x12 & n882 ) | ( n881 & n882 ) ;
  assign n884 = n881 & ~n883 ;
  assign n885 = x8 & n884 ;
  assign n886 = ( x5 & x6 ) | ( x5 & n885 ) | ( x6 & n885 ) ;
  assign n887 = ~x5 & n886 ;
  assign n919 = x4 & n887 ;
  assign n920 = x2 | n919 ;
  assign n921 = ~n918 & n920 ;
  assign n922 = x3 & ~n921 ;
  assign n868 = x7 & x8 ;
  assign n869 = ~x6 & n868 ;
  assign n873 = ( x13 & n137 ) | ( x13 & n869 ) | ( n137 & n869 ) ;
  assign n870 = x4 & x6 ;
  assign n871 = ( x5 & n811 ) | ( x5 & n870 ) | ( n811 & n870 ) ;
  assign n872 = ~n811 & n871 ;
  assign n874 = ~x13 & n872 ;
  assign n875 = ( n869 & ~n873 ) | ( n869 & n874 ) | ( ~n873 & n874 ) ;
  assign n876 = x9 & n875 ;
  assign n877 = ( x10 & x12 ) | ( x10 & n876 ) | ( x12 & n876 ) ;
  assign n878 = ~x12 & n877 ;
  assign n923 = ~x2 & n878 ;
  assign n924 = x3 | n923 ;
  assign n925 = ~n922 & n924 ;
  assign n926 = x11 & n925 ;
  assign n865 = x6 | n213 ;
  assign n866 = ( ~x5 & x7 ) | ( ~x5 & n865 ) | ( x7 & n865 ) ;
  assign n867 = x5 | n866 ;
  assign n927 = n867 & ~n926 ;
  assign n928 = ( n864 & ~n926 ) | ( n864 & n927 ) | ( ~n926 & n927 ) ;
  assign n929 = x7 | n655 ;
  assign n930 = n862 | n929 ;
  assign n934 = x10 & ~x12 ;
  assign n935 = ~x13 & n934 ;
  assign n936 = n772 & n935 ;
  assign n937 = ( n213 & n761 ) | ( n213 & n936 ) | ( n761 & n936 ) ;
  assign n938 = ~n213 & n937 ;
  assign n939 = ( x0 & x9 ) | ( x0 & ~x10 ) | ( x9 & ~x10 ) ;
  assign n940 = ( x4 & ~x10 ) | ( x4 & n939 ) | ( ~x10 & n939 ) ;
  assign n941 = x10 & n940 ;
  assign n942 = n940 & ~n941 ;
  assign n943 = ( x10 & ~n941 ) | ( x10 & n942 ) | ( ~n941 & n942 ) ;
  assign n944 = x8 & ~x13 ;
  assign n945 = ( x12 & n943 ) | ( x12 & n944 ) | ( n943 & n944 ) ;
  assign n946 = ~n943 & n945 ;
  assign n947 = x2 & x7 ;
  assign n948 = ( x5 & ~n946 ) | ( x5 & n947 ) | ( ~n946 & n947 ) ;
  assign n949 = n946 & n948 ;
  assign n975 = ( x1 & x3 ) | ( x1 & ~n949 ) | ( x3 & ~n949 ) ;
  assign n950 = ( x13 & ~n87 ) | ( x13 & n692 ) | ( ~n87 & n692 ) ;
  assign n951 = n692 & ~n950 ;
  assign n972 = ( x2 & ~x12 ) | ( x2 & n951 ) | ( ~x12 & n951 ) ;
  assign n964 = x13 & n761 ;
  assign n965 = x10 & n964 ;
  assign n966 = ~x1 & x4 ;
  assign n967 = n965 & n966 ;
  assign n968 = ~n36 & n967 ;
  assign n957 = ~x9 & x13 ;
  assign n958 = ~x10 & n957 ;
  assign n959 = ~x1 & n87 ;
  assign n960 = n958 & n959 ;
  assign n961 = ( x1 & x13 ) | ( x1 & ~n960 ) | ( x13 & ~n960 ) ;
  assign n952 = ( x4 & x9 ) | ( x4 & ~x10 ) | ( x9 & ~x10 ) ;
  assign n953 = ( x5 & ~x10 ) | ( x5 & n952 ) | ( ~x10 & n952 ) ;
  assign n954 = x10 & n953 ;
  assign n955 = n953 & ~n954 ;
  assign n956 = ( x10 & ~n954 ) | ( x10 & n955 ) | ( ~n954 & n955 ) ;
  assign n962 = n956 & ~n960 ;
  assign n963 = ( ~x1 & n961 ) | ( ~x1 & n962 ) | ( n961 & n962 ) ;
  assign n969 = ( x7 & ~n963 ) | ( x7 & n968 ) | ( ~n963 & n968 ) ;
  assign n970 = x8 & ~n969 ;
  assign n971 = ( x8 & n968 ) | ( x8 & ~n970 ) | ( n968 & ~n970 ) ;
  assign n973 = ( x2 & x12 ) | ( x2 & ~n971 ) | ( x12 & ~n971 ) ;
  assign n974 = n972 & ~n973 ;
  assign n976 = x3 & n974 ;
  assign n977 = ( n949 & n975 ) | ( n949 & n976 ) | ( n975 & n976 ) ;
  assign n978 = ( x5 & ~n213 ) | ( x5 & n824 ) | ( ~n213 & n824 ) ;
  assign n979 = ~x5 & n978 ;
  assign n980 = x7 & n445 ;
  assign n981 = ( n935 & ~n979 ) | ( n935 & n980 ) | ( ~n979 & n980 ) ;
  assign n982 = n979 & n981 ;
  assign n983 = ( ~n938 & n977 ) | ( ~n938 & n982 ) | ( n977 & n982 ) ;
  assign n984 = x6 | n982 ;
  assign n985 = ( n938 & n983 ) | ( n938 & n984 ) | ( n983 & n984 ) ;
  assign n986 = x11 & n985 ;
  assign n931 = x5 | n213 ;
  assign n932 = ( ~x4 & x6 ) | ( ~x4 & n931 ) | ( x6 & n931 ) ;
  assign n933 = x4 | n932 ;
  assign n987 = n933 & ~n986 ;
  assign n988 = ( n930 & ~n986 ) | ( n930 & n987 ) | ( ~n986 & n987 ) ;
  assign n1072 = x8 & n539 ;
  assign n1073 = ~x5 & x7 ;
  assign n1074 = ~x6 & n1073 ;
  assign n1077 = ( x12 & n1072 ) | ( x12 & ~n1074 ) | ( n1072 & ~n1074 ) ;
  assign n1075 = ( x5 & ~n692 ) | ( x5 & n870 ) | ( ~n692 & n870 ) ;
  assign n1076 = n692 & n1075 ;
  assign n1078 = ~x12 & n1076 ;
  assign n1079 = ( n1072 & ~n1077 ) | ( n1072 & n1078 ) | ( ~n1077 & n1078 ) ;
  assign n1088 = ( x2 & ~x13 ) | ( x2 & n1079 ) | ( ~x13 & n1079 ) ;
  assign n1080 = x2 & ~n137 ;
  assign n1081 = ( x0 & x1 ) | ( x0 & n1080 ) | ( x1 & n1080 ) ;
  assign n1082 = ~x0 & n1081 ;
  assign n1083 = ~x9 & x12 ;
  assign n1084 = x10 & n1083 ;
  assign n1085 = x6 & ~n811 ;
  assign n1086 = ( ~n1082 & n1084 ) | ( ~n1082 & n1085 ) | ( n1084 & n1085 ) ;
  assign n1087 = n1082 & n1086 ;
  assign n1089 = ~x13 & n1087 ;
  assign n1090 = ( ~x2 & n1088 ) | ( ~x2 & n1089 ) | ( n1088 & n1089 ) ;
  assign n1091 = ~x3 & n1090 ;
  assign n1002 = x1 & ~x13 ;
  assign n1003 = x10 | x12 ;
  assign n1004 = ( x1 & ~n1002 ) | ( x1 & n1003 ) | ( ~n1002 & n1003 ) ;
  assign n1005 = x8 | n1004 ;
  assign n1006 = ( ~x6 & x9 ) | ( ~x6 & n1005 ) | ( x9 & n1005 ) ;
  assign n1007 = x6 | n1006 ;
  assign n1008 = x5 & x9 ;
  assign n1009 = ( x10 & x13 ) | ( x10 & n1008 ) | ( x13 & n1008 ) ;
  assign n1010 = ~x13 & n1009 ;
  assign n1011 = ( x1 & x5 ) | ( x1 & ~n1010 ) | ( x5 & ~n1010 ) ;
  assign n1012 = n958 & n1011 ;
  assign n1013 = ( n958 & n1010 ) | ( n958 & ~n1012 ) | ( n1010 & ~n1012 ) ;
  assign n1017 = ( ~x4 & x12 ) | ( ~x4 & n1013 ) | ( x12 & n1013 ) ;
  assign n1014 = x10 | n137 ;
  assign n1015 = ( ~x9 & x13 ) | ( ~x9 & n1014 ) | ( x13 & n1014 ) ;
  assign n1016 = x9 | n1015 ;
  assign n1018 = x12 | n1016 ;
  assign n1019 = ( ~n1013 & n1017 ) | ( ~n1013 & n1018 ) | ( n1017 & n1018 ) ;
  assign n1041 = ( x6 & x8 ) | ( x6 & n1019 ) | ( x8 & n1019 ) ;
  assign n990 = x6 & x9 ;
  assign n1029 = x10 & n990 ;
  assign n1030 = ( x4 & ~n32 ) | ( x4 & n1029 ) | ( ~n32 & n1029 ) ;
  assign n1031 = n32 & n1030 ;
  assign n1023 = x6 & n539 ;
  assign n1024 = x0 & ~x4 ;
  assign n1025 = x0 & ~n1024 ;
  assign n1026 = n1023 & n1025 ;
  assign n1020 = ( x6 & x9 ) | ( x6 & x10 ) | ( x9 & x10 ) ;
  assign n1021 = x6 & ~n1020 ;
  assign n1022 = ( x9 & ~n1020 ) | ( x9 & n1021 ) | ( ~n1020 & n1021 ) ;
  assign n1027 = ( n1022 & ~n1024 ) | ( n1022 & n1025 ) | ( ~n1024 & n1025 ) ;
  assign n1028 = ( ~x4 & n1026 ) | ( ~x4 & n1027 ) | ( n1026 & n1027 ) ;
  assign n1032 = ( ~x13 & n1028 ) | ( ~x13 & n1031 ) | ( n1028 & n1031 ) ;
  assign n1033 = x12 & ~n1032 ;
  assign n1034 = ( x12 & n1031 ) | ( x12 & ~n1033 ) | ( n1031 & ~n1033 ) ;
  assign n1038 = ( x1 & x5 ) | ( x1 & ~n1034 ) | ( x5 & ~n1034 ) ;
  assign n1035 = n32 & n258 ;
  assign n1036 = ( x4 & ~n72 ) | ( x4 & n1035 ) | ( ~n72 & n1035 ) ;
  assign n1037 = ~x4 & n1036 ;
  assign n1039 = x1 & n1037 ;
  assign n1040 = ( n1034 & n1038 ) | ( n1034 & n1039 ) | ( n1038 & n1039 ) ;
  assign n1042 = x8 & n1040 ;
  assign n1043 = ( ~n1019 & n1041 ) | ( ~n1019 & n1042 ) | ( n1041 & n1042 ) ;
  assign n1044 = ( x4 & x5 ) | ( x4 & ~n1043 ) | ( x5 & ~n1043 ) ;
  assign n1045 = ~n1007 & n1044 ;
  assign n1046 = ( n1007 & ~n1043 ) | ( n1007 & n1045 ) | ( ~n1043 & n1045 ) ;
  assign n1059 = ( x2 & x7 ) | ( x2 & n1046 ) | ( x7 & n1046 ) ;
  assign n1048 = ( x8 & x10 ) | ( x8 & n158 ) | ( x10 & n158 ) ;
  assign n1049 = ( x1 & x8 ) | ( x1 & ~n158 ) | ( x8 & ~n158 ) ;
  assign n1050 = ( x4 & x10 ) | ( x4 & n1049 ) | ( x10 & n1049 ) ;
  assign n1051 = ~n1048 & n1050 ;
  assign n1052 = x13 & ~n1051 ;
  assign n1047 = x4 | x8 ;
  assign n1053 = x10 & ~n1047 ;
  assign n1054 = x13 | n1053 ;
  assign n1055 = ~n1052 & n1054 ;
  assign n1056 = ( x12 & ~n434 ) | ( x12 & n1055 ) | ( ~n434 & n1055 ) ;
  assign n1057 = n1055 & ~n1056 ;
  assign n1058 = n258 & n1057 ;
  assign n1060 = x2 & n1058 ;
  assign n1061 = ( ~n1046 & n1059 ) | ( ~n1046 & n1060 ) | ( n1059 & n1060 ) ;
  assign n1062 = x7 & x9 ;
  assign n1063 = ( x8 & x10 ) | ( x8 & ~n1062 ) | ( x10 & ~n1062 ) ;
  assign n1064 = ( ~x7 & x8 ) | ( ~x7 & n1062 ) | ( x8 & n1062 ) ;
  assign n1065 = ( ~x9 & x10 ) | ( ~x9 & n1064 ) | ( x10 & n1064 ) ;
  assign n1066 = n1063 & ~n1065 ;
  assign n1067 = ( x13 & ~n333 ) | ( x13 & n1066 ) | ( ~n333 & n1066 ) ;
  assign n1068 = n1066 & ~n1067 ;
  assign n1069 = ~x5 & n1068 ;
  assign n1070 = ( x2 & x4 ) | ( x2 & n1069 ) | ( x4 & n1069 ) ;
  assign n1071 = ~x2 & n1070 ;
  assign n1092 = n1061 | n1071 ;
  assign n1093 = x3 & n1092 ;
  assign n1094 = n1091 | n1093 ;
  assign n1095 = x11 & n1094 ;
  assign n989 = x1 | x13 ;
  assign n991 = ( x1 & ~n989 ) | ( x1 & n990 ) | ( ~n989 & n990 ) ;
  assign n992 = ( x4 & n86 ) | ( x4 & ~n991 ) | ( n86 & ~n991 ) ;
  assign n993 = n991 & n992 ;
  assign n996 = ( ~x2 & x12 ) | ( ~x2 & n993 ) | ( x12 & n993 ) ;
  assign n994 = ( ~x5 & x13 ) | ( ~x5 & n865 ) | ( x13 & n865 ) ;
  assign n995 = x5 | n994 ;
  assign n997 = x12 | n995 ;
  assign n998 = ( ~n993 & n996 ) | ( ~n993 & n997 ) | ( n996 & n997 ) ;
  assign n999 = x10 | n998 ;
  assign n1000 = ( ~x8 & x11 ) | ( ~x8 & n999 ) | ( x11 & n999 ) ;
  assign n1001 = x8 | n1000 ;
  assign n1096 = n1001 & ~n1095 ;
  assign n1097 = ( x7 & ~n1095 ) | ( x7 & n1096 ) | ( ~n1095 & n1096 ) ;
  assign n1409 = ~x3 & n310 ;
  assign n1410 = ( x4 & ~x5 ) | ( x4 & n1409 ) | ( ~x5 & n1409 ) ;
  assign n1411 = ( n310 & n1409 ) | ( n310 & n1410 ) | ( n1409 & n1410 ) ;
  assign n1134 = x9 & n554 ;
  assign n1412 = n72 | n1134 ;
  assign n1413 = ( n868 & n1134 ) | ( n868 & ~n1412 ) | ( n1134 & ~n1412 ) ;
  assign n1420 = ~x6 & n1413 ;
  assign n1414 = x5 | n224 ;
  assign n1415 = x4 | n1414 ;
  assign n1417 = n67 & ~n811 ;
  assign n1322 = x6 | x7 ;
  assign n1416 = ( x6 & ~n460 ) | ( x6 & n1322 ) | ( ~n460 & n1322 ) ;
  assign n1418 = x0 & n1416 ;
  assign n1419 = ~n1417 & n1418 ;
  assign n1421 = n1415 & n1419 ;
  assign n1422 = ( ~n1413 & n1420 ) | ( ~n1413 & n1421 ) | ( n1420 & n1421 ) ;
  assign n1436 = x6 & n773 ;
  assign n1437 = ( x5 & n773 ) | ( x5 & n1436 ) | ( n773 & n1436 ) ;
  assign n1438 = ~x7 & n1437 ;
  assign n1423 = x5 & ~x11 ;
  assign n1424 = ( ~x5 & x9 ) | ( ~x5 & n1423 ) | ( x9 & n1423 ) ;
  assign n1425 = ( x9 & x10 ) | ( x9 & n1424 ) | ( x10 & n1424 ) ;
  assign n1426 = ( n72 & n1424 ) | ( n72 & ~n1425 ) | ( n1424 & ~n1425 ) ;
  assign n1433 = x3 & ~n1426 ;
  assign n1427 = n72 | n426 ;
  assign n1428 = ( n426 & ~n1134 ) | ( n426 & n1427 ) | ( ~n1134 & n1427 ) ;
  assign n1429 = ( x0 & ~n72 ) | ( x0 & n316 ) | ( ~n72 & n316 ) ;
  assign n1430 = ( ~x0 & n1134 ) | ( ~x0 & n1429 ) | ( n1134 & n1429 ) ;
  assign n1431 = x5 & ~n1430 ;
  assign n1432 = ( x5 & n1429 ) | ( x5 & ~n1431 ) | ( n1429 & ~n1431 ) ;
  assign n1434 = n1428 & ~n1432 ;
  assign n1435 = ( n1426 & n1433 ) | ( n1426 & n1434 ) | ( n1433 & n1434 ) ;
  assign n1439 = x6 & ~n1435 ;
  assign n1440 = x7 & ~n1439 ;
  assign n1441 = n1438 | n1440 ;
  assign n1533 = x8 | n1441 ;
  assign n1442 = ( x5 & ~x6 ) | ( x5 & x10 ) | ( ~x6 & x10 ) ;
  assign n1443 = x3 & n1442 ;
  assign n1444 = ( ~x3 & x5 ) | ( ~x3 & n1443 ) | ( x5 & n1443 ) ;
  assign n1449 = x0 & ~n1444 ;
  assign n1445 = x5 & x7 ;
  assign n1446 = x6 & n1445 ;
  assign n1447 = x8 & n554 ;
  assign n1448 = n1446 & n1447 ;
  assign n1450 = n110 & ~n1448 ;
  assign n1451 = ( n1444 & n1449 ) | ( n1444 & n1450 ) | ( n1449 & n1450 ) ;
  assign n1479 = ( ~x4 & x9 ) | ( ~x4 & n1451 ) | ( x9 & n1451 ) ;
  assign n1452 = x6 | n460 ;
  assign n1453 = x2 & ~x8 ;
  assign n1454 = ( x7 & n554 ) | ( x7 & n1453 ) | ( n554 & n1453 ) ;
  assign n1455 = ~x7 & n1454 ;
  assign n1456 = n1452 & ~n1455 ;
  assign n1457 = ( x0 & n1452 ) | ( x0 & ~n1456 ) | ( n1452 & ~n1456 ) ;
  assign n1458 = ( x0 & x3 ) | ( x0 & n1457 ) | ( x3 & n1457 ) ;
  assign n1459 = ( n37 & n1457 ) | ( n37 & ~n1458 ) | ( n1457 & ~n1458 ) ;
  assign n1476 = x5 & ~n1459 ;
  assign n1460 = x0 & x1 ;
  assign n1461 = ( x2 & x3 ) | ( x2 & n1460 ) | ( x3 & n1460 ) ;
  assign n1462 = ~x3 & n1461 ;
  assign n1463 = ( x0 & n868 ) | ( x0 & ~n1462 ) | ( n868 & ~n1462 ) ;
  assign n1464 = x3 & n1463 ;
  assign n1465 = ( x3 & n1462 ) | ( x3 & ~n1464 ) | ( n1462 & ~n1464 ) ;
  assign n1466 = ~x10 & n1465 ;
  assign n1467 = ( x5 & n1465 ) | ( x5 & n1466 ) | ( n1465 & n1466 ) ;
  assign n1468 = ( x3 & ~x5 ) | ( x3 & x10 ) | ( ~x5 & x10 ) ;
  assign n1469 = ( x5 & n224 ) | ( x5 & n1468 ) | ( n224 & n1468 ) ;
  assign n1470 = x3 | n1462 ;
  assign n1471 = ( ~x0 & n1462 ) | ( ~x0 & n1470 ) | ( n1462 & n1470 ) ;
  assign n1472 = ~x11 & n1471 ;
  assign n1473 = ( ~n1452 & n1471 ) | ( ~n1452 & n1472 ) | ( n1471 & n1472 ) ;
  assign n1474 = x0 & ~n1473 ;
  assign n1475 = ( n1469 & n1473 ) | ( n1469 & ~n1474 ) | ( n1473 & ~n1474 ) ;
  assign n1477 = n1467 | n1475 ;
  assign n1478 = ( n1459 & n1476 ) | ( n1459 & ~n1477 ) | ( n1476 & ~n1477 ) ;
  assign n1480 = x4 | n1478 ;
  assign n1481 = ( n1451 & ~n1479 ) | ( n1451 & n1480 ) | ( ~n1479 & n1480 ) ;
  assign n1098 = x1 & x2 ;
  assign n1482 = x0 & n1098 ;
  assign n1483 = n130 & n1482 ;
  assign n1484 = ( x5 & x9 ) | ( x5 & n1483 ) | ( x9 & n1483 ) ;
  assign n1485 = ~x9 & n1484 ;
  assign n1486 = ( x9 & ~x11 ) | ( x9 & n1485 ) | ( ~x11 & n1485 ) ;
  assign n1487 = n811 | n1486 ;
  assign n1488 = ( ~n811 & n1485 ) | ( ~n811 & n1487 ) | ( n1485 & n1487 ) ;
  assign n1530 = ~x10 & n1488 ;
  assign n1497 = ( ~x3 & x9 ) | ( ~x3 & n761 ) | ( x9 & n761 ) ;
  assign n1498 = x7 & ~n1497 ;
  assign n1499 = ~x7 & n110 ;
  assign n1500 = ( x10 & n1498 ) | ( x10 & ~n1499 ) | ( n1498 & ~n1499 ) ;
  assign n1501 = ( ~x7 & x10 ) | ( ~x7 & n1500 ) | ( x10 & n1500 ) ;
  assign n1496 = ( x5 & x11 ) | ( x5 & n67 ) | ( x11 & n67 ) ;
  assign n1502 = n1496 & n1500 ;
  assign n1503 = ( x7 & n1501 ) | ( x7 & n1502 ) | ( n1501 & n1502 ) ;
  assign n1504 = ( x7 & n460 ) | ( x7 & n1503 ) | ( n460 & n1503 ) ;
  assign n1505 = x2 & n1503 ;
  assign n1506 = ( ~n460 & n1504 ) | ( ~n460 & n1505 ) | ( n1504 & n1505 ) ;
  assign n1489 = n36 & ~n460 ;
  assign n1490 = x4 & ~n1489 ;
  assign n1491 = ( x0 & ~n1489 ) | ( x0 & n1490 ) | ( ~n1489 & n1490 ) ;
  assign n1492 = ( x4 & n86 ) | ( x4 & ~n1482 ) | ( n86 & ~n1482 ) ;
  assign n1493 = n1482 & n1492 ;
  assign n1494 = x7 | n460 ;
  assign n1495 = ( n460 & ~n1493 ) | ( n460 & n1494 ) | ( ~n1493 & n1494 ) ;
  assign n1507 = ( x6 & ~n1491 ) | ( x6 & n1495 ) | ( ~n1491 & n1495 ) ;
  assign n1508 = n1506 & ~n1507 ;
  assign n1509 = ( x6 & n1506 ) | ( x6 & ~n1508 ) | ( n1506 & ~n1508 ) ;
  assign n1516 = ~x8 & n67 ;
  assign n1517 = ~n36 & n1516 ;
  assign n1514 = ( x4 & n86 ) | ( x4 & n868 ) | ( n86 & n868 ) ;
  assign n1515 = ~n868 & n1514 ;
  assign n1518 = ( x1 & n1515 ) | ( x1 & n1517 ) | ( n1515 & n1517 ) ;
  assign n1519 = x2 & ~n1518 ;
  assign n1520 = ( x2 & n1517 ) | ( x2 & ~n1519 ) | ( n1517 & ~n1519 ) ;
  assign n1521 = x0 & n1520 ;
  assign n1510 = ( x3 & ~x5 ) | ( x3 & n295 ) | ( ~x5 & n295 ) ;
  assign n1511 = ~x3 & n1510 ;
  assign n1512 = ( ~x9 & n93 ) | ( ~x9 & n1511 ) | ( n93 & n1511 ) ;
  assign n1513 = ~n1511 & n1512 ;
  assign n1522 = n1513 | n1521 ;
  assign n1523 = ( ~x7 & n1521 ) | ( ~x7 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1524 = ( n1417 & ~n1493 ) | ( n1417 & n1523 ) | ( ~n1493 & n1523 ) ;
  assign n1525 = x10 & ~n1523 ;
  assign n1526 = ( n1493 & n1524 ) | ( n1493 & ~n1525 ) | ( n1524 & ~n1525 ) ;
  assign n1527 = ( n72 & n1493 ) | ( n72 & ~n1526 ) | ( n1493 & ~n1526 ) ;
  assign n1528 = x11 & ~n1526 ;
  assign n1529 = ( ~n1493 & n1527 ) | ( ~n1493 & n1528 ) | ( n1527 & n1528 ) ;
  assign n1531 = n1509 & n1529 ;
  assign n1532 = ( ~n1488 & n1530 ) | ( ~n1488 & n1531 ) | ( n1530 & n1531 ) ;
  assign n1534 = n1481 & n1532 ;
  assign n1535 = ( n1441 & ~n1533 ) | ( n1441 & n1534 ) | ( ~n1533 & n1534 ) ;
  assign n1536 = ( n1411 & n1422 ) | ( n1411 & n1535 ) | ( n1422 & n1535 ) ;
  assign n1537 = x1 & n1535 ;
  assign n1538 = ( ~n1411 & n1536 ) | ( ~n1411 & n1537 ) | ( n1536 & n1537 ) ;
  assign n1539 = x12 & ~n1538 ;
  assign n1226 = x6 & ~x8 ;
  assign n1227 = ( x4 & n426 ) | ( x4 & ~n1226 ) | ( n426 & ~n1226 ) ;
  assign n1228 = n1226 & n1227 ;
  assign n1229 = ( ~x6 & n70 ) | ( ~x6 & n1228 ) | ( n70 & n1228 ) ;
  assign n1230 = x7 & ~n1229 ;
  assign n1231 = ( x7 & n1228 ) | ( x7 & ~n1230 ) | ( n1228 & ~n1230 ) ;
  assign n1255 = ( x3 & x10 ) | ( x3 & ~n1231 ) | ( x10 & ~n1231 ) ;
  assign n1159 = x5 | x6 ;
  assign n1237 = x5 & n811 ;
  assign n1238 = ( ~x5 & n1159 ) | ( ~x5 & n1237 ) | ( n1159 & n1237 ) ;
  assign n1239 = ( x6 & x7 ) | ( x6 & x9 ) | ( x7 & x9 ) ;
  assign n1240 = ( x6 & ~x7 ) | ( x6 & x11 ) | ( ~x7 & x11 ) ;
  assign n1241 = n1239 | n1240 ;
  assign n1242 = ( ~x9 & n1239 ) | ( ~x9 & n1241 ) | ( n1239 & n1241 ) ;
  assign n1249 = ( ~x2 & x10 ) | ( ~x2 & n1242 ) | ( x10 & n1242 ) ;
  assign n1243 = x4 & n990 ;
  assign n1244 = x2 & n1243 ;
  assign n1245 = x9 & ~n1244 ;
  assign n1246 = ( x7 & n1244 ) | ( x7 & ~n1245 ) | ( n1244 & ~n1245 ) ;
  assign n1247 = x8 & n1246 ;
  assign n1248 = x5 & n1247 ;
  assign n1250 = ~x10 & n1248 ;
  assign n1251 = ( x2 & n1249 ) | ( x2 & ~n1250 ) | ( n1249 & ~n1250 ) ;
  assign n1252 = ( x2 & n1238 ) | ( x2 & n1251 ) | ( n1238 & n1251 ) ;
  assign n1200 = ( x7 & x9 ) | ( x7 & ~x11 ) | ( x9 & ~x11 ) ;
  assign n1232 = ( ~x7 & x8 ) | ( ~x7 & n1200 ) | ( x8 & n1200 ) ;
  assign n1233 = ( ~x8 & x11 ) | ( ~x8 & n1200 ) | ( x11 & n1200 ) ;
  assign n1234 = n1232 & n1233 ;
  assign n1235 = ( x5 & n870 ) | ( x5 & n1234 ) | ( n870 & n1234 ) ;
  assign n1236 = ~n1234 & n1235 ;
  assign n1253 = ( x2 & n1236 ) | ( x2 & ~n1251 ) | ( n1236 & ~n1251 ) ;
  assign n1254 = n1252 & ~n1253 ;
  assign n1256 = x3 & ~n1254 ;
  assign n1257 = ( n1231 & n1255 ) | ( n1231 & n1256 ) | ( n1255 & n1256 ) ;
  assign n1261 = x6 & n1134 ;
  assign n1262 = n868 & n1261 ;
  assign n1258 = ~x8 & n773 ;
  assign n1124 = x7 & n539 ;
  assign n1259 = x8 & ~n1124 ;
  assign n1260 = n1258 | n1259 ;
  assign n1263 = ( ~x2 & n1260 ) | ( ~x2 & n1262 ) | ( n1260 & n1262 ) ;
  assign n1264 = x6 | n1263 ;
  assign n1265 = ( ~x6 & n1262 ) | ( ~x6 & n1264 ) | ( n1262 & n1264 ) ;
  assign n1313 = x3 & ~x11 ;
  assign n1314 = ( x3 & ~x5 ) | ( x3 & n1313 ) | ( ~x5 & n1313 ) ;
  assign n1315 = x7 & n72 ;
  assign n1311 = x6 & ~x10 ;
  assign n1312 = ( ~x5 & x6 ) | ( ~x5 & n1311 ) | ( x6 & n1311 ) ;
  assign n1316 = x7 | n1312 ;
  assign n1317 = ( n1314 & n1315 ) | ( n1314 & n1316 ) | ( n1315 & n1316 ) ;
  assign n1363 = x8 & ~n1317 ;
  assign n1318 = x8 & ~x10 ;
  assign n1319 = ( n761 & ~n1062 ) | ( n761 & n1318 ) | ( ~n1062 & n1318 ) ;
  assign n1320 = ( x10 & n1318 ) | ( x10 & n1319 ) | ( n1318 & n1319 ) ;
  assign n1332 = x6 | n1320 ;
  assign n1321 = ( ~x7 & x8 ) | ( ~x7 & x9 ) | ( x8 & x9 ) ;
  assign n1323 = ( x9 & ~n1321 ) | ( x9 & n1322 ) | ( ~n1321 & n1322 ) ;
  assign n1324 = ( x9 & ~x10 ) | ( x9 & x11 ) | ( ~x10 & x11 ) ;
  assign n1325 = x8 & n1324 ;
  assign n1326 = ( ~x8 & x11 ) | ( ~x8 & n1325 ) | ( x11 & n1325 ) ;
  assign n1327 = ( x8 & ~x10 ) | ( x8 & n1326 ) | ( ~x10 & n1326 ) ;
  assign n1328 = x6 & n1326 ;
  assign n1329 = ( ~x8 & n1327 ) | ( ~x8 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = ~x9 & n1329 ;
  assign n1331 = ( n1226 & n1329 ) | ( n1226 & n1330 ) | ( n1329 & n1330 ) ;
  assign n1333 = n1323 & n1331 ;
  assign n1334 = ( n1320 & ~n1332 ) | ( n1320 & n1333 ) | ( ~n1332 & n1333 ) ;
  assign n1335 = ( ~x8 & x9 ) | ( ~x8 & n1334 ) | ( x9 & n1334 ) ;
  assign n1336 = x3 & n1334 ;
  assign n1337 = ( x8 & n1335 ) | ( x8 & n1336 ) | ( n1335 & n1336 ) ;
  assign n1348 = ( x4 & x5 ) | ( x4 & ~n1337 ) | ( x5 & ~n1337 ) ;
  assign n1340 = ( x10 & ~n445 ) | ( x10 & n773 ) | ( ~n445 & n773 ) ;
  assign n1342 = ( ~x7 & x8 ) | ( ~x7 & x11 ) | ( x8 & x11 ) ;
  assign n1341 = ( x4 & ~n72 ) | ( x4 & n771 ) | ( ~n72 & n771 ) ;
  assign n1343 = ~x8 & n1341 ;
  assign n1344 = ( x7 & n1342 ) | ( x7 & ~n1343 ) | ( n1342 & ~n1343 ) ;
  assign n1345 = ( x7 & n1340 ) | ( x7 & n1344 ) | ( n1340 & n1344 ) ;
  assign n1338 = x11 & ~n445 ;
  assign n1339 = ( n72 & ~n554 ) | ( n72 & n1338 ) | ( ~n554 & n1338 ) ;
  assign n1346 = ( ~x7 & n1339 ) | ( ~x7 & n1344 ) | ( n1339 & n1344 ) ;
  assign n1347 = n1345 & n1346 ;
  assign n1349 = x5 | n1347 ;
  assign n1350 = ( n1337 & n1348 ) | ( n1337 & n1349 ) | ( n1348 & n1349 ) ;
  assign n1353 = ( x4 & ~x9 ) | ( x4 & n1226 ) | ( ~x9 & n1226 ) ;
  assign n1180 = x5 & x8 ;
  assign n1351 = x11 & ~n1180 ;
  assign n1352 = ( x6 & ~n1180 ) | ( x6 & n1351 ) | ( ~n1180 & n1351 ) ;
  assign n1354 = x9 | n1352 ;
  assign n1355 = ( n1226 & ~n1353 ) | ( n1226 & n1354 ) | ( ~n1353 & n1354 ) ;
  assign n1356 = x7 & n1355 ;
  assign n1357 = x6 | n67 ;
  assign n1358 = ~x7 & n1357 ;
  assign n1359 = n1356 | n1358 ;
  assign n1360 = x10 | n1359 ;
  assign n1361 = ~n869 & n1360 ;
  assign n1362 = ( ~n1134 & n1360 ) | ( ~n1134 & n1361 ) | ( n1360 & n1361 ) ;
  assign n1364 = n1350 & n1362 ;
  assign n1365 = ( n1317 & n1363 ) | ( n1317 & n1364 ) | ( n1363 & n1364 ) ;
  assign n1366 = ( x4 & x6 ) | ( x4 & ~x11 ) | ( x6 & ~x11 ) ;
  assign n1367 = ( x5 & x6 ) | ( x5 & x11 ) | ( x6 & x11 ) ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1369 = x7 & x10 ;
  assign n1370 = ( x9 & ~n1368 ) | ( x9 & n1369 ) | ( ~n1368 & n1369 ) ;
  assign n1371 = n1368 & n1370 ;
  assign n1372 = x9 & ~n1062 ;
  assign n1373 = x6 & n1372 ;
  assign n1374 = ( x5 & n1062 ) | ( x5 & ~n1372 ) | ( n1062 & ~n1372 ) ;
  assign n1375 = ( x7 & n1373 ) | ( x7 & ~n1374 ) | ( n1373 & ~n1374 ) ;
  assign n1380 = ( x3 & x10 ) | ( x3 & n1375 ) | ( x10 & n1375 ) ;
  assign n1376 = ( x9 & ~x11 ) | ( x9 & n496 ) | ( ~x11 & n496 ) ;
  assign n1377 = ( n94 & n1062 ) | ( n94 & ~n1376 ) | ( n1062 & ~n1376 ) ;
  assign n1378 = x6 & n1377 ;
  assign n1379 = ( ~n881 & n1377 ) | ( ~n881 & n1378 ) | ( n1377 & n1378 ) ;
  assign n1381 = x10 | n1379 ;
  assign n1382 = ( ~n1375 & n1380 ) | ( ~n1375 & n1381 ) | ( n1380 & n1381 ) ;
  assign n1385 = ( x4 & ~x9 ) | ( x4 & n773 ) | ( ~x9 & n773 ) ;
  assign n1386 = ( x9 & n1047 ) | ( x9 & n1385 ) | ( n1047 & n1385 ) ;
  assign n1387 = ( x8 & ~n68 ) | ( x8 & n1386 ) | ( ~n68 & n1386 ) ;
  assign n1388 = x6 & n1386 ;
  assign n1389 = ( n68 & n1387 ) | ( n68 & n1388 ) | ( n1387 & n1388 ) ;
  assign n1392 = ( x6 & ~x8 ) | ( x6 & x10 ) | ( ~x8 & x10 ) ;
  assign n1390 = ( ~x3 & x9 ) | ( ~x3 & x10 ) | ( x9 & x10 ) ;
  assign n1391 = ( x3 & n1008 ) | ( x3 & n1390 ) | ( n1008 & n1390 ) ;
  assign n1393 = ( x6 & x8 ) | ( x6 & n1391 ) | ( x8 & n1391 ) ;
  assign n1394 = n1392 & ~n1393 ;
  assign n1395 = x5 | n1394 ;
  assign n1396 = ( ~n1389 & n1394 ) | ( ~n1389 & n1395 ) | ( n1394 & n1395 ) ;
  assign n1397 = x7 | n1396 ;
  assign n1383 = ~x10 & n1226 ;
  assign n1384 = ( ~x10 & n823 ) | ( ~x10 & n1383 ) | ( n823 & n1383 ) ;
  assign n1398 = ~x9 & n1384 ;
  assign n1399 = x7 & ~n1398 ;
  assign n1400 = n1397 & ~n1399 ;
  assign n1401 = ( n1371 & n1382 ) | ( n1371 & ~n1400 ) | ( n1382 & ~n1400 ) ;
  assign n1402 = x8 | n1400 ;
  assign n1403 = ( n1371 & ~n1401 ) | ( n1371 & n1402 ) | ( ~n1401 & n1402 ) ;
  assign n1404 = ( x2 & ~n1365 ) | ( x2 & n1403 ) | ( ~n1365 & n1403 ) ;
  assign n1266 = x7 & ~x8 ;
  assign n1267 = ( x8 & ~n69 ) | ( x8 & n1266 ) | ( ~n69 & n1266 ) ;
  assign n1308 = n586 | n1267 ;
  assign n1270 = ( x6 & x11 ) | ( x6 & ~n811 ) | ( x11 & ~n811 ) ;
  assign n1268 = x7 & n1072 ;
  assign n1269 = x5 & n1268 ;
  assign n1271 = x11 & n1269 ;
  assign n1272 = ( ~x6 & n1270 ) | ( ~x6 & n1271 ) | ( n1270 & n1271 ) ;
  assign n1273 = x3 | n539 ;
  assign n1274 = ( ~n87 & n539 ) | ( ~n87 & n1273 ) | ( n539 & n1273 ) ;
  assign n1275 = ( x3 & x4 ) | ( x3 & n110 ) | ( x4 & n110 ) ;
  assign n1276 = ( ~x4 & n554 ) | ( ~x4 & n1275 ) | ( n554 & n1275 ) ;
  assign n1277 = x7 & n1275 ;
  assign n1278 = ( x4 & n1276 ) | ( x4 & n1277 ) | ( n1276 & n1277 ) ;
  assign n1279 = x10 | n1062 ;
  assign n1280 = ( x8 & n1062 ) | ( x8 & n1279 ) | ( n1062 & n1279 ) ;
  assign n1281 = x4 & ~x11 ;
  assign n1282 = ( ~n15 & n1280 ) | ( ~n15 & n1281 ) | ( n1280 & n1281 ) ;
  assign n1286 = x5 & n1282 ;
  assign n1283 = ( x7 & n773 ) | ( x7 & ~n879 ) | ( n773 & ~n879 ) ;
  assign n1284 = x3 | x11 ;
  assign n1285 = ( x3 & ~n445 ) | ( x3 & n1284 ) | ( ~n445 & n1284 ) ;
  assign n1287 = n1283 & n1285 ;
  assign n1288 = ( ~n1282 & n1286 ) | ( ~n1282 & n1287 ) | ( n1286 & n1287 ) ;
  assign n1289 = ( ~n1274 & n1278 ) | ( ~n1274 & n1288 ) | ( n1278 & n1288 ) ;
  assign n1290 = x8 & n1288 ;
  assign n1291 = ( n1274 & n1289 ) | ( n1274 & n1290 ) | ( n1289 & n1290 ) ;
  assign n1305 = x6 | n1291 ;
  assign n1292 = ~x4 & n905 ;
  assign n1293 = ( x4 & ~x5 ) | ( x4 & n1292 ) | ( ~x5 & n1292 ) ;
  assign n1294 = ( x3 & n905 ) | ( x3 & ~n1293 ) | ( n905 & ~n1293 ) ;
  assign n1295 = ~n1292 & n1294 ;
  assign n1297 = ( x8 & ~x9 ) | ( x8 & n1295 ) | ( ~x9 & n1295 ) ;
  assign n1296 = ( ~x7 & n744 ) | ( ~x7 & n1062 ) | ( n744 & n1062 ) ;
  assign n1298 = x8 & n1296 ;
  assign n1299 = ( ~n1295 & n1297 ) | ( ~n1295 & n1298 ) | ( n1297 & n1298 ) ;
  assign n1301 = x7 & ~n863 ;
  assign n1300 = ( x6 & n445 ) | ( x6 & n870 ) | ( n445 & n870 ) ;
  assign n1302 = ( x3 & n1300 ) | ( x3 & ~n1301 ) | ( n1300 & ~n1301 ) ;
  assign n1303 = x5 & n1302 ;
  assign n1304 = ( x5 & n1301 ) | ( x5 & ~n1303 ) | ( n1301 & ~n1303 ) ;
  assign n1306 = n1299 | n1304 ;
  assign n1307 = ( ~n1291 & n1305 ) | ( ~n1291 & n1306 ) | ( n1305 & n1306 ) ;
  assign n1309 = n1272 | n1307 ;
  assign n1310 = ( ~n586 & n1308 ) | ( ~n586 & n1309 ) | ( n1308 & n1309 ) ;
  assign n1405 = ( ~x2 & n1310 ) | ( ~x2 & n1403 ) | ( n1310 & n1403 ) ;
  assign n1406 = n1404 | n1405 ;
  assign n1407 = n86 & ~n1406 ;
  assign n1408 = ( n1265 & n1406 ) | ( n1265 & ~n1407 ) | ( n1406 & ~n1407 ) ;
  assign n1540 = n1257 | n1408 ;
  assign n1541 = ~x12 & n1540 ;
  assign n1542 = n1539 | n1541 ;
  assign n1543 = x13 | n1542 ;
  assign n1106 = x7 & ~n158 ;
  assign n1099 = ( n583 & n773 ) | ( n583 & ~n1098 ) | ( n773 & ~n1098 ) ;
  assign n1100 = ~x7 & n773 ;
  assign n1101 = ( n1098 & n1099 ) | ( n1098 & n1100 ) | ( n1099 & n1100 ) ;
  assign n1103 = x6 & n736 ;
  assign n1102 = x2 & x3 ;
  assign n1104 = x1 & n1102 ;
  assign n1105 = n1103 & n1104 ;
  assign n1107 = n1101 | n1105 ;
  assign n1108 = ( n158 & n1106 ) | ( n158 & ~n1107 ) | ( n1106 & ~n1107 ) ;
  assign n1130 = ( x5 & ~x8 ) | ( x5 & n1108 ) | ( ~x8 & n1108 ) ;
  assign n1111 = ( x1 & x10 ) | ( x1 & x11 ) | ( x10 & x11 ) ;
  assign n1112 = ( ~x1 & n774 ) | ( ~x1 & n1111 ) | ( n774 & n1111 ) ;
  assign n1113 = ( ~x1 & x10 ) | ( ~x1 & x11 ) | ( x10 & x11 ) ;
  assign n1114 = ~x6 & x11 ;
  assign n1115 = ( x1 & n1113 ) | ( x1 & n1114 ) | ( n1113 & n1114 ) ;
  assign n1116 = x4 & ~n1115 ;
  assign n1117 = n990 & n1102 ;
  assign n1118 = ( n1115 & n1116 ) | ( n1115 & n1117 ) | ( n1116 & n1117 ) ;
  assign n1119 = x5 & n1118 ;
  assign n1120 = ( n1112 & n1118 ) | ( n1112 & n1119 ) | ( n1118 & n1119 ) ;
  assign n1121 = ( n495 & n966 ) | ( n495 & n1098 ) | ( n966 & n1098 ) ;
  assign n1122 = x3 & ~n1121 ;
  assign n1123 = ( x3 & n966 ) | ( x3 & ~n1122 ) | ( n966 & ~n1122 ) ;
  assign n1125 = ~x5 & n1123 ;
  assign n1126 = ( ~n539 & n1124 ) | ( ~n539 & n1125 ) | ( n1124 & n1125 ) ;
  assign n1127 = ( x7 & n1120 ) | ( x7 & ~n1126 ) | ( n1120 & ~n1126 ) ;
  assign n1109 = ~x10 & n139 ;
  assign n1110 = ~x9 & n1109 ;
  assign n1128 = ( x7 & n1110 ) | ( x7 & n1126 ) | ( n1110 & n1126 ) ;
  assign n1129 = n1127 & ~n1128 ;
  assign n1131 = x8 | n1129 ;
  assign n1132 = ( n1108 & ~n1130 ) | ( n1108 & n1131 ) | ( ~n1130 & n1131 ) ;
  assign n1145 = ( ~x7 & n761 ) | ( ~x7 & n773 ) | ( n761 & n773 ) ;
  assign n1141 = n966 | n1098 ;
  assign n1142 = ( n15 & n966 ) | ( n15 & n1141 ) | ( n966 & n1141 ) ;
  assign n1143 = x10 & n1142 ;
  assign n1144 = ~x5 & n1143 ;
  assign n1146 = ~n761 & n1144 ;
  assign n1147 = ( x7 & n1145 ) | ( x7 & ~n1146 ) | ( n1145 & ~n1146 ) ;
  assign n1135 = x8 & n1134 ;
  assign n1136 = x7 & ~n1135 ;
  assign n1137 = n1100 | n1136 ;
  assign n1133 = x5 & n636 ;
  assign n1138 = ( n130 & n1133 ) | ( n130 & n1137 ) | ( n1133 & n1137 ) ;
  assign n1139 = x2 & ~n1138 ;
  assign n1140 = ( x2 & n1137 ) | ( x2 & ~n1139 ) | ( n1137 & ~n1139 ) ;
  assign n1151 = ( ~x5 & x6 ) | ( ~x5 & x7 ) | ( x6 & x7 ) ;
  assign n1152 = ( x5 & x7 ) | ( x5 & ~n460 ) | ( x7 & ~n460 ) ;
  assign n1153 = n1151 | n1152 ;
  assign n1148 = ~x10 & n67 ;
  assign n1149 = ~x8 & n1148 ;
  assign n1150 = x3 & n1149 ;
  assign n1154 = ( x5 & n1150 ) | ( x5 & n1153 ) | ( n1150 & n1153 ) ;
  assign n1155 = ~x6 & n1154 ;
  assign n1156 = ( x6 & n1153 ) | ( x6 & n1155 ) | ( n1153 & n1155 ) ;
  assign n1157 = ( x5 & ~x6 ) | ( x5 & n23 ) | ( ~x6 & n23 ) ;
  assign n1158 = ( n22 & n23 ) | ( n22 & n1157 ) | ( n23 & n1157 ) ;
  assign n1161 = x10 & n881 ;
  assign n1160 = ( ~x3 & n112 ) | ( ~x3 & n1159 ) | ( n112 & n1159 ) ;
  assign n1162 = x1 & n1160 ;
  assign n1163 = ( ~n881 & n1161 ) | ( ~n881 & n1162 ) | ( n1161 & n1162 ) ;
  assign n1164 = ( x1 & n495 ) | ( x1 & n881 ) | ( n495 & n881 ) ;
  assign n1165 = ~x3 & n881 ;
  assign n1166 = ( ~x1 & n1164 ) | ( ~x1 & n1165 ) | ( n1164 & n1165 ) ;
  assign n1167 = ( x8 & x9 ) | ( x8 & n87 ) | ( x9 & n87 ) ;
  assign n1168 = ~x6 & x9 ;
  assign n1169 = ( ~n87 & n1167 ) | ( ~n87 & n1168 ) | ( n1167 & n1168 ) ;
  assign n1181 = ( x6 & ~n1102 ) | ( x6 & n1180 ) | ( ~n1102 & n1180 ) ;
  assign n1182 = n1102 & n1181 ;
  assign n1183 = ( x5 & x7 ) | ( x5 & ~n1182 ) | ( x7 & ~n1182 ) ;
  assign n1184 = x9 & n1183 ;
  assign n1185 = ( x9 & n1182 ) | ( x9 & ~n1184 ) | ( n1182 & ~n1184 ) ;
  assign n1187 = ( x1 & x4 ) | ( x1 & ~n1185 ) | ( x4 & ~n1185 ) ;
  assign n1186 = ~n36 & n445 ;
  assign n1188 = x1 & n1186 ;
  assign n1189 = ( n1185 & n1187 ) | ( n1185 & n1188 ) | ( n1187 & n1188 ) ;
  assign n1190 = ( ~x7 & n1169 ) | ( ~x7 & n1189 ) | ( n1169 & n1189 ) ;
  assign n1177 = ( x1 & ~x9 ) | ( x1 & n495 ) | ( ~x9 & n495 ) ;
  assign n1174 = x6 & n1047 ;
  assign n1170 = ( x1 & ~x4 ) | ( x1 & x8 ) | ( ~x4 & x8 ) ;
  assign n1171 = x4 | x11 ;
  assign n1172 = ( x1 & ~n1170 ) | ( x1 & n1171 ) | ( ~n1170 & n1171 ) ;
  assign n1173 = ~x5 & x11 ;
  assign n1175 = n1172 & n1173 ;
  assign n1176 = ( ~n1047 & n1174 ) | ( ~n1047 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1178 = x9 | n1176 ;
  assign n1179 = ( n495 & ~n1177 ) | ( n495 & n1178 ) | ( ~n1177 & n1178 ) ;
  assign n1191 = ( x7 & ~n1179 ) | ( x7 & n1189 ) | ( ~n1179 & n1189 ) ;
  assign n1192 = n1190 | n1191 ;
  assign n1202 = x1 & ~n632 ;
  assign n1203 = ( x4 & ~n632 ) | ( x4 & n1202 ) | ( ~n632 & n1202 ) ;
  assign n1201 = ( ~n880 & n1142 ) | ( ~n880 & n1200 ) | ( n1142 & n1200 ) ;
  assign n1204 = n445 & n1102 ;
  assign n1205 = ( x1 & x4 ) | ( x1 & n1204 ) | ( x4 & n1204 ) ;
  assign n1206 = ~x4 & n1205 ;
  assign n1207 = ( x1 & x3 ) | ( x1 & ~n1206 ) | ( x3 & ~n1206 ) ;
  assign n1208 = x4 & n1207 ;
  assign n1209 = ( x4 & n1206 ) | ( x4 & ~n1208 ) | ( n1206 & ~n1208 ) ;
  assign n1210 = n1201 | n1209 ;
  assign n1211 = n1203 | n1210 ;
  assign n1212 = ~x5 & n1211 ;
  assign n1193 = ( ~x7 & x9 ) | ( ~x7 & x11 ) | ( x9 & x11 ) ;
  assign n1194 = ( x7 & n761 ) | ( x7 & n1193 ) | ( n761 & n1193 ) ;
  assign n1195 = x6 & ~n1194 ;
  assign n1196 = x5 & n1195 ;
  assign n1197 = x2 & x4 ;
  assign n1198 = ( x3 & ~n1196 ) | ( x3 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1199 = n1196 & n1198 ;
  assign n1213 = n1199 | n1212 ;
  assign n1214 = ( x1 & n1212 ) | ( x1 & n1213 ) | ( n1212 & n1213 ) ;
  assign n1215 = ( ~n1166 & n1192 ) | ( ~n1166 & n1214 ) | ( n1192 & n1214 ) ;
  assign n1216 = x10 & ~n1214 ;
  assign n1217 = ( n1166 & n1215 ) | ( n1166 & ~n1216 ) | ( n1215 & ~n1216 ) ;
  assign n1218 = ( n1158 & n1163 ) | ( n1158 & ~n1217 ) | ( n1163 & ~n1217 ) ;
  assign n1219 = x2 & ~n1217 ;
  assign n1220 = ( ~n1158 & n1218 ) | ( ~n1158 & n1219 ) | ( n1218 & n1219 ) ;
  assign n1221 = n158 & n1220 ;
  assign n1222 = ( n1156 & n1220 ) | ( n1156 & n1221 ) | ( n1220 & n1221 ) ;
  assign n1223 = n1140 & n1222 ;
  assign n1224 = ( ~n1132 & n1147 ) | ( ~n1132 & n1223 ) | ( n1147 & n1223 ) ;
  assign n1225 = n1132 & n1224 ;
  assign n1544 = x12 | n1225 ;
  assign n1545 = x13 & n1544 ;
  assign n1546 = n1543 & ~n1545 ;
  assign y0 = n129 ;
  assign y1 = n207 ;
  assign y2 = n290 ;
  assign y3 = n386 ;
  assign y4 = n483 ;
  assign y5 = n550 ;
  assign y6 = n581 ;
  assign y7 = n654 ;
  assign y8 = ~n735 ;
  assign y9 = ~n860 ;
  assign y10 = ~n928 ;
  assign y11 = ~n988 ;
  assign y12 = ~n1097 ;
  assign y13 = n1546 ;
endmodule
