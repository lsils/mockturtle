module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 ;
  wire n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 ;
  assign n51 = x6 | x8 ;
  assign n52 = x7 | n51 ;
  assign n53 = x9 | n52 ;
  assign n54 = x10 & x11 ;
  assign n55 = ( x10 & x12 ) | ( x10 & n54 ) | ( x12 & n54 ) ;
  assign n56 = ~x1 & x2 ;
  assign n57 = x0 & n56 ;
  assign n58 = x0 & x2 ;
  assign n59 = x1 & n58 ;
  assign n60 = ~x34 & x35 ;
  assign n61 = x33 & n57 ;
  assign n62 = ( x34 & n60 ) | ( x34 & n61 ) | ( n60 & n61 ) ;
  assign n63 = x6 & x8 ;
  assign n64 = ( x6 & x7 ) | ( x6 & n63 ) | ( x7 & n63 ) ;
  assign n65 = n62 | n64 ;
  assign n66 = ( n59 & n62 ) | ( n59 & n65 ) | ( n62 & n65 ) ;
  assign n67 = x9 & ~x32 ;
  assign n68 = x10 & x33 ;
  assign n69 = x34 | n68 ;
  assign n70 = ( x11 & n68 ) | ( x11 & n69 ) | ( n68 & n69 ) ;
  assign n71 = x35 | n70 ;
  assign n72 = ( x12 & n70 ) | ( x12 & n71 ) | ( n70 & n71 ) ;
  assign n73 = x36 | n72 ;
  assign n74 = ( x13 & n72 ) | ( x13 & n73 ) | ( n72 & n73 ) ;
  assign n75 = x6 & x29 ;
  assign n76 = x30 | n75 ;
  assign n77 = ( x7 & n75 ) | ( x7 & n76 ) | ( n75 & n76 ) ;
  assign n78 = x31 | n77 ;
  assign n79 = ( x8 & n77 ) | ( x8 & n78 ) | ( n77 & n78 ) ;
  assign n80 = n74 | n79 ;
  assign n81 = ( x9 & ~n67 ) | ( x9 & n80 ) | ( ~n67 & n80 ) ;
  assign n82 = ( ~n59 & n66 ) | ( ~n59 & n81 ) | ( n66 & n81 ) ;
  assign n83 = n57 | n82 ;
  assign n84 = ( ~n57 & n66 ) | ( ~n57 & n83 ) | ( n66 & n83 ) ;
  assign n85 = ( x33 & x34 ) | ( x33 & x35 ) | ( x34 & x35 ) ;
  assign n86 = ( x33 & x34 ) | ( x33 & ~n85 ) | ( x34 & ~n85 ) ;
  assign n87 = ( x35 & ~n85 ) | ( x35 & n86 ) | ( ~n85 & n86 ) ;
  assign n88 = ~x36 & n87 ;
  assign n89 = x36 & ~n87 ;
  assign n90 = n88 | n89 ;
  assign n91 = ( x29 & x30 ) | ( x29 & x31 ) | ( x30 & x31 ) ;
  assign n92 = ( x29 & x30 ) | ( x29 & ~n91 ) | ( x30 & ~n91 ) ;
  assign n93 = ( x31 & ~n91 ) | ( x31 & n92 ) | ( ~n91 & n92 ) ;
  assign n94 = ~x32 & n93 ;
  assign n95 = x32 & ~n93 ;
  assign n96 = n94 | n95 ;
  assign n97 = ~n90 & n96 ;
  assign n98 = n90 & n96 ;
  assign n99 = ( n90 & n97 ) | ( n90 & ~n98 ) | ( n97 & ~n98 ) ;
  assign n100 = ( x10 & x11 ) | ( x10 & x12 ) | ( x11 & x12 ) ;
  assign n101 = ( x10 & x11 ) | ( x10 & ~n100 ) | ( x11 & ~n100 ) ;
  assign n102 = ( x12 & ~n100 ) | ( x12 & n101 ) | ( ~n100 & n101 ) ;
  assign n103 = ~x13 & n102 ;
  assign n104 = x13 & ~n102 ;
  assign n105 = n103 | n104 ;
  assign n106 = ( x6 & x7 ) | ( x6 & x8 ) | ( x7 & x8 ) ;
  assign n107 = ( x6 & x7 ) | ( x6 & ~n106 ) | ( x7 & ~n106 ) ;
  assign n108 = ( x8 & ~n106 ) | ( x8 & n107 ) | ( ~n106 & n107 ) ;
  assign n109 = ~x9 & n108 ;
  assign n110 = x9 & ~n108 ;
  assign n111 = n109 | n110 ;
  assign n112 = n105 | n111 ;
  assign n113 = n105 & ~n111 ;
  assign n114 = ( ~n105 & n112 ) | ( ~n105 & n113 ) | ( n112 & n113 ) ;
  assign n115 = x3 & ~x40 ;
  assign n116 = x34 & ~x48 ;
  assign n117 = x3 | n116 ;
  assign n118 = ~n115 & n117 ;
  assign n119 = ( ~x3 & x35 ) | ( ~x3 & n118 ) | ( x35 & n118 ) ;
  assign n120 = x48 & ~n119 ;
  assign n121 = ( x48 & n118 ) | ( x48 & ~n120 ) | ( n118 & ~n120 ) ;
  assign n122 = x3 & ~x4 ;
  assign n123 = x0 & x1 ;
  assign n124 = ( ~x3 & n122 ) | ( ~x3 & n123 ) | ( n122 & n123 ) ;
  assign n125 = ~x0 & x5 ;
  assign n126 = ~x4 & n125 ;
  assign n127 = ( ~x37 & n124 ) | ( ~x37 & n126 ) | ( n124 & n126 ) ;
  assign n128 = ( x36 & ~n124 ) | ( x36 & n126 ) | ( ~n124 & n126 ) ;
  assign n129 = ~n127 & n128 ;
  assign n130 = n124 | n129 ;
  assign n131 = ( n121 & n129 ) | ( n121 & n130 ) | ( n129 & n130 ) ;
  assign n132 = ~x0 & x2 ;
  assign n133 = x1 & n132 ;
  assign n134 = x13 & n133 ;
  assign n135 = x0 | x3 ;
  assign n136 = ( x0 & ~x2 ) | ( x0 & x3 ) | ( ~x2 & x3 ) ;
  assign n137 = ( x2 & n123 ) | ( x2 & n136 ) | ( n123 & n136 ) ;
  assign n138 = n133 | n137 ;
  assign n139 = x13 & ~n138 ;
  assign n140 = ( x0 & ~n135 ) | ( x0 & n139 ) | ( ~n135 & n139 ) ;
  assign n141 = x2 | x3 ;
  assign n142 = ( x11 & n137 ) | ( x11 & n141 ) | ( n137 & n141 ) ;
  assign n143 = x2 & ~x13 ;
  assign n144 = x3 & x38 ;
  assign n145 = x2 | n144 ;
  assign n146 = ~n143 & n145 ;
  assign n147 = n137 & n146 ;
  assign n148 = ( ~n141 & n142 ) | ( ~n141 & n147 ) | ( n142 & n147 ) ;
  assign n149 = n140 | n148 ;
  assign n150 = ( n133 & ~n134 ) | ( n133 & n149 ) | ( ~n134 & n149 ) ;
  assign n151 = ( x24 & ~n131 ) | ( x24 & n150 ) | ( ~n131 & n150 ) ;
  assign n152 = ( x25 & n131 ) | ( x25 & n150 ) | ( n131 & n150 ) ;
  assign n153 = n151 | n152 ;
  assign n154 = ( x22 & ~n131 ) | ( x22 & n150 ) | ( ~n131 & n150 ) ;
  assign n155 = ( x23 & n131 ) | ( x23 & n150 ) | ( n131 & n150 ) ;
  assign n156 = n154 & n155 ;
  assign n157 = n153 & ~n156 ;
  assign n158 = x3 & ~x13 ;
  assign n159 = x31 & ~x48 ;
  assign n160 = x3 | n159 ;
  assign n161 = ~n158 & n160 ;
  assign n162 = ( ~x3 & x32 ) | ( ~x3 & n161 ) | ( x32 & n161 ) ;
  assign n163 = x48 & ~n162 ;
  assign n164 = ( x48 & n161 ) | ( x48 & ~n163 ) | ( n161 & ~n163 ) ;
  assign n165 = ( x33 & ~n124 ) | ( x33 & n125 ) | ( ~n124 & n125 ) ;
  assign n166 = ( ~x37 & n124 ) | ( ~x37 & n125 ) | ( n124 & n125 ) ;
  assign n167 = n165 & ~n166 ;
  assign n168 = n124 | n167 ;
  assign n169 = ( n164 & n167 ) | ( n164 & n168 ) | ( n167 & n168 ) ;
  assign n170 = x10 & n133 ;
  assign n171 = x10 & ~n138 ;
  assign n172 = ( x0 & ~n135 ) | ( x0 & n171 ) | ( ~n135 & n171 ) ;
  assign n173 = ( x8 & n137 ) | ( x8 & n141 ) | ( n137 & n141 ) ;
  assign n174 = x10 | x12 ;
  assign n175 = x11 | n174 ;
  assign n176 = x2 & ~n175 ;
  assign n177 = x3 & x11 ;
  assign n178 = x2 | n177 ;
  assign n179 = ~n176 & n178 ;
  assign n180 = n137 & n179 ;
  assign n181 = ( ~n141 & n173 ) | ( ~n141 & n180 ) | ( n173 & n180 ) ;
  assign n182 = n172 | n181 ;
  assign n183 = ( n133 & ~n170 ) | ( n133 & n182 ) | ( ~n170 & n182 ) ;
  assign n184 = ( x24 & ~n169 ) | ( x24 & n183 ) | ( ~n169 & n183 ) ;
  assign n185 = ( x25 & n169 ) | ( x25 & n183 ) | ( n169 & n183 ) ;
  assign n186 = n184 | n185 ;
  assign n187 = ( x22 & ~n169 ) | ( x22 & n183 ) | ( ~n169 & n183 ) ;
  assign n188 = ( x23 & n169 ) | ( x23 & n183 ) | ( n169 & n183 ) ;
  assign n189 = n187 & n188 ;
  assign n190 = n186 & ~n189 ;
  assign n191 = x3 & ~x38 ;
  assign n192 = x32 & ~x48 ;
  assign n193 = x3 | n192 ;
  assign n194 = ~n191 & n193 ;
  assign n195 = ( ~x3 & x33 ) | ( ~x3 & n194 ) | ( x33 & n194 ) ;
  assign n196 = x48 & ~n195 ;
  assign n197 = ( x48 & n194 ) | ( x48 & ~n196 ) | ( n194 & ~n196 ) ;
  assign n198 = ( x34 & ~n124 ) | ( x34 & n126 ) | ( ~n124 & n126 ) ;
  assign n199 = ~n127 & n198 ;
  assign n200 = n124 | n199 ;
  assign n201 = ( n197 & n199 ) | ( n197 & n200 ) | ( n199 & n200 ) ;
  assign n202 = x11 & n133 ;
  assign n203 = x11 & ~n138 ;
  assign n204 = ( x0 & ~n135 ) | ( x0 & n203 ) | ( ~n135 & n203 ) ;
  assign n205 = ( x9 & n137 ) | ( x9 & n141 ) | ( n137 & n141 ) ;
  assign n206 = x11 & x12 ;
  assign n207 = ( x2 & ~x11 ) | ( x2 & x12 ) | ( ~x11 & x12 ) ;
  assign n208 = ~x3 & x12 ;
  assign n209 = ( x2 & x12 ) | ( x2 & n208 ) | ( x12 & n208 ) ;
  assign n210 = ( n206 & n207 ) | ( n206 & ~n209 ) | ( n207 & ~n209 ) ;
  assign n211 = n137 & n210 ;
  assign n212 = ( ~n141 & n205 ) | ( ~n141 & n211 ) | ( n205 & n211 ) ;
  assign n213 = n204 | n212 ;
  assign n214 = ( n133 & ~n202 ) | ( n133 & n213 ) | ( ~n202 & n213 ) ;
  assign n215 = ( x24 & ~n201 ) | ( x24 & n214 ) | ( ~n201 & n214 ) ;
  assign n216 = ( x25 & n201 ) | ( x25 & n214 ) | ( n201 & n214 ) ;
  assign n217 = n215 | n216 ;
  assign n218 = ( x22 & ~n201 ) | ( x22 & n214 ) | ( ~n201 & n214 ) ;
  assign n219 = ( x23 & n201 ) | ( x23 & n214 ) | ( n201 & n214 ) ;
  assign n220 = n218 & n219 ;
  assign n221 = n217 & ~n220 ;
  assign n222 = n190 & n221 ;
  assign n223 = x3 & ~x39 ;
  assign n224 = x33 & ~x48 ;
  assign n225 = x3 | n224 ;
  assign n226 = ~n223 & n225 ;
  assign n227 = ( ~x3 & x34 ) | ( ~x3 & n226 ) | ( x34 & n226 ) ;
  assign n228 = x48 & ~n227 ;
  assign n229 = ( x48 & n226 ) | ( x48 & ~n228 ) | ( n226 & ~n228 ) ;
  assign n230 = ( x35 & ~n124 ) | ( x35 & n126 ) | ( ~n124 & n126 ) ;
  assign n231 = ~n127 & n230 ;
  assign n232 = n124 | n231 ;
  assign n233 = ( n229 & n231 ) | ( n229 & n232 ) | ( n231 & n232 ) ;
  assign n234 = x12 & n133 ;
  assign n235 = x12 & ~n138 ;
  assign n236 = ( x0 & ~n135 ) | ( x0 & n235 ) | ( ~n135 & n235 ) ;
  assign n237 = ( x10 & n137 ) | ( x10 & n141 ) | ( n137 & n141 ) ;
  assign n238 = x2 & x12 ;
  assign n239 = x3 & x13 ;
  assign n240 = x2 | n239 ;
  assign n241 = ~n238 & n240 ;
  assign n242 = n137 & n241 ;
  assign n243 = ( ~n141 & n237 ) | ( ~n141 & n242 ) | ( n237 & n242 ) ;
  assign n244 = n236 | n243 ;
  assign n245 = ( n133 & ~n234 ) | ( n133 & n244 ) | ( ~n234 & n244 ) ;
  assign n246 = ( x24 & ~n233 ) | ( x24 & n245 ) | ( ~n233 & n245 ) ;
  assign n247 = ( x25 & n233 ) | ( x25 & n245 ) | ( n233 & n245 ) ;
  assign n248 = n246 | n247 ;
  assign n249 = ( x22 & ~n233 ) | ( x22 & n245 ) | ( ~n233 & n245 ) ;
  assign n250 = ( x23 & n233 ) | ( x23 & n245 ) | ( n233 & n245 ) ;
  assign n251 = n249 & n250 ;
  assign n252 = n248 & ~n251 ;
  assign n253 = n222 & n252 ;
  assign n254 = n157 & n253 ;
  assign n255 = x3 & ~x12 ;
  assign n256 = x30 & ~x48 ;
  assign n257 = x3 | n256 ;
  assign n258 = ~n255 & n257 ;
  assign n259 = ( ~x3 & x31 ) | ( ~x3 & n258 ) | ( x31 & n258 ) ;
  assign n260 = x48 & ~n259 ;
  assign n261 = ( x48 & n258 ) | ( x48 & ~n260 ) | ( n258 & ~n260 ) ;
  assign n262 = ( ~x0 & x4 ) | ( ~x0 & n125 ) | ( x4 & n125 ) ;
  assign n263 = ( ~x37 & n124 ) | ( ~x37 & n262 ) | ( n124 & n262 ) ;
  assign n264 = ( x32 & ~n124 ) | ( x32 & n262 ) | ( ~n124 & n262 ) ;
  assign n265 = ~n263 & n264 ;
  assign n266 = n124 | n265 ;
  assign n267 = ( n261 & n265 ) | ( n261 & n266 ) | ( n265 & n266 ) ;
  assign n268 = x9 & n133 ;
  assign n269 = x0 | x2 ;
  assign n270 = x9 & ~n138 ;
  assign n271 = ( x0 & ~n269 ) | ( x0 & n270 ) | ( ~n269 & n270 ) ;
  assign n272 = ( x7 & n137 ) | ( x7 & n141 ) | ( n137 & n141 ) ;
  assign n273 = x2 & ~x9 ;
  assign n274 = x3 & x10 ;
  assign n275 = x2 | n274 ;
  assign n276 = ~n273 & n275 ;
  assign n277 = n137 & n276 ;
  assign n278 = ( ~n141 & n272 ) | ( ~n141 & n277 ) | ( n272 & n277 ) ;
  assign n279 = n271 | n278 ;
  assign n280 = ( n133 & ~n268 ) | ( n133 & n279 ) | ( ~n268 & n279 ) ;
  assign n281 = ( x24 & ~n267 ) | ( x24 & n280 ) | ( ~n267 & n280 ) ;
  assign n282 = ( x25 & n267 ) | ( x25 & n280 ) | ( n267 & n280 ) ;
  assign n283 = n281 | n282 ;
  assign n284 = ( x22 & ~n267 ) | ( x22 & n280 ) | ( ~n267 & n280 ) ;
  assign n285 = ( x23 & n267 ) | ( x23 & n280 ) | ( n267 & n280 ) ;
  assign n286 = n284 & n285 ;
  assign n287 = n283 & ~n286 ;
  assign n288 = x3 & ~x9 ;
  assign n289 = x27 & ~x48 ;
  assign n290 = x3 | n289 ;
  assign n291 = ~n288 & n290 ;
  assign n292 = ( ~x3 & x28 ) | ( ~x3 & n291 ) | ( x28 & n291 ) ;
  assign n293 = x48 & ~n292 ;
  assign n294 = ( x48 & n291 ) | ( x48 & ~n293 ) | ( n291 & ~n293 ) ;
  assign n295 = ( x29 & ~n124 ) | ( x29 & n262 ) | ( ~n124 & n262 ) ;
  assign n296 = ~n263 & n295 ;
  assign n297 = n124 | n296 ;
  assign n298 = ( n294 & n296 ) | ( n294 & n297 ) | ( n296 & n297 ) ;
  assign n299 = x6 & n133 ;
  assign n300 = x6 & ~n138 ;
  assign n301 = ( x0 & ~n269 ) | ( x0 & n300 ) | ( ~n269 & n300 ) ;
  assign n302 = ( x20 & n137 ) | ( x20 & n141 ) | ( n137 & n141 ) ;
  assign n303 = x2 & ~n52 ;
  assign n304 = x3 & x7 ;
  assign n305 = x2 | n304 ;
  assign n306 = ~n303 & n305 ;
  assign n307 = n137 & n306 ;
  assign n308 = ( ~n141 & n302 ) | ( ~n141 & n307 ) | ( n302 & n307 ) ;
  assign n309 = n301 | n308 ;
  assign n310 = ( n133 & ~n299 ) | ( n133 & n309 ) | ( ~n299 & n309 ) ;
  assign n311 = ( x24 & ~n298 ) | ( x24 & n310 ) | ( ~n298 & n310 ) ;
  assign n312 = ( x25 & n298 ) | ( x25 & n310 ) | ( n298 & n310 ) ;
  assign n313 = n311 | n312 ;
  assign n314 = ( x22 & ~n298 ) | ( x22 & n310 ) | ( ~n298 & n310 ) ;
  assign n315 = ( x23 & n298 ) | ( x23 & n310 ) | ( n298 & n310 ) ;
  assign n316 = n314 & n315 ;
  assign n317 = n313 & ~n316 ;
  assign n318 = x3 & ~x10 ;
  assign n319 = x28 & ~x48 ;
  assign n320 = x3 | n319 ;
  assign n321 = ~n318 & n320 ;
  assign n322 = ( ~x3 & x29 ) | ( ~x3 & n321 ) | ( x29 & n321 ) ;
  assign n323 = x48 & ~n322 ;
  assign n324 = ( x48 & n321 ) | ( x48 & ~n323 ) | ( n321 & ~n323 ) ;
  assign n325 = ( x30 & ~n124 ) | ( x30 & n262 ) | ( ~n124 & n262 ) ;
  assign n326 = ~n263 & n325 ;
  assign n327 = n124 | n326 ;
  assign n328 = ( n324 & n326 ) | ( n324 & n327 ) | ( n326 & n327 ) ;
  assign n329 = x7 & n133 ;
  assign n330 = x7 & ~n138 ;
  assign n331 = ( x0 & ~n269 ) | ( x0 & n330 ) | ( ~n269 & n330 ) ;
  assign n332 = ( x21 & n137 ) | ( x21 & n141 ) | ( n137 & n141 ) ;
  assign n333 = x7 & x8 ;
  assign n334 = ( x2 & ~x7 ) | ( x2 & x8 ) | ( ~x7 & x8 ) ;
  assign n335 = ~x3 & x8 ;
  assign n336 = ( x2 & x8 ) | ( x2 & n335 ) | ( x8 & n335 ) ;
  assign n337 = ( n333 & n334 ) | ( n333 & ~n336 ) | ( n334 & ~n336 ) ;
  assign n338 = n137 & n337 ;
  assign n339 = ( ~n141 & n332 ) | ( ~n141 & n338 ) | ( n332 & n338 ) ;
  assign n340 = n331 | n339 ;
  assign n341 = ( n133 & ~n329 ) | ( n133 & n340 ) | ( ~n329 & n340 ) ;
  assign n342 = ( x24 & ~n328 ) | ( x24 & n341 ) | ( ~n328 & n341 ) ;
  assign n343 = ( x25 & n328 ) | ( x25 & n341 ) | ( n328 & n341 ) ;
  assign n344 = n342 | n343 ;
  assign n345 = ( x22 & ~n328 ) | ( x22 & n341 ) | ( ~n328 & n341 ) ;
  assign n346 = ( x23 & n328 ) | ( x23 & n341 ) | ( n328 & n341 ) ;
  assign n347 = n345 & n346 ;
  assign n348 = n344 & ~n347 ;
  assign n349 = n317 & n348 ;
  assign n350 = x3 & ~x11 ;
  assign n351 = x29 & ~x48 ;
  assign n352 = x3 | n351 ;
  assign n353 = ~n350 & n352 ;
  assign n354 = ( ~x3 & x30 ) | ( ~x3 & n353 ) | ( x30 & n353 ) ;
  assign n355 = x48 & ~n354 ;
  assign n356 = ( x48 & n353 ) | ( x48 & ~n355 ) | ( n353 & ~n355 ) ;
  assign n357 = ( x31 & ~n124 ) | ( x31 & n262 ) | ( ~n124 & n262 ) ;
  assign n358 = ~n263 & n357 ;
  assign n359 = n124 | n358 ;
  assign n360 = ( n356 & n358 ) | ( n356 & n359 ) | ( n358 & n359 ) ;
  assign n361 = x8 & n133 ;
  assign n362 = x8 & ~n138 ;
  assign n363 = ( x0 & ~n269 ) | ( x0 & n362 ) | ( ~n269 & n362 ) ;
  assign n364 = ( x6 & n137 ) | ( x6 & n141 ) | ( n137 & n141 ) ;
  assign n365 = x2 & x8 ;
  assign n366 = x3 & x9 ;
  assign n367 = x2 | n366 ;
  assign n368 = ~n365 & n367 ;
  assign n369 = n137 & n368 ;
  assign n370 = ( ~n141 & n364 ) | ( ~n141 & n369 ) | ( n364 & n369 ) ;
  assign n371 = n363 | n370 ;
  assign n372 = ( n133 & ~n361 ) | ( n133 & n371 ) | ( ~n361 & n371 ) ;
  assign n373 = ( x24 & ~n360 ) | ( x24 & n372 ) | ( ~n360 & n372 ) ;
  assign n374 = ( x25 & n360 ) | ( x25 & n372 ) | ( n360 & n372 ) ;
  assign n375 = n373 | n374 ;
  assign n376 = ( x22 & ~n360 ) | ( x22 & n372 ) | ( ~n360 & n372 ) ;
  assign n377 = ( x23 & n360 ) | ( x23 & n372 ) | ( n360 & n372 ) ;
  assign n378 = n376 & n377 ;
  assign n379 = n375 & ~n378 ;
  assign n380 = n349 & n379 ;
  assign n381 = n287 & n380 ;
  assign n382 = n254 & n381 ;
  assign n383 = n349 & ~n378 ;
  assign n384 = n317 & n379 ;
  assign n385 = ( ~n286 & n348 ) | ( ~n286 & n384 ) | ( n348 & n384 ) ;
  assign n386 = n286 & n385 ;
  assign n387 = n316 | n347 ;
  assign n388 = ( n313 & n316 ) | ( n313 & n387 ) | ( n316 & n387 ) ;
  assign n389 = n386 | n388 ;
  assign n390 = ( n349 & ~n383 ) | ( n349 & n389 ) | ( ~n383 & n389 ) ;
  assign n391 = n222 & ~n251 ;
  assign n392 = n190 & n252 ;
  assign n393 = ( ~n156 & n221 ) | ( ~n156 & n392 ) | ( n221 & n392 ) ;
  assign n394 = n156 & n393 ;
  assign n395 = n189 | n220 ;
  assign n396 = ( n186 & n189 ) | ( n186 & n395 ) | ( n189 & n395 ) ;
  assign n397 = n394 | n396 ;
  assign n398 = ( n222 & ~n391 ) | ( n222 & n397 ) | ( ~n391 & n397 ) ;
  assign n399 = n390 | n398 ;
  assign n400 = ( n381 & n390 ) | ( n381 & n399 ) | ( n390 & n399 ) ;
  assign n401 = ~x2 & x26 ;
  assign n402 = ( x0 & x1 ) | ( x0 & n401 ) | ( x1 & n401 ) ;
  assign n403 = ~x0 & n402 ;
  assign n404 = x47 & n403 ;
  assign n405 = n245 & ~n404 ;
  assign n406 = ( n245 & n252 ) | ( n245 & n405 ) | ( n252 & n405 ) ;
  assign n407 = ( ~n245 & n252 ) | ( ~n245 & n405 ) | ( n252 & n405 ) ;
  assign n408 = ( n245 & ~n406 ) | ( n245 & n407 ) | ( ~n406 & n407 ) ;
  assign n409 = n150 & ~n404 ;
  assign n410 = ( n150 & n157 ) | ( n150 & n409 ) | ( n157 & n409 ) ;
  assign n411 = ( ~n150 & n157 ) | ( ~n150 & n409 ) | ( n157 & n409 ) ;
  assign n412 = ( n150 & ~n410 ) | ( n150 & n411 ) | ( ~n410 & n411 ) ;
  assign n413 = n408 & n412 ;
  assign n414 = x46 & n413 ;
  assign n415 = ( n156 & n404 ) | ( n156 & ~n408 ) | ( n404 & ~n408 ) ;
  assign n416 = n251 & ~n404 ;
  assign n417 = ( n156 & ~n415 ) | ( n156 & n416 ) | ( ~n415 & n416 ) ;
  assign n418 = n414 | n417 ;
  assign n419 = x0 & ~x4 ;
  assign n420 = ( x1 & x2 ) | ( x1 & n419 ) | ( x2 & n419 ) ;
  assign n421 = ~x1 & n420 ;
  assign n422 = n169 | n233 ;
  assign n423 = n201 | n422 ;
  assign n424 = x23 & n131 ;
  assign n425 = x23 & ~n424 ;
  assign n426 = ~n423 & n425 ;
  assign n427 = n169 & n233 ;
  assign n428 = n201 & n427 ;
  assign n429 = ( ~n424 & n425 ) | ( ~n424 & n428 ) | ( n425 & n428 ) ;
  assign n430 = ( n131 & n426 ) | ( n131 & n429 ) | ( n426 & n429 ) ;
  assign n431 = n404 & ~n430 ;
  assign n432 = n254 & ~n404 ;
  assign n433 = ( n404 & ~n431 ) | ( n404 & n432 ) | ( ~n431 & n432 ) ;
  assign n434 = x46 & n433 ;
  assign n435 = n398 & ~n404 ;
  assign n436 = n434 | n435 ;
  assign n437 = ~x0 & n436 ;
  assign n438 = n64 | n437 ;
  assign n439 = ( n421 & n437 ) | ( n421 & n438 ) | ( n437 & n438 ) ;
  assign n440 = x13 | n175 ;
  assign n441 = ( n421 & ~n439 ) | ( n421 & n440 ) | ( ~n439 & n440 ) ;
  assign n442 = x0 & n441 ;
  assign n443 = ( x0 & n439 ) | ( x0 & ~n442 ) | ( n439 & ~n442 ) ;
  assign n444 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n445 = x5 & n444 ;
  assign n446 = ( x0 & ~x5 ) | ( x0 & n445 ) | ( ~x5 & n445 ) ;
  assign n447 = ~n421 & n446 ;
  assign n448 = x46 & ~n412 ;
  assign n449 = ( ~x46 & n412 ) | ( ~x46 & n447 ) | ( n412 & n447 ) ;
  assign n450 = ( ~n447 & n448 ) | ( ~n447 & n449 ) | ( n448 & n449 ) ;
  assign n451 = x2 & x22 ;
  assign n452 = ( ~x2 & n123 ) | ( ~x2 & n451 ) | ( n123 & n451 ) ;
  assign n453 = ( x1 & x2 ) | ( x1 & ~n452 ) | ( x2 & ~n452 ) ;
  assign n454 = ~x3 & n453 ;
  assign n455 = ( x3 & ~n452 ) | ( x3 & n454 ) | ( ~n452 & n454 ) ;
  assign n456 = ( x13 & ~n57 ) | ( x13 & n455 ) | ( ~n57 & n455 ) ;
  assign n457 = x5 & n111 ;
  assign n458 = ~x5 & n64 ;
  assign n459 = ( x5 & ~n457 ) | ( x5 & n458 ) | ( ~n457 & n458 ) ;
  assign n460 = ( x3 & ~n57 ) | ( x3 & n459 ) | ( ~n57 & n459 ) ;
  assign n461 = ( x3 & ~n55 ) | ( x3 & n57 ) | ( ~n55 & n57 ) ;
  assign n462 = ~n460 & n461 ;
  assign n463 = n455 & n462 ;
  assign n464 = ( ~x13 & n456 ) | ( ~x13 & n463 ) | ( n456 & n463 ) ;
  assign n465 = x23 & x25 ;
  assign n466 = ( ~x2 & x24 ) | ( ~x2 & n465 ) | ( x24 & n465 ) ;
  assign n467 = x2 & n466 ;
  assign n468 = ~x6 & n467 ;
  assign n469 = x2 & x23 ;
  assign n470 = ( x24 & x25 ) | ( x24 & n469 ) | ( x25 & n469 ) ;
  assign n471 = ~x25 & n470 ;
  assign n472 = ( x2 & x24 ) | ( x2 & n465 ) | ( x24 & n465 ) ;
  assign n473 = ~x24 & n472 ;
  assign n474 = x23 & ~x25 ;
  assign n475 = ( x2 & x24 ) | ( x2 & n474 ) | ( x24 & n474 ) ;
  assign n476 = ~x24 & n475 ;
  assign n477 = ~x9 & n476 ;
  assign n478 = x2 & x25 ;
  assign n479 = ( x23 & x24 ) | ( x23 & n478 ) | ( x24 & n478 ) ;
  assign n480 = ~x23 & n479 ;
  assign n481 = x10 & n480 ;
  assign n482 = ( x2 & x23 ) | ( x2 & x25 ) | ( x23 & x25 ) ;
  assign n483 = x24 & n482 ;
  assign n484 = ( x2 & ~x24 ) | ( x2 & n483 ) | ( ~x24 & n483 ) ;
  assign n485 = x2 & ~x24 ;
  assign n486 = ( x23 & ~x25 ) | ( x23 & n485 ) | ( ~x25 & n485 ) ;
  assign n487 = ~x23 & n486 ;
  assign n488 = x21 & n487 ;
  assign n489 = ~x24 & x25 ;
  assign n490 = ( x2 & x23 ) | ( x2 & n489 ) | ( x23 & n489 ) ;
  assign n491 = ~x23 & n490 ;
  assign n492 = n488 | n491 ;
  assign n493 = ( x12 & n488 ) | ( x12 & n492 ) | ( n488 & n492 ) ;
  assign n494 = x11 | n493 ;
  assign n495 = ( ~n484 & n493 ) | ( ~n484 & n494 ) | ( n493 & n494 ) ;
  assign n496 = n481 | n495 ;
  assign n497 = ( n476 & ~n477 ) | ( n476 & n496 ) | ( ~n477 & n496 ) ;
  assign n498 = x8 | n497 ;
  assign n499 = ( n473 & n497 ) | ( n473 & n498 ) | ( n497 & n498 ) ;
  assign n500 = x7 | n499 ;
  assign n501 = ( n471 & n499 ) | ( n471 & n500 ) | ( n499 & n500 ) ;
  assign n502 = x3 | n501 ;
  assign n503 = ( n467 & ~n468 ) | ( n467 & n502 ) | ( ~n468 & n502 ) ;
  assign n504 = ~x44 & n467 ;
  assign n505 = x45 & n487 ;
  assign n506 = n491 | n505 ;
  assign n507 = ( x38 & n505 ) | ( x38 & n506 ) | ( n505 & n506 ) ;
  assign n508 = x39 | n507 ;
  assign n509 = ( ~n484 & n507 ) | ( ~n484 & n508 ) | ( n507 & n508 ) ;
  assign n510 = x40 | n509 ;
  assign n511 = ( n480 & n509 ) | ( n480 & n510 ) | ( n509 & n510 ) ;
  assign n512 = x41 | n511 ;
  assign n513 = ( n476 & n511 ) | ( n476 & n512 ) | ( n511 & n512 ) ;
  assign n514 = x42 | n513 ;
  assign n515 = ( n473 & n513 ) | ( n473 & n514 ) | ( n513 & n514 ) ;
  assign n516 = x43 | n515 ;
  assign n517 = ( n471 & n515 ) | ( n471 & n516 ) | ( n515 & n516 ) ;
  assign n518 = x3 & ~n517 ;
  assign n519 = ( ~n467 & n504 ) | ( ~n467 & n518 ) | ( n504 & n518 ) ;
  assign n520 = x2 | n412 ;
  assign n521 = ( ~x1 & x3 ) | ( ~x1 & n520 ) | ( x3 & n520 ) ;
  assign n522 = x1 | n521 ;
  assign n523 = ( n503 & n519 ) | ( n503 & ~n522 ) | ( n519 & ~n522 ) ;
  assign n524 = ~n452 & n522 ;
  assign n525 = ( n503 & ~n523 ) | ( n503 & n524 ) | ( ~n523 & n524 ) ;
  assign n526 = ( n450 & ~n464 ) | ( n450 & n525 ) | ( ~n464 & n525 ) ;
  assign n527 = n447 & ~n526 ;
  assign n528 = ( n447 & n450 ) | ( n447 & ~n527 ) | ( n450 & ~n527 ) ;
  assign n529 = ~x1 & x3 ;
  assign n530 = x9 | n452 ;
  assign n531 = ( x1 & n529 ) | ( x1 & ~n530 ) | ( n529 & ~n530 ) ;
  assign n532 = n280 & ~n404 ;
  assign n533 = ( n280 & n287 ) | ( n280 & n532 ) | ( n287 & n532 ) ;
  assign n534 = ( ~n280 & n287 ) | ( ~n280 & n532 ) | ( n287 & n532 ) ;
  assign n535 = ( n280 & ~n533 ) | ( n280 & n534 ) | ( ~n533 & n534 ) ;
  assign n536 = x41 & n487 ;
  assign n537 = n491 | n536 ;
  assign n538 = ( x10 & n536 ) | ( x10 & n537 ) | ( n536 & n537 ) ;
  assign n539 = x11 | n538 ;
  assign n540 = ( ~n484 & n538 ) | ( ~n484 & n539 ) | ( n538 & n539 ) ;
  assign n541 = x12 | n540 ;
  assign n542 = ( n480 & n540 ) | ( n480 & n541 ) | ( n540 & n541 ) ;
  assign n543 = x13 | n542 ;
  assign n544 = ( n476 & n542 ) | ( n476 & n543 ) | ( n542 & n543 ) ;
  assign n545 = x38 | n544 ;
  assign n546 = ( n473 & n544 ) | ( n473 & n545 ) | ( n544 & n545 ) ;
  assign n547 = x39 | n546 ;
  assign n548 = ( n471 & n546 ) | ( n471 & n547 ) | ( n546 & n547 ) ;
  assign n549 = x40 | n548 ;
  assign n550 = ( n467 & n548 ) | ( n467 & n549 ) | ( n548 & n549 ) ;
  assign n551 = ( x3 & ~n452 ) | ( x3 & n550 ) | ( ~n452 & n550 ) ;
  assign n552 = x17 & n487 ;
  assign n553 = n491 | n552 ;
  assign n554 = ( x8 & n552 ) | ( x8 & n553 ) | ( n552 & n553 ) ;
  assign n555 = x7 | n554 ;
  assign n556 = ( ~n484 & n554 ) | ( ~n484 & n555 ) | ( n554 & n555 ) ;
  assign n557 = x6 | n556 ;
  assign n558 = ( n480 & n556 ) | ( n480 & n557 ) | ( n556 & n557 ) ;
  assign n559 = x21 | n558 ;
  assign n560 = ( n476 & n558 ) | ( n476 & n559 ) | ( n558 & n559 ) ;
  assign n561 = x20 | n560 ;
  assign n562 = ( n473 & n560 ) | ( n473 & n561 ) | ( n560 & n561 ) ;
  assign n563 = x19 | n562 ;
  assign n564 = ( n471 & n562 ) | ( n471 & n563 ) | ( n562 & n563 ) ;
  assign n565 = x18 | n564 ;
  assign n566 = ( n467 & n564 ) | ( n467 & n565 ) | ( n564 & n565 ) ;
  assign n567 = ( x3 & n452 ) | ( x3 & ~n566 ) | ( n452 & ~n566 ) ;
  assign n568 = ~n551 & n567 ;
  assign n569 = ( x1 & x3 ) | ( x1 & ~n568 ) | ( x3 & ~n568 ) ;
  assign n570 = ~n535 & n569 ;
  assign n571 = ( n535 & ~n568 ) | ( n535 & n570 ) | ( ~n568 & n570 ) ;
  assign n572 = ~n531 & n571 ;
  assign n573 = ( ~n434 & n435 ) | ( ~n434 & n535 ) | ( n435 & n535 ) ;
  assign n574 = ( n434 & ~n435 ) | ( n434 & n573 ) | ( ~n435 & n573 ) ;
  assign n575 = ( ~n535 & n573 ) | ( ~n535 & n574 ) | ( n573 & n574 ) ;
  assign n576 = n421 & n446 ;
  assign n577 = ( n446 & n575 ) | ( n446 & ~n576 ) | ( n575 & ~n576 ) ;
  assign n578 = ( n446 & n572 ) | ( n446 & ~n576 ) | ( n572 & ~n576 ) ;
  assign n579 = ( n572 & n577 ) | ( n572 & ~n578 ) | ( n577 & ~n578 ) ;
  assign n580 = ( x0 & ~x1 ) | ( x0 & n58 ) | ( ~x1 & n58 ) ;
  assign n581 = n381 | n390 ;
  assign n582 = ( n390 & n435 ) | ( n390 & n581 ) | ( n435 & n581 ) ;
  assign n583 = n435 & n535 ;
  assign n584 = n286 & ~n404 ;
  assign n585 = ~n583 & n584 ;
  assign n586 = n341 & ~n403 ;
  assign n587 = ( n341 & n348 ) | ( n341 & n586 ) | ( n348 & n586 ) ;
  assign n588 = ( ~n341 & n348 ) | ( ~n341 & n586 ) | ( n348 & n586 ) ;
  assign n589 = ( n341 & ~n587 ) | ( n341 & n588 ) | ( ~n587 & n588 ) ;
  assign n590 = n372 & ~n404 ;
  assign n591 = ( n372 & n379 ) | ( n372 & n590 ) | ( n379 & n590 ) ;
  assign n592 = ( ~n372 & n379 ) | ( ~n372 & n590 ) | ( n379 & n590 ) ;
  assign n593 = ( n372 & ~n591 ) | ( n372 & n592 ) | ( ~n591 & n592 ) ;
  assign n594 = n589 & n593 ;
  assign n595 = ( n583 & n585 ) | ( n583 & n594 ) | ( n585 & n594 ) ;
  assign n596 = n378 & ~n404 ;
  assign n597 = n589 & n596 ;
  assign n598 = n403 & ~n597 ;
  assign n599 = ( n347 & n597 ) | ( n347 & ~n598 ) | ( n597 & ~n598 ) ;
  assign n600 = n595 | n599 ;
  assign n601 = n535 & n589 ;
  assign n602 = ( ~n433 & n593 ) | ( ~n433 & n601 ) | ( n593 & n601 ) ;
  assign n603 = n433 & n602 ;
  assign n604 = n381 & n433 ;
  assign n605 = ( x46 & n603 ) | ( x46 & n604 ) | ( n603 & n604 ) ;
  assign n606 = ~n604 & n605 ;
  assign n607 = ( ~n603 & n605 ) | ( ~n603 & n606 ) | ( n605 & n606 ) ;
  assign n608 = ( n582 & ~n600 ) | ( n582 & n607 ) | ( ~n600 & n607 ) ;
  assign n609 = ( n582 & n600 ) | ( n582 & ~n607 ) | ( n600 & ~n607 ) ;
  assign n610 = ( ~n582 & n608 ) | ( ~n582 & n609 ) | ( n608 & n609 ) ;
  assign n611 = ~n580 & n610 ;
  assign n612 = ( x11 & x12 ) | ( x11 & n59 ) | ( x12 & n59 ) ;
  assign n613 = ( x11 & x12 ) | ( x11 & ~x13 ) | ( x12 & ~x13 ) ;
  assign n614 = n612 & ~n613 ;
  assign n615 = x6 & x7 ;
  assign n616 = x8 | n615 ;
  assign n617 = x6 & ~x9 ;
  assign n618 = ( x8 & n615 ) | ( x8 & n617 ) | ( n615 & n617 ) ;
  assign n619 = n616 & ~n618 ;
  assign n620 = ( ~x1 & n614 ) | ( ~x1 & n619 ) | ( n614 & n619 ) ;
  assign n621 = x0 & ~n620 ;
  assign n622 = ( x0 & n614 ) | ( x0 & ~n621 ) | ( n614 & ~n621 ) ;
  assign n623 = n611 | n622 ;
  assign n624 = n214 & ~n404 ;
  assign n625 = ( n214 & n221 ) | ( n214 & n624 ) | ( n221 & n624 ) ;
  assign n626 = ( ~n214 & n221 ) | ( ~n214 & n624 ) | ( n221 & n624 ) ;
  assign n627 = ( n214 & ~n625 ) | ( n214 & n626 ) | ( ~n625 & n626 ) ;
  assign n628 = ( n414 & n417 ) | ( n414 & ~n627 ) | ( n417 & ~n627 ) ;
  assign n629 = ( n414 & n417 ) | ( n414 & ~n628 ) | ( n417 & ~n628 ) ;
  assign n630 = ( n627 & n628 ) | ( n627 & ~n629 ) | ( n628 & ~n629 ) ;
  assign n631 = n156 & ~n404 ;
  assign n632 = x46 & n412 ;
  assign n633 = ( n408 & ~n631 ) | ( n408 & n632 ) | ( ~n631 & n632 ) ;
  assign n634 = ( n408 & n632 ) | ( n408 & ~n633 ) | ( n632 & ~n633 ) ;
  assign n635 = ( n631 & n633 ) | ( n631 & ~n634 ) | ( n633 & ~n634 ) ;
  assign n636 = n183 & ~n404 ;
  assign n637 = ( n183 & n190 ) | ( n183 & n636 ) | ( n190 & n636 ) ;
  assign n638 = ( ~n183 & n190 ) | ( ~n183 & n636 ) | ( n190 & n636 ) ;
  assign n639 = ( n183 & ~n637 ) | ( n183 & n638 ) | ( ~n637 & n638 ) ;
  assign n640 = x46 & n627 ;
  assign n641 = n413 & n640 ;
  assign n642 = ( n251 & n404 ) | ( n251 & ~n627 ) | ( n404 & ~n627 ) ;
  assign n643 = n220 & ~n404 ;
  assign n644 = ( n251 & ~n642 ) | ( n251 & n643 ) | ( ~n642 & n643 ) ;
  assign n645 = ( n408 & n627 ) | ( n408 & n644 ) | ( n627 & n644 ) ;
  assign n646 = n631 & ~n645 ;
  assign n647 = ( n631 & n644 ) | ( n631 & ~n646 ) | ( n644 & ~n646 ) ;
  assign n648 = ( ~n639 & n641 ) | ( ~n639 & n647 ) | ( n641 & n647 ) ;
  assign n649 = ( n641 & n647 ) | ( n641 & ~n648 ) | ( n647 & ~n648 ) ;
  assign n650 = ( n639 & n648 ) | ( n639 & ~n649 ) | ( n648 & ~n649 ) ;
  assign n651 = ( ~n630 & n635 ) | ( ~n630 & n650 ) | ( n635 & n650 ) ;
  assign n652 = n436 & n650 ;
  assign n653 = ( n630 & n651 ) | ( n630 & n652 ) | ( n651 & n652 ) ;
  assign n654 = ~n421 & n653 ;
  assign n655 = x10 | n57 ;
  assign n656 = x3 & ~n90 ;
  assign n657 = n57 & ~n656 ;
  assign n658 = n655 & ~n657 ;
  assign n659 = n455 & n658 ;
  assign n660 = ~x19 & n467 ;
  assign n661 = ~x7 & n480 ;
  assign n662 = x8 & ~n484 ;
  assign n663 = x18 & n487 ;
  assign n664 = n491 | n663 ;
  assign n665 = ( x9 & n663 ) | ( x9 & n664 ) | ( n663 & n664 ) ;
  assign n666 = n662 | n665 ;
  assign n667 = ( n480 & ~n661 ) | ( n480 & n666 ) | ( ~n661 & n666 ) ;
  assign n668 = x6 | n667 ;
  assign n669 = ( n476 & n667 ) | ( n476 & n668 ) | ( n667 & n668 ) ;
  assign n670 = x21 | n669 ;
  assign n671 = ( n473 & n669 ) | ( n473 & n670 ) | ( n669 & n670 ) ;
  assign n672 = x20 | n671 ;
  assign n673 = ( n471 & n671 ) | ( n471 & n672 ) | ( n671 & n672 ) ;
  assign n674 = x3 | n673 ;
  assign n675 = ( n467 & ~n660 ) | ( n467 & n674 ) | ( ~n660 & n674 ) ;
  assign n676 = ~x41 & n467 ;
  assign n677 = x42 & n487 ;
  assign n678 = n491 | n677 ;
  assign n679 = ( x11 & n677 ) | ( x11 & n678 ) | ( n677 & n678 ) ;
  assign n680 = x12 | n679 ;
  assign n681 = ( ~n484 & n679 ) | ( ~n484 & n680 ) | ( n679 & n680 ) ;
  assign n682 = x13 | n681 ;
  assign n683 = ( n480 & n681 ) | ( n480 & n682 ) | ( n681 & n682 ) ;
  assign n684 = x38 | n683 ;
  assign n685 = ( n476 & n683 ) | ( n476 & n684 ) | ( n683 & n684 ) ;
  assign n686 = x39 | n685 ;
  assign n687 = ( n473 & n685 ) | ( n473 & n686 ) | ( n685 & n686 ) ;
  assign n688 = x40 | n687 ;
  assign n689 = ( n471 & n687 ) | ( n471 & n688 ) | ( n687 & n688 ) ;
  assign n690 = x3 & ~n689 ;
  assign n691 = ( ~n467 & n676 ) | ( ~n467 & n690 ) | ( n676 & n690 ) ;
  assign n692 = x2 | n639 ;
  assign n693 = ( ~x1 & x3 ) | ( ~x1 & n692 ) | ( x3 & n692 ) ;
  assign n694 = x1 | n693 ;
  assign n695 = ( n675 & n691 ) | ( n675 & ~n694 ) | ( n691 & ~n694 ) ;
  assign n696 = ~n452 & n694 ;
  assign n697 = ( n675 & ~n695 ) | ( n675 & n696 ) | ( ~n695 & n696 ) ;
  assign n698 = n447 & n697 ;
  assign n699 = ( ~n455 & n659 ) | ( ~n455 & n698 ) | ( n659 & n698 ) ;
  assign n700 = ~n446 & n650 ;
  assign n701 = n699 | n700 ;
  assign n702 = ( n653 & ~n654 ) | ( n653 & n701 ) | ( ~n654 & n701 ) ;
  assign n703 = ~n446 & n635 ;
  assign n704 = ~n436 & n635 ;
  assign n705 = ( n421 & ~n436 ) | ( n421 & n635 ) | ( ~n436 & n635 ) ;
  assign n706 = ( n703 & ~n704 ) | ( n703 & n705 ) | ( ~n704 & n705 ) ;
  assign n707 = ( x12 & ~n57 ) | ( x12 & n455 ) | ( ~n57 & n455 ) ;
  assign n708 = x5 & n96 ;
  assign n709 = x8 & ~x9 ;
  assign n710 = x6 | n440 ;
  assign n711 = ( x8 & ~n709 ) | ( x8 & n710 ) | ( ~n709 & n710 ) ;
  assign n712 = x7 & ~n711 ;
  assign n713 = x5 | n712 ;
  assign n714 = ~n708 & n713 ;
  assign n715 = ( x3 & ~n57 ) | ( x3 & n714 ) | ( ~n57 & n714 ) ;
  assign n716 = ( x3 & n57 ) | ( x3 & n440 ) | ( n57 & n440 ) ;
  assign n717 = ~n715 & n716 ;
  assign n718 = n455 & n717 ;
  assign n719 = ( ~x12 & n707 ) | ( ~x12 & n718 ) | ( n707 & n718 ) ;
  assign n720 = ~x21 & n467 ;
  assign n721 = ~x8 & n476 ;
  assign n722 = x9 & n480 ;
  assign n723 = x20 & n487 ;
  assign n724 = n491 | n723 ;
  assign n725 = ( x11 & n723 ) | ( x11 & n724 ) | ( n723 & n724 ) ;
  assign n726 = x10 | n725 ;
  assign n727 = ( ~n484 & n725 ) | ( ~n484 & n726 ) | ( n725 & n726 ) ;
  assign n728 = n722 | n727 ;
  assign n729 = ( n476 & ~n721 ) | ( n476 & n728 ) | ( ~n721 & n728 ) ;
  assign n730 = x7 | n729 ;
  assign n731 = ( n473 & n729 ) | ( n473 & n730 ) | ( n729 & n730 ) ;
  assign n732 = x6 | n731 ;
  assign n733 = ( n471 & n731 ) | ( n471 & n732 ) | ( n731 & n732 ) ;
  assign n734 = x3 | n733 ;
  assign n735 = ( n467 & ~n720 ) | ( n467 & n734 ) | ( ~n720 & n734 ) ;
  assign n736 = ~x43 & n467 ;
  assign n737 = x44 & n487 ;
  assign n738 = n491 | n737 ;
  assign n739 = ( x13 & n737 ) | ( x13 & n738 ) | ( n737 & n738 ) ;
  assign n740 = x38 | n739 ;
  assign n741 = ( ~n484 & n739 ) | ( ~n484 & n740 ) | ( n739 & n740 ) ;
  assign n742 = x39 | n741 ;
  assign n743 = ( n480 & n741 ) | ( n480 & n742 ) | ( n741 & n742 ) ;
  assign n744 = x40 | n743 ;
  assign n745 = ( n476 & n743 ) | ( n476 & n744 ) | ( n743 & n744 ) ;
  assign n746 = x41 | n745 ;
  assign n747 = ( n473 & n745 ) | ( n473 & n746 ) | ( n745 & n746 ) ;
  assign n748 = x42 | n747 ;
  assign n749 = ( n471 & n747 ) | ( n471 & n748 ) | ( n747 & n748 ) ;
  assign n750 = x3 & ~n749 ;
  assign n751 = ( ~n467 & n736 ) | ( ~n467 & n750 ) | ( n736 & n750 ) ;
  assign n752 = x2 | n408 ;
  assign n753 = ( ~x1 & x3 ) | ( ~x1 & n752 ) | ( x3 & n752 ) ;
  assign n754 = x1 | n753 ;
  assign n755 = ( n735 & n751 ) | ( n735 & ~n754 ) | ( n751 & ~n754 ) ;
  assign n756 = ~n452 & n754 ;
  assign n757 = ( n735 & ~n755 ) | ( n735 & n756 ) | ( ~n755 & n756 ) ;
  assign n758 = ( n706 & ~n719 ) | ( n706 & n757 ) | ( ~n719 & n757 ) ;
  assign n759 = n447 & ~n758 ;
  assign n760 = ( n447 & n706 ) | ( n447 & ~n759 ) | ( n706 & ~n759 ) ;
  assign n761 = n446 & n630 ;
  assign n762 = x11 | n57 ;
  assign n763 = x3 & ~n105 ;
  assign n764 = n57 & ~n763 ;
  assign n765 = n762 & ~n764 ;
  assign n766 = n455 & n765 ;
  assign n767 = ~x20 & n467 ;
  assign n768 = ~x8 & n480 ;
  assign n769 = x9 & ~n484 ;
  assign n770 = x19 & n487 ;
  assign n771 = n491 | n770 ;
  assign n772 = ( x10 & n770 ) | ( x10 & n771 ) | ( n770 & n771 ) ;
  assign n773 = n769 | n772 ;
  assign n774 = ( n480 & ~n768 ) | ( n480 & n773 ) | ( ~n768 & n773 ) ;
  assign n775 = x7 | n774 ;
  assign n776 = ( n476 & n774 ) | ( n476 & n775 ) | ( n774 & n775 ) ;
  assign n777 = x6 | n776 ;
  assign n778 = ( n473 & n776 ) | ( n473 & n777 ) | ( n776 & n777 ) ;
  assign n779 = x21 | n778 ;
  assign n780 = ( n471 & n778 ) | ( n471 & n779 ) | ( n778 & n779 ) ;
  assign n781 = x3 | n780 ;
  assign n782 = ( n467 & ~n767 ) | ( n467 & n781 ) | ( ~n767 & n781 ) ;
  assign n783 = ~x42 & n467 ;
  assign n784 = x43 & n487 ;
  assign n785 = n491 | n784 ;
  assign n786 = ( x12 & n784 ) | ( x12 & n785 ) | ( n784 & n785 ) ;
  assign n787 = x13 | n786 ;
  assign n788 = ( ~n484 & n786 ) | ( ~n484 & n787 ) | ( n786 & n787 ) ;
  assign n789 = x38 | n788 ;
  assign n790 = ( n480 & n788 ) | ( n480 & n789 ) | ( n788 & n789 ) ;
  assign n791 = x39 | n790 ;
  assign n792 = ( n476 & n790 ) | ( n476 & n791 ) | ( n790 & n791 ) ;
  assign n793 = x40 | n792 ;
  assign n794 = ( n473 & n792 ) | ( n473 & n793 ) | ( n792 & n793 ) ;
  assign n795 = x41 | n794 ;
  assign n796 = ( n471 & n794 ) | ( n471 & n795 ) | ( n794 & n795 ) ;
  assign n797 = x3 & ~n796 ;
  assign n798 = ( ~n467 & n783 ) | ( ~n467 & n797 ) | ( n783 & n797 ) ;
  assign n799 = x2 | n627 ;
  assign n800 = ( ~x1 & x3 ) | ( ~x1 & n799 ) | ( x3 & n799 ) ;
  assign n801 = x1 | n800 ;
  assign n802 = ( n782 & n798 ) | ( n782 & ~n801 ) | ( n798 & ~n801 ) ;
  assign n803 = ~n452 & n801 ;
  assign n804 = ( n782 & ~n802 ) | ( n782 & n803 ) | ( ~n802 & n803 ) ;
  assign n805 = n447 & n804 ;
  assign n806 = ( ~n455 & n766 ) | ( ~n455 & n805 ) | ( n766 & n805 ) ;
  assign n807 = ( n421 & n436 ) | ( n421 & ~n635 ) | ( n436 & ~n635 ) ;
  assign n808 = n630 | n807 ;
  assign n809 = ( ~n421 & n630 ) | ( ~n421 & n807 ) | ( n630 & n807 ) ;
  assign n810 = ( n421 & ~n808 ) | ( n421 & n809 ) | ( ~n808 & n809 ) ;
  assign n811 = n806 | n810 ;
  assign n812 = ( n630 & ~n761 ) | ( n630 & n811 ) | ( ~n761 & n811 ) ;
  assign n813 = x39 & n487 ;
  assign n814 = n491 | n813 ;
  assign n815 = ( x8 & n813 ) | ( x8 & n814 ) | ( n813 & n814 ) ;
  assign n816 = n481 | n815 ;
  assign n817 = n769 | n816 ;
  assign n818 = x11 | n817 ;
  assign n819 = ( n476 & n817 ) | ( n476 & n818 ) | ( n817 & n818 ) ;
  assign n820 = x12 | n819 ;
  assign n821 = ( n473 & n819 ) | ( n473 & n820 ) | ( n819 & n820 ) ;
  assign n822 = x13 | n821 ;
  assign n823 = ( n471 & n821 ) | ( n471 & n822 ) | ( n821 & n822 ) ;
  assign n824 = x38 | n823 ;
  assign n825 = ( n467 & n823 ) | ( n467 & n824 ) | ( n823 & n824 ) ;
  assign n826 = ( x3 & ~n452 ) | ( x3 & n825 ) | ( ~n452 & n825 ) ;
  assign n827 = x15 & n487 ;
  assign n828 = n491 | n827 ;
  assign n829 = ( x6 & n827 ) | ( x6 & n828 ) | ( n827 & n828 ) ;
  assign n830 = x21 | n829 ;
  assign n831 = ( ~n484 & n829 ) | ( ~n484 & n830 ) | ( n829 & n830 ) ;
  assign n832 = x20 | n831 ;
  assign n833 = ( n480 & n831 ) | ( n480 & n832 ) | ( n831 & n832 ) ;
  assign n834 = x19 | n833 ;
  assign n835 = ( n476 & n833 ) | ( n476 & n834 ) | ( n833 & n834 ) ;
  assign n836 = x18 | n835 ;
  assign n837 = ( n473 & n835 ) | ( n473 & n836 ) | ( n835 & n836 ) ;
  assign n838 = x17 | n837 ;
  assign n839 = ( n471 & n837 ) | ( n471 & n838 ) | ( n837 & n838 ) ;
  assign n840 = x16 | n839 ;
  assign n841 = ( n467 & n839 ) | ( n467 & n840 ) | ( n839 & n840 ) ;
  assign n842 = ( x3 & n452 ) | ( x3 & ~n841 ) | ( n452 & ~n841 ) ;
  assign n843 = ~n826 & n842 ;
  assign n844 = ( x1 & x3 ) | ( x1 & ~n843 ) | ( x3 & ~n843 ) ;
  assign n845 = ~n589 & n844 ;
  assign n846 = ( n589 & ~n843 ) | ( n589 & n845 ) | ( ~n843 & n845 ) ;
  assign n847 = n433 & n535 ;
  assign n848 = x46 & n593 ;
  assign n849 = n847 & n848 ;
  assign n850 = n584 | n596 ;
  assign n851 = ( n593 & n596 ) | ( n593 & n850 ) | ( n596 & n850 ) ;
  assign n852 = ( n535 & n593 ) | ( n535 & n851 ) | ( n593 & n851 ) ;
  assign n853 = n435 & ~n852 ;
  assign n854 = ( n435 & n851 ) | ( n435 & ~n853 ) | ( n851 & ~n853 ) ;
  assign n855 = ( ~n589 & n849 ) | ( ~n589 & n854 ) | ( n849 & n854 ) ;
  assign n856 = ( n849 & n854 ) | ( n849 & ~n855 ) | ( n854 & ~n855 ) ;
  assign n857 = ( n589 & n855 ) | ( n589 & ~n856 ) | ( n855 & ~n856 ) ;
  assign n858 = ~n446 & n857 ;
  assign n859 = ( n583 & ~n585 ) | ( n583 & n593 ) | ( ~n585 & n593 ) ;
  assign n860 = ( n583 & n585 ) | ( n583 & ~n593 ) | ( n585 & ~n593 ) ;
  assign n861 = ( ~n583 & n859 ) | ( ~n583 & n860 ) | ( n859 & n860 ) ;
  assign n862 = ~x46 & n847 ;
  assign n863 = ( n847 & ~n861 ) | ( n847 & n862 ) | ( ~n861 & n862 ) ;
  assign n864 = ( n847 & n861 ) | ( n847 & ~n862 ) | ( n861 & ~n862 ) ;
  assign n865 = ( ~n847 & n863 ) | ( ~n847 & n864 ) | ( n863 & n864 ) ;
  assign n866 = x46 | n582 ;
  assign n867 = ( n582 & n604 ) | ( n582 & n866 ) | ( n604 & n866 ) ;
  assign n868 = n865 & ~n867 ;
  assign n869 = n857 & n868 ;
  assign n870 = ( n421 & n857 ) | ( n421 & n868 ) | ( n857 & n868 ) ;
  assign n871 = ( n858 & ~n869 ) | ( n858 & n870 ) | ( ~n869 & n870 ) ;
  assign n872 = x7 | n452 ;
  assign n873 = ( x1 & n529 ) | ( x1 & ~n872 ) | ( n529 & ~n872 ) ;
  assign n874 = ( n447 & n871 ) | ( n447 & ~n873 ) | ( n871 & ~n873 ) ;
  assign n875 = n846 & ~n874 ;
  assign n876 = ( n846 & n871 ) | ( n846 & ~n875 ) | ( n871 & ~n875 ) ;
  assign n877 = n310 & ~n403 ;
  assign n878 = ( n310 & n317 ) | ( n310 & n877 ) | ( n317 & n877 ) ;
  assign n879 = ( ~n310 & n317 ) | ( ~n310 & n877 ) | ( n317 & n877 ) ;
  assign n880 = ( n310 & ~n878 ) | ( n310 & n879 ) | ( ~n878 & n879 ) ;
  assign n881 = x46 & n603 ;
  assign n882 = ( n600 & n880 ) | ( n600 & n881 ) | ( n880 & n881 ) ;
  assign n883 = ( n600 & n881 ) | ( n600 & ~n882 ) | ( n881 & ~n882 ) ;
  assign n884 = ( n880 & ~n882 ) | ( n880 & n883 ) | ( ~n882 & n883 ) ;
  assign n885 = ( ~n857 & n865 ) | ( ~n857 & n884 ) | ( n865 & n884 ) ;
  assign n886 = n867 & n884 ;
  assign n887 = ( n857 & n885 ) | ( n857 & n886 ) | ( n885 & n886 ) ;
  assign n888 = ~n421 & n887 ;
  assign n889 = x6 | n452 ;
  assign n890 = ( x1 & n529 ) | ( x1 & ~n889 ) | ( n529 & ~n889 ) ;
  assign n891 = x14 & n487 ;
  assign n892 = x21 | n891 ;
  assign n893 = ( n491 & n891 ) | ( n491 & n892 ) | ( n891 & n892 ) ;
  assign n894 = x20 | n893 ;
  assign n895 = ( ~n484 & n893 ) | ( ~n484 & n894 ) | ( n893 & n894 ) ;
  assign n896 = x19 | n895 ;
  assign n897 = ( n480 & n895 ) | ( n480 & n896 ) | ( n895 & n896 ) ;
  assign n898 = x18 | n897 ;
  assign n899 = ( n476 & n897 ) | ( n476 & n898 ) | ( n897 & n898 ) ;
  assign n900 = x17 | n899 ;
  assign n901 = ( n473 & n899 ) | ( n473 & n900 ) | ( n899 & n900 ) ;
  assign n902 = x16 | n901 ;
  assign n903 = ( n471 & n901 ) | ( n471 & n902 ) | ( n901 & n902 ) ;
  assign n904 = x15 | n903 ;
  assign n905 = ( n467 & n903 ) | ( n467 & n904 ) | ( n903 & n904 ) ;
  assign n906 = ( ~x3 & x4 ) | ( ~x3 & n905 ) | ( x4 & n905 ) ;
  assign n907 = x38 & n487 ;
  assign n908 = n491 | n907 ;
  assign n909 = ( x7 & n907 ) | ( x7 & n908 ) | ( n907 & n908 ) ;
  assign n910 = n662 | n909 ;
  assign n911 = n722 | n910 ;
  assign n912 = x10 | n911 ;
  assign n913 = ( n476 & n911 ) | ( n476 & n912 ) | ( n911 & n912 ) ;
  assign n914 = x11 | n913 ;
  assign n915 = ( n473 & n913 ) | ( n473 & n914 ) | ( n913 & n914 ) ;
  assign n916 = x12 | n915 ;
  assign n917 = ( n471 & n915 ) | ( n471 & n916 ) | ( n915 & n916 ) ;
  assign n918 = x13 | n917 ;
  assign n919 = ( n467 & n917 ) | ( n467 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( x3 & x4 ) | ( x3 & n919 ) | ( x4 & n919 ) ;
  assign n921 = n906 | n920 ;
  assign n922 = x6 & n921 ;
  assign n923 = ( ~x4 & n921 ) | ( ~x4 & n922 ) | ( n921 & n922 ) ;
  assign n924 = x1 | n880 ;
  assign n925 = x3 | n924 ;
  assign n926 = ~n452 & n925 ;
  assign n927 = ( n923 & n925 ) | ( n923 & n926 ) | ( n925 & n926 ) ;
  assign n928 = ~n890 & n927 ;
  assign n929 = n447 & n928 ;
  assign n930 = ~n446 & n884 ;
  assign n931 = n929 | n930 ;
  assign n932 = ( n887 & ~n888 ) | ( n887 & n931 ) | ( ~n888 & n931 ) ;
  assign n933 = x40 & n487 ;
  assign n934 = n491 | n933 ;
  assign n935 = ( x9 & n933 ) | ( x9 & n934 ) | ( n933 & n934 ) ;
  assign n936 = x10 | n935 ;
  assign n937 = ( ~n484 & n935 ) | ( ~n484 & n936 ) | ( n935 & n936 ) ;
  assign n938 = x11 | n937 ;
  assign n939 = ( n480 & n937 ) | ( n480 & n938 ) | ( n937 & n938 ) ;
  assign n940 = x12 | n939 ;
  assign n941 = ( n476 & n939 ) | ( n476 & n940 ) | ( n939 & n940 ) ;
  assign n942 = x13 | n941 ;
  assign n943 = ( n473 & n941 ) | ( n473 & n942 ) | ( n941 & n942 ) ;
  assign n944 = x38 | n943 ;
  assign n945 = ( n471 & n943 ) | ( n471 & n944 ) | ( n943 & n944 ) ;
  assign n946 = x39 | n945 ;
  assign n947 = ( n467 & n945 ) | ( n467 & n946 ) | ( n945 & n946 ) ;
  assign n948 = ( x3 & ~n452 ) | ( x3 & n947 ) | ( ~n452 & n947 ) ;
  assign n949 = x16 & n487 ;
  assign n950 = n491 | n949 ;
  assign n951 = ( x7 & n949 ) | ( x7 & n950 ) | ( n949 & n950 ) ;
  assign n952 = x6 | n951 ;
  assign n953 = ( ~n484 & n951 ) | ( ~n484 & n952 ) | ( n951 & n952 ) ;
  assign n954 = x21 | n953 ;
  assign n955 = ( n480 & n953 ) | ( n480 & n954 ) | ( n953 & n954 ) ;
  assign n956 = x20 | n955 ;
  assign n957 = ( n476 & n955 ) | ( n476 & n956 ) | ( n955 & n956 ) ;
  assign n958 = x19 | n957 ;
  assign n959 = ( n473 & n957 ) | ( n473 & n958 ) | ( n957 & n958 ) ;
  assign n960 = x18 | n959 ;
  assign n961 = ( n471 & n959 ) | ( n471 & n960 ) | ( n959 & n960 ) ;
  assign n962 = x17 | n961 ;
  assign n963 = ( n467 & n961 ) | ( n467 & n962 ) | ( n961 & n962 ) ;
  assign n964 = ( x3 & n452 ) | ( x3 & ~n963 ) | ( n452 & ~n963 ) ;
  assign n965 = ~n948 & n964 ;
  assign n966 = ( x1 & x3 ) | ( x1 & ~n965 ) | ( x3 & ~n965 ) ;
  assign n967 = ~n593 & n966 ;
  assign n968 = ( n593 & ~n965 ) | ( n593 & n967 ) | ( ~n965 & n967 ) ;
  assign n969 = ~n446 & n865 ;
  assign n970 = ( n421 & n865 ) | ( n421 & ~n867 ) | ( n865 & ~n867 ) ;
  assign n971 = ( ~n868 & n969 ) | ( ~n868 & n970 ) | ( n969 & n970 ) ;
  assign n972 = x8 | n452 ;
  assign n973 = ( x1 & n529 ) | ( x1 & ~n972 ) | ( n529 & ~n972 ) ;
  assign n974 = ( n447 & n971 ) | ( n447 & ~n973 ) | ( n971 & ~n973 ) ;
  assign n975 = n968 & ~n974 ;
  assign n976 = ( n968 & n971 ) | ( n968 & ~n975 ) | ( n971 & ~n975 ) ;
  assign n977 = n579 | n932 ;
  assign n978 = ( ~n876 & n976 ) | ( ~n876 & n977 ) | ( n976 & n977 ) ;
  assign n979 = n876 | n978 ;
  assign n980 = n528 | n760 ;
  assign n981 = ( ~n702 & n812 ) | ( ~n702 & n980 ) | ( n812 & n980 ) ;
  assign n982 = n702 | n981 ;
  assign n983 = n979 | n982 ;
  assign n984 = n876 | n932 ;
  assign n985 = x47 & ~n984 ;
  assign n986 = x26 & n983 ;
  assign n987 = ( n984 & n985 ) | ( n984 & n986 ) | ( n985 & n986 ) ;
  assign n988 = ~x47 & x49 ;
  assign n989 = x26 & n988 ;
  assign n990 = ( n702 & n760 ) | ( n702 & n812 ) | ( n760 & n812 ) ;
  assign n991 = ( n702 & n760 ) | ( n702 & ~n990 ) | ( n760 & ~n990 ) ;
  assign n992 = ( n812 & ~n990 ) | ( n812 & n991 ) | ( ~n990 & n991 ) ;
  assign n993 = ~n528 & n992 ;
  assign n994 = n528 & ~n992 ;
  assign n995 = n993 | n994 ;
  assign n996 = n876 & ~n932 ;
  assign n997 = x26 & ~x47 ;
  assign n998 = ( ~n876 & n932 ) | ( ~n876 & n997 ) | ( n932 & n997 ) ;
  assign n999 = ( n996 & ~n997 ) | ( n996 & n998 ) | ( ~n997 & n998 ) ;
  assign n1000 = ~n579 & n976 ;
  assign n1001 = n579 | n976 ;
  assign n1002 = ( ~n976 & n1000 ) | ( ~n976 & n1001 ) | ( n1000 & n1001 ) ;
  assign n1003 = ( n995 & n999 ) | ( n995 & n1002 ) | ( n999 & n1002 ) ;
  assign n1004 = ( n999 & n1002 ) | ( n999 & ~n1003 ) | ( n1002 & ~n1003 ) ;
  assign n1005 = ( n995 & ~n1003 ) | ( n995 & n1004 ) | ( ~n1003 & n1004 ) ;
  assign n1006 = n989 | n1005 ;
  assign n1007 = n989 & n1005 ;
  assign n1008 = n1006 & ~n1007 ;
  assign n1009 = ( n876 & n932 ) | ( n876 & ~n1002 ) | ( n932 & ~n1002 ) ;
  assign n1010 = ( n876 & n932 ) | ( n876 & ~n1009 ) | ( n932 & ~n1009 ) ;
  assign n1011 = ( n1002 & n1009 ) | ( n1002 & ~n1010 ) | ( n1009 & ~n1010 ) ;
  assign n1012 = n995 & ~n1011 ;
  assign n1013 = ~n995 & n1011 ;
  assign n1014 = n1012 | n1013 ;
  assign y0 = ~n53 ;
  assign y1 = ~n55 ;
  assign y2 = ~n84 ;
  assign y3 = ~n99 ;
  assign y4 = ~n114 ;
  assign y5 = n382 ;
  assign y6 = n400 ;
  assign y7 = n418 ;
  assign y8 = n443 ;
  assign y9 = n528 ;
  assign y10 = n579 ;
  assign y11 = n623 ;
  assign y12 = n702 ;
  assign y13 = n760 ;
  assign y14 = n812 ;
  assign y15 = n876 ;
  assign y16 = n932 ;
  assign y17 = n976 ;
  assign y18 = n983 ;
  assign y19 = ~n987 ;
  assign y20 = ~n1008 ;
  assign y21 = ~n1014 ;
endmodule
