module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , y0 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 ;
  output y0 ;
  wire n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
  assign n10 = x6 & ~x7 ;
  assign n11 = x6 | x7 ;
  assign n12 = ( ~x6 & n10 ) | ( ~x6 & n11 ) | ( n10 & n11 ) ;
  assign n13 = ~x8 & n12 ;
  assign n14 = x1 & ~n13 ;
  assign n15 = ~x6 & x7 ;
  assign n16 = x7 | x8 ;
  assign n17 = ( ~x7 & n15 ) | ( ~x7 & n16 ) | ( n15 & n16 ) ;
  assign n18 = x0 & n17 ;
  assign n19 = x1 | n18 ;
  assign n20 = ~n14 & n19 ;
  assign n21 = ( x1 & ~x5 ) | ( x1 & n10 ) | ( ~x5 & n10 ) ;
  assign n22 = ( x5 & ~x6 ) | ( x5 & n10 ) | ( ~x6 & n10 ) ;
  assign n23 = n21 | n22 ;
  assign n24 = ( ~x0 & n20 ) | ( ~x0 & n23 ) | ( n20 & n23 ) ;
  assign n25 = x4 & ~n24 ;
  assign n26 = ( x4 & n20 ) | ( x4 & ~n25 ) | ( n20 & ~n25 ) ;
  assign n27 = ( ~x2 & x3 ) | ( ~x2 & n26 ) | ( x3 & n26 ) ;
  assign n28 = ( x1 & x2 ) | ( x1 & ~x8 ) | ( x2 & ~x8 ) ;
  assign n29 = ( x2 & x4 ) | ( x2 & x8 ) | ( x4 & x8 ) ;
  assign n30 = n28 & ~n29 ;
  assign n31 = ( x5 & x6 ) | ( x5 & ~n30 ) | ( x6 & ~n30 ) ;
  assign n32 = x4 & ~x7 ;
  assign n33 = x1 & x2 ;
  assign n34 = x1 & ~n33 ;
  assign n35 = n32 & n34 ;
  assign n36 = x0 & ~x4 ;
  assign n37 = x0 | x7 ;
  assign n38 = ( ~x0 & n36 ) | ( ~x0 & n37 ) | ( n36 & n37 ) ;
  assign n39 = ( ~n33 & n34 ) | ( ~n33 & n38 ) | ( n34 & n38 ) ;
  assign n40 = ( x2 & n35 ) | ( x2 & n39 ) | ( n35 & n39 ) ;
  assign n41 = x6 & n40 ;
  assign n42 = ( n30 & n31 ) | ( n30 & n41 ) | ( n31 & n41 ) ;
  assign n43 = x1 & x6 ;
  assign n44 = x6 & ~n43 ;
  assign n45 = ~x2 & n44 ;
  assign n46 = ( x4 & n43 ) | ( x4 & ~n44 ) | ( n43 & ~n44 ) ;
  assign n47 = ( x1 & n45 ) | ( x1 & ~n46 ) | ( n45 & ~n46 ) ;
  assign n48 = ( x0 & n42 ) | ( x0 & n47 ) | ( n42 & n47 ) ;
  assign n49 = x7 & ~n48 ;
  assign n50 = ( x7 & n42 ) | ( x7 & ~n49 ) | ( n42 & ~n49 ) ;
  assign n51 = ~x3 & n50 ;
  assign n52 = ( n26 & ~n27 ) | ( n26 & n51 ) | ( ~n27 & n51 ) ;
  assign n53 = ( x0 & x3 ) | ( x0 & x6 ) | ( x3 & x6 ) ;
  assign n54 = x0 & ~n53 ;
  assign n55 = ( x3 & ~n53 ) | ( x3 & n54 ) | ( ~n53 & n54 ) ;
  assign n56 = ( x2 & x5 ) | ( x2 & n55 ) | ( x5 & n55 ) ;
  assign n57 = x2 & ~x4 ;
  assign n58 = ( x3 & ~x7 ) | ( x3 & n57 ) | ( ~x7 & n57 ) ;
  assign n59 = ~x3 & n58 ;
  assign n60 = ( ~x0 & n12 ) | ( ~x0 & n59 ) | ( n12 & n59 ) ;
  assign n61 = x1 | n60 ;
  assign n62 = ( ~x1 & n59 ) | ( ~x1 & n61 ) | ( n59 & n61 ) ;
  assign n63 = x5 & n62 ;
  assign n64 = ( ~x2 & n56 ) | ( ~x2 & n63 ) | ( n56 & n63 ) ;
  assign n65 = ( x1 & x2 ) | ( x1 & x3 ) | ( x2 & x3 ) ;
  assign n66 = ~x3 & n65 ;
  assign n67 = ( ~x2 & n65 ) | ( ~x2 & n66 ) | ( n65 & n66 ) ;
  assign n68 = ( ~x0 & x4 ) | ( ~x0 & n67 ) | ( x4 & n67 ) ;
  assign n69 = x5 & ~n68 ;
  assign n70 = ( x5 & n67 ) | ( x5 & ~n69 ) | ( n67 & ~n69 ) ;
  assign n71 = ( ~x2 & x4 ) | ( ~x2 & x5 ) | ( x4 & x5 ) ;
  assign n72 = ( x2 & x3 ) | ( x2 & x4 ) | ( x3 & x4 ) ;
  assign n73 = ~n71 & n72 ;
  assign n74 = ~n70 & n73 ;
  assign n75 = ( ~n11 & n70 ) | ( ~n11 & n74 ) | ( n70 & n74 ) ;
  assign n76 = ( x3 & x4 ) | ( x3 & n12 ) | ( x4 & n12 ) ;
  assign n77 = ( x3 & x4 ) | ( x3 & x5 ) | ( x4 & x5 ) ;
  assign n78 = n76 & ~n77 ;
  assign n79 = ( x8 & n75 ) | ( x8 & n78 ) | ( n75 & n78 ) ;
  assign n80 = ~n64 & n79 ;
  assign n81 = ( x8 & n64 ) | ( x8 & n80 ) | ( n64 & n80 ) ;
  assign n82 = ( x4 & ~x5 ) | ( x4 & x8 ) | ( ~x5 & x8 ) ;
  assign n83 = ( x4 & x5 ) | ( x4 & x6 ) | ( x5 & x6 ) ;
  assign n84 = n82 & ~n83 ;
  assign n85 = ~x2 & n84 ;
  assign n86 = ~x2 & x8 ;
  assign n87 = ( x1 & x6 ) | ( x1 & n86 ) | ( x6 & n86 ) ;
  assign n88 = ~x1 & n87 ;
  assign n89 = ( x3 & ~x6 ) | ( x3 & n57 ) | ( ~x6 & n57 ) ;
  assign n90 = ( ~x1 & x6 ) | ( ~x1 & n57 ) | ( x6 & n57 ) ;
  assign n91 = n89 | n90 ;
  assign n92 = ( ~x5 & x8 ) | ( ~x5 & n91 ) | ( x8 & n91 ) ;
  assign n93 = x2 & x3 ;
  assign n94 = x3 & ~n93 ;
  assign n95 = x4 & n94 ;
  assign n96 = ( x6 & ~n93 ) | ( x6 & n94 ) | ( ~n93 & n94 ) ;
  assign n97 = ( x2 & n95 ) | ( x2 & n96 ) | ( n95 & n96 ) ;
  assign n98 = ~x8 & n97 ;
  assign n99 = ( n91 & ~n92 ) | ( n91 & n98 ) | ( ~n92 & n98 ) ;
  assign n100 = n88 | n99 ;
  assign n101 = ( n84 & ~n85 ) | ( n84 & n100 ) | ( ~n85 & n100 ) ;
  assign n102 = ( x0 & ~x7 ) | ( x0 & n101 ) | ( ~x7 & n101 ) ;
  assign n103 = ( x2 & x4 ) | ( x2 & ~x7 ) | ( x4 & ~x7 ) ;
  assign n104 = ( x2 & x7 ) | ( x2 & x8 ) | ( x7 & x8 ) ;
  assign n105 = n103 & ~n104 ;
  assign n106 = x5 & n105 ;
  assign n107 = x3 & n106 ;
  assign n108 = ~x7 & x8 ;
  assign n109 = x6 & ~n108 ;
  assign n110 = x1 & x3 ;
  assign n111 = x6 | n110 ;
  assign n112 = ~n109 & n111 ;
  assign n113 = ( ~x4 & n107 ) | ( ~x4 & n112 ) | ( n107 & n112 ) ;
  assign n114 = x2 & ~n113 ;
  assign n115 = ( x2 & n107 ) | ( x2 & ~n114 ) | ( n107 & ~n114 ) ;
  assign n116 = ~x0 & n115 ;
  assign n117 = ( n101 & ~n102 ) | ( n101 & n116 ) | ( ~n102 & n116 ) ;
  assign n118 = x5 & n17 ;
  assign n119 = ~x4 & n118 ;
  assign n120 = ( ~x3 & n38 ) | ( ~x3 & n119 ) | ( n38 & n119 ) ;
  assign n121 = x8 & ~n120 ;
  assign n122 = ( x8 & n119 ) | ( x8 & ~n121 ) | ( n119 & ~n121 ) ;
  assign n123 = x4 & x6 ;
  assign n124 = x3 & ~x5 ;
  assign n125 = ( x4 & x6 ) | ( x4 & ~n124 ) | ( x6 & ~n124 ) ;
  assign n126 = ( ~n123 & n124 ) | ( ~n123 & n125 ) | ( n124 & n125 ) ;
  assign n127 = ( ~x8 & n122 ) | ( ~x8 & n126 ) | ( n122 & n126 ) ;
  assign n128 = x7 & ~n127 ;
  assign n129 = ( x7 & n122 ) | ( x7 & ~n128 ) | ( n122 & ~n128 ) ;
  assign n130 = x2 & n129 ;
  assign n131 = ( x2 & x3 ) | ( x2 & x5 ) | ( x3 & x5 ) ;
  assign n132 = ~x3 & n131 ;
  assign n133 = ( ~x2 & n131 ) | ( ~x2 & n132 ) | ( n131 & n132 ) ;
  assign n134 = ~x0 & n133 ;
  assign n135 = ~x4 & n134 ;
  assign n136 = ( x6 & x7 ) | ( x6 & ~x8 ) | ( x7 & ~x8 ) ;
  assign n137 = ( x4 & x6 ) | ( x4 & x8 ) | ( x6 & x8 ) ;
  assign n138 = ~n136 & n137 ;
  assign n139 = ( x2 & ~x5 ) | ( x2 & n138 ) | ( ~x5 & n138 ) ;
  assign n140 = x2 & ~x7 ;
  assign n141 = x2 | x6 ;
  assign n142 = ( ~x2 & n140 ) | ( ~x2 & n141 ) | ( n140 & n141 ) ;
  assign n143 = x0 & x3 ;
  assign n144 = x3 & ~n143 ;
  assign n145 = n142 & n144 ;
  assign n146 = ~x4 & x6 ;
  assign n147 = ( ~n143 & n144 ) | ( ~n143 & n146 ) | ( n144 & n146 ) ;
  assign n148 = ( x0 & n145 ) | ( x0 & n147 ) | ( n145 & n147 ) ;
  assign n149 = ~x5 & n148 ;
  assign n150 = ( ~x2 & n139 ) | ( ~x2 & n149 ) | ( n139 & n149 ) ;
  assign n151 = n135 | n150 ;
  assign n152 = ( n129 & ~n130 ) | ( n129 & n151 ) | ( ~n130 & n151 ) ;
  assign n153 = ~x1 & n152 ;
  assign n154 = ( x0 & x3 ) | ( x0 & ~x6 ) | ( x3 & ~x6 ) ;
  assign n155 = ( x3 & x6 ) | ( x3 & x7 ) | ( x6 & x7 ) ;
  assign n156 = ~n154 & n155 ;
  assign n157 = ( x4 & x5 ) | ( x4 & n156 ) | ( x5 & n156 ) ;
  assign n158 = ( x3 & x5 ) | ( x3 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n159 = ( x2 & x5 ) | ( x2 & x7 ) | ( x5 & x7 ) ;
  assign n160 = n158 & ~n159 ;
  assign n161 = x1 & ~n160 ;
  assign n162 = x5 & n12 ;
  assign n163 = x1 | n162 ;
  assign n164 = ~n161 & n163 ;
  assign n165 = x4 & n164 ;
  assign n166 = ( ~x5 & n157 ) | ( ~x5 & n165 ) | ( n157 & n165 ) ;
  assign n167 = x0 & ~x7 ;
  assign n168 = x1 & n167 ;
  assign n169 = ( x3 & ~x5 ) | ( x3 & n168 ) | ( ~x5 & n168 ) ;
  assign n170 = x7 & ~n169 ;
  assign n171 = ( x7 & n168 ) | ( x7 & ~n170 ) | ( n168 & ~n170 ) ;
  assign n172 = ( ~x6 & n166 ) | ( ~x6 & n171 ) | ( n166 & n171 ) ;
  assign n173 = x2 & ~n172 ;
  assign n174 = ( x2 & n166 ) | ( x2 & ~n173 ) | ( n166 & ~n173 ) ;
  assign n175 = ( ~x1 & x4 ) | ( ~x1 & x7 ) | ( x4 & x7 ) ;
  assign n176 = ( x1 & x3 ) | ( x1 & x4 ) | ( x3 & x4 ) ;
  assign n177 = n175 & ~n176 ;
  assign n178 = ~n47 & n177 ;
  assign n179 = x0 & x5 ;
  assign n180 = ( n47 & n178 ) | ( n47 & n179 ) | ( n178 & n179 ) ;
  assign n181 = ~x1 & x7 ;
  assign n182 = ( x2 & ~x5 ) | ( x2 & n181 ) | ( ~x5 & n181 ) ;
  assign n183 = ( x5 & ~x7 ) | ( x5 & n181 ) | ( ~x7 & n181 ) ;
  assign n184 = n182 | n183 ;
  assign n185 = ( x3 & n146 ) | ( x3 & ~n184 ) | ( n146 & ~n184 ) ;
  assign n186 = n184 & n185 ;
  assign n187 = ( ~x8 & n180 ) | ( ~x8 & n186 ) | ( n180 & n186 ) ;
  assign n188 = ~n174 & n187 ;
  assign n189 = ( ~x8 & n174 ) | ( ~x8 & n188 ) | ( n174 & n188 ) ;
  assign n190 = x3 & x4 ;
  assign n191 = ( x1 & x2 ) | ( x1 & n190 ) | ( x2 & n190 ) ;
  assign n192 = x3 | x4 ;
  assign n193 = ( x1 & x2 ) | ( x1 & n192 ) | ( x2 & n192 ) ;
  assign n194 = ~n191 & n193 ;
  assign n195 = ~x3 & x4 ;
  assign n196 = ( x3 & ~x4 ) | ( x3 & n12 ) | ( ~x4 & n12 ) ;
  assign n197 = ( x8 & n195 ) | ( x8 & n196 ) | ( n195 & n196 ) ;
  assign n198 = x2 & n197 ;
  assign n199 = x5 & ~x7 ;
  assign n200 = ( x3 & x6 ) | ( x3 & n199 ) | ( x6 & n199 ) ;
  assign n201 = ~x6 & n200 ;
  assign n202 = ( x4 & x5 ) | ( x4 & ~n12 ) | ( x5 & ~n12 ) ;
  assign n203 = n76 & ~n202 ;
  assign n204 = n201 | n203 ;
  assign n205 = ( n197 & ~n198 ) | ( n197 & n204 ) | ( ~n198 & n204 ) ;
  assign n206 = ( ~x0 & x1 ) | ( ~x0 & n205 ) | ( x1 & n205 ) ;
  assign n207 = ( x0 & x3 ) | ( x0 & n57 ) | ( x3 & n57 ) ;
  assign n208 = ( x0 & x3 ) | ( x0 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n209 = n207 & ~n208 ;
  assign n210 = ( x0 & x2 ) | ( x0 & ~x5 ) | ( x2 & ~x5 ) ;
  assign n211 = ~x0 & x8 ;
  assign n212 = ( x2 & x5 ) | ( x2 & x8 ) | ( x5 & x8 ) ;
  assign n213 = ( n210 & n211 ) | ( n210 & ~n212 ) | ( n211 & ~n212 ) ;
  assign n214 = ( x3 & n209 ) | ( x3 & n213 ) | ( n209 & n213 ) ;
  assign n215 = x4 & ~n214 ;
  assign n216 = ( x4 & n209 ) | ( x4 & ~n215 ) | ( n209 & ~n215 ) ;
  assign n217 = ~x1 & n216 ;
  assign n218 = ( n205 & ~n206 ) | ( n205 & n217 ) | ( ~n206 & n217 ) ;
  assign n219 = ( x0 & ~x5 ) | ( x0 & n218 ) | ( ~x5 & n218 ) ;
  assign n220 = n194 & ~n219 ;
  assign n221 = ( n194 & n218 ) | ( n194 & ~n220 ) | ( n218 & ~n220 ) ;
  assign n222 = n189 | n221 ;
  assign n223 = ( n152 & ~n153 ) | ( n152 & n222 ) | ( ~n153 & n222 ) ;
  assign n224 = n117 | n223 ;
  assign n225 = ( ~n52 & n81 ) | ( ~n52 & n224 ) | ( n81 & n224 ) ;
  assign n226 = n52 | n225 ;
  assign y0 = n226 ;
endmodule
