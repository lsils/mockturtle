module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 ;
  wire n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 ;
  assign n46 = ~x18 & x19 ;
  assign n47 = x21 & n46 ;
  assign n48 = x26 & n47 ;
  assign n49 = ~x29 & x30 ;
  assign n50 = ( x28 & n48 ) | ( x28 & n49 ) | ( n48 & n49 ) ;
  assign n51 = ~x28 & n50 ;
  assign n52 = ~x0 & x18 ;
  assign n59 = ~x20 & x21 ;
  assign n60 = ( x19 & n52 ) | ( x19 & n59 ) | ( n52 & n59 ) ;
  assign n61 = ~x19 & n60 ;
  assign n62 = ( x28 & n49 ) | ( x28 & n61 ) | ( n49 & n61 ) ;
  assign n63 = ~x28 & n62 ;
  assign n53 = x19 & x21 ;
  assign n54 = ( x20 & ~n52 ) | ( x20 & n53 ) | ( ~n52 & n53 ) ;
  assign n55 = n52 & n54 ;
  assign n56 = x24 & x30 ;
  assign n57 = ( x29 & n55 ) | ( x29 & n56 ) | ( n55 & n56 ) ;
  assign n58 = ~x29 & n57 ;
  assign n67 = x10 & x21 ;
  assign n68 = ( x18 & x19 ) | ( x18 & n67 ) | ( x19 & n67 ) ;
  assign n69 = ~x18 & n68 ;
  assign n70 = x25 & ~x29 ;
  assign n71 = ( x28 & n69 ) | ( x28 & n70 ) | ( n69 & n70 ) ;
  assign n72 = ~x28 & n71 ;
  assign n73 = x30 & n72 ;
  assign n64 = x24 & n47 ;
  assign n65 = ( x28 & n49 ) | ( x28 & n64 ) | ( n49 & n64 ) ;
  assign n66 = ~x28 & n65 ;
  assign n74 = ~x18 & x20 ;
  assign n75 = ( x0 & ~x19 ) | ( x0 & n74 ) | ( ~x19 & n74 ) ;
  assign n76 = ~x0 & n75 ;
  assign n77 = x21 & n76 ;
  assign n78 = ( x24 & x29 ) | ( x24 & n77 ) | ( x29 & n77 ) ;
  assign n79 = ~x29 & n78 ;
  assign n80 = x30 & n79 ;
  assign n81 = n66 | n80 ;
  assign n82 = n73 | n81 ;
  assign n83 = n58 | n82 ;
  assign n84 = ( ~n51 & n63 ) | ( ~n51 & n83 ) | ( n63 & n83 ) ;
  assign n85 = n51 | n84 ;
  assign n86 = n58 | n80 ;
  assign n87 = n51 | n73 ;
  assign n88 = n51 | n58 ;
  assign n89 = n66 | n88 ;
  assign n90 = ~x19 & x20 ;
  assign n91 = ( x0 & x18 ) | ( x0 & n90 ) | ( x18 & n90 ) ;
  assign n92 = ~x18 & n91 ;
  assign n93 = x21 & n92 ;
  assign n94 = ( x29 & n56 ) | ( x29 & n93 ) | ( n56 & n93 ) ;
  assign n95 = ~x29 & n94 ;
  assign n102 = x0 & x19 ;
  assign n103 = x18 & n102 ;
  assign n104 = x20 & n103 ;
  assign n105 = x21 & x30 ;
  assign n106 = ( x29 & n104 ) | ( x29 & n105 ) | ( n104 & n105 ) ;
  assign n107 = ~x29 & n106 ;
  assign n96 = x0 & ~x19 ;
  assign n97 = x18 & n96 ;
  assign n98 = ~x28 & n97 ;
  assign n99 = ( x20 & x21 ) | ( x20 & n98 ) | ( x21 & n98 ) ;
  assign n100 = ~x20 & n99 ;
  assign n101 = n49 & n100 ;
  assign n108 = x0 & x21 ;
  assign n109 = ( x18 & x19 ) | ( x18 & n108 ) | ( x19 & n108 ) ;
  assign n110 = ~x18 & n109 ;
  assign n111 = x28 & x30 ;
  assign n112 = ( x29 & n110 ) | ( x29 & n111 ) | ( n110 & n111 ) ;
  assign n113 = ~x29 & n112 ;
  assign n114 = n101 | n113 ;
  assign n115 = ( ~n95 & n107 ) | ( ~n95 & n114 ) | ( n107 & n114 ) ;
  assign n116 = n95 | n115 ;
  assign n243 = x10 & x18 ;
  assign n244 = ( x0 & x11 ) | ( x0 & n243 ) | ( x11 & n243 ) ;
  assign n245 = ~x11 & n244 ;
  assign n246 = x19 & ~x21 ;
  assign n247 = ( x20 & n245 ) | ( x20 & n246 ) | ( n245 & n246 ) ;
  assign n248 = ~x20 & n247 ;
  assign n249 = x25 & n248 ;
  assign n250 = ( x29 & x30 ) | ( x29 & n249 ) | ( x30 & n249 ) ;
  assign n251 = ~x30 & n250 ;
  assign n266 = x3 & x19 ;
  assign n267 = ( ~x0 & x18 ) | ( ~x0 & n266 ) | ( x18 & n266 ) ;
  assign n268 = x0 & n267 ;
  assign n269 = x20 & x27 ;
  assign n270 = ( x21 & n268 ) | ( x21 & n269 ) | ( n268 & n269 ) ;
  assign n271 = ~x21 & n270 ;
  assign n272 = ~x29 & n271 ;
  assign n273 = ~x30 & n272 ;
  assign n138 = x0 & ~x5 ;
  assign n258 = x19 & n138 ;
  assign n259 = x18 & n258 ;
  assign n260 = x20 & ~x27 ;
  assign n261 = ( x21 & n259 ) | ( x21 & n260 ) | ( n259 & n260 ) ;
  assign n262 = ~x21 & n261 ;
  assign n263 = x30 & n262 ;
  assign n264 = ( x28 & x29 ) | ( x28 & n263 ) | ( x29 & n263 ) ;
  assign n265 = ~x28 & n264 ;
  assign n274 = ~x4 & x19 ;
  assign n275 = ( x0 & x18 ) | ( x0 & n274 ) | ( x18 & n274 ) ;
  assign n276 = ~x0 & n275 ;
  assign n277 = ( x21 & n260 ) | ( x21 & n276 ) | ( n260 & n276 ) ;
  assign n278 = ~x21 & n277 ;
  assign n279 = x28 & n278 ;
  assign n280 = ( x29 & x30 ) | ( x29 & n279 ) | ( x30 & n279 ) ;
  assign n281 = ~x30 & n280 ;
  assign n282 = n265 | n281 ;
  assign n283 = n273 | n282 ;
  assign n252 = ~x21 & x26 ;
  assign n253 = ( x20 & n103 ) | ( x20 & n252 ) | ( n103 & n252 ) ;
  assign n254 = ~x20 & n253 ;
  assign n255 = ~x30 & n254 ;
  assign n256 = ( x28 & x29 ) | ( x28 & n255 ) | ( x29 & n255 ) ;
  assign n257 = ~x28 & n256 ;
  assign n284 = x11 & x19 ;
  assign n285 = ( ~x0 & x18 ) | ( ~x0 & n284 ) | ( x18 & n284 ) ;
  assign n286 = x0 & n285 ;
  assign n287 = ( x20 & n252 ) | ( x20 & n286 ) | ( n252 & n286 ) ;
  assign n288 = ~x20 & n287 ;
  assign n289 = ( x29 & n111 ) | ( x29 & n288 ) | ( n111 & n288 ) ;
  assign n290 = ~x29 & n289 ;
  assign n291 = ( x11 & x18 ) | ( x11 & n102 ) | ( x18 & n102 ) ;
  assign n292 = ~x11 & n291 ;
  assign n293 = ( x20 & n252 ) | ( x20 & n292 ) | ( n252 & n292 ) ;
  assign n294 = ~x20 & n293 ;
  assign n295 = ( x29 & n111 ) | ( x29 & n294 ) | ( n111 & n294 ) ;
  assign n296 = ~x29 & n295 ;
  assign n297 = n290 | n296 ;
  assign n298 = n257 | n297 ;
  assign n299 = ( ~n251 & n283 ) | ( ~n251 & n298 ) | ( n283 & n298 ) ;
  assign n300 = n251 | n299 ;
  assign n117 = x0 & ~x3 ;
  assign n118 = ( x2 & ~x18 ) | ( x2 & n117 ) | ( ~x18 & n117 ) ;
  assign n119 = ~x2 & n118 ;
  assign n120 = ~x21 & n119 ;
  assign n121 = ( x19 & x20 ) | ( x19 & n120 ) | ( x20 & n120 ) ;
  assign n122 = ~x19 & n121 ;
  assign n123 = ( x29 & n111 ) | ( x29 & n122 ) | ( n111 & n122 ) ;
  assign n124 = ~x29 & n123 ;
  assign n133 = ~x28 & n92 ;
  assign n134 = ( x21 & x23 ) | ( x21 & n133 ) | ( x23 & n133 ) ;
  assign n135 = ~x21 & n134 ;
  assign n136 = ~x30 & n135 ;
  assign n137 = x29 & n136 ;
  assign n125 = x2 & ~x18 ;
  assign n126 = ( x0 & x3 ) | ( x0 & n125 ) | ( x3 & n125 ) ;
  assign n127 = ~x3 & n126 ;
  assign n128 = ~x20 & n127 ;
  assign n129 = ( x19 & ~x21 ) | ( x19 & n128 ) | ( ~x21 & n128 ) ;
  assign n130 = ~x19 & n129 ;
  assign n131 = ( x29 & n111 ) | ( x29 & n130 ) | ( n111 & n130 ) ;
  assign n132 = ~x29 & n131 ;
  assign n139 = ~x15 & n138 ;
  assign n140 = x11 & n139 ;
  assign n141 = x18 & x20 ;
  assign n142 = ( x19 & n140 ) | ( x19 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ~x19 & n142 ;
  assign n144 = x21 & n143 ;
  assign n145 = ( x26 & x28 ) | ( x26 & n144 ) | ( x28 & n144 ) ;
  assign n146 = ~x28 & n145 ;
  assign n147 = n49 & n146 ;
  assign n158 = ~x11 & n138 ;
  assign n159 = ~x15 & n158 ;
  assign n160 = ( x19 & n141 ) | ( x19 & n159 ) | ( n141 & n159 ) ;
  assign n161 = ~x19 & n160 ;
  assign n162 = x21 & n161 ;
  assign n163 = ( x26 & x28 ) | ( x26 & n162 ) | ( x28 & n162 ) ;
  assign n164 = ~x28 & n163 ;
  assign n165 = n49 & n164 ;
  assign n148 = x11 & n138 ;
  assign n149 = x10 & n148 ;
  assign n150 = ~x19 & n149 ;
  assign n151 = ( x15 & x18 ) | ( x15 & n150 ) | ( x18 & n150 ) ;
  assign n152 = ~x15 & n151 ;
  assign n153 = x20 & x25 ;
  assign n154 = ( x21 & ~n152 ) | ( x21 & n153 ) | ( ~n152 & n153 ) ;
  assign n155 = n152 & n154 ;
  assign n156 = ( x28 & n49 ) | ( x28 & n155 ) | ( n49 & n155 ) ;
  assign n157 = ~x28 & n156 ;
  assign n166 = ( x3 & ~x18 ) | ( x3 & n138 ) | ( ~x18 & n138 ) ;
  assign n167 = ~x3 & n166 ;
  assign n168 = ~x20 & n167 ;
  assign n169 = ( x19 & ~x21 ) | ( x19 & n168 ) | ( ~x21 & n168 ) ;
  assign n170 = ~x19 & n169 ;
  assign n171 = ~x30 & n170 ;
  assign n172 = ( x28 & x29 ) | ( x28 & n171 ) | ( x29 & n171 ) ;
  assign n173 = ~x28 & n172 ;
  assign n174 = n157 | n173 ;
  assign n175 = ( ~n147 & n165 ) | ( ~n147 & n174 ) | ( n165 & n174 ) ;
  assign n176 = n147 | n175 ;
  assign n177 = n132 | n176 ;
  assign n178 = ( ~n124 & n137 ) | ( ~n124 & n177 ) | ( n137 & n177 ) ;
  assign n179 = n124 | n178 ;
  assign n212 = x22 & x30 ;
  assign n213 = ( x29 & n93 ) | ( x29 & n212 ) | ( n93 & n212 ) ;
  assign n214 = ~x29 & n213 ;
  assign n215 = x10 & ~x18 ;
  assign n216 = ( x0 & x11 ) | ( x0 & n215 ) | ( x11 & n215 ) ;
  assign n217 = ~x11 & n216 ;
  assign n218 = x21 & n217 ;
  assign n219 = ( x19 & x20 ) | ( x19 & n218 ) | ( x20 & n218 ) ;
  assign n220 = ~x19 & n219 ;
  assign n221 = x25 & x30 ;
  assign n222 = ( x29 & n220 ) | ( x29 & n221 ) | ( n220 & n221 ) ;
  assign n223 = ~x29 & n222 ;
  assign n224 = n214 | n223 ;
  assign n187 = x11 & ~x19 ;
  assign n188 = ( x0 & x18 ) | ( x0 & n187 ) | ( x18 & n187 ) ;
  assign n189 = ~x18 & n188 ;
  assign n190 = x20 & x26 ;
  assign n191 = ( x21 & ~n189 ) | ( x21 & n190 ) | ( ~n189 & n190 ) ;
  assign n192 = n189 & n191 ;
  assign n193 = n49 & n192 ;
  assign n180 = ( x15 & n46 ) | ( x15 & n138 ) | ( n46 & n138 ) ;
  assign n181 = ~x15 & n180 ;
  assign n182 = x20 & x22 ;
  assign n183 = ( x21 & ~n181 ) | ( x21 & n182 ) | ( ~n181 & n182 ) ;
  assign n184 = n181 & n183 ;
  assign n185 = ( x28 & n49 ) | ( x28 & n184 ) | ( n49 & n184 ) ;
  assign n186 = ~x28 & n185 ;
  assign n194 = x10 & n158 ;
  assign n195 = ~x19 & n194 ;
  assign n196 = ( x15 & x18 ) | ( x15 & n195 ) | ( x18 & n195 ) ;
  assign n197 = ~x15 & n196 ;
  assign n198 = ( x21 & n153 ) | ( x21 & ~n197 ) | ( n153 & ~n197 ) ;
  assign n199 = n197 & n198 ;
  assign n200 = ( x28 & n49 ) | ( x28 & n199 ) | ( n49 & n199 ) ;
  assign n201 = ~x28 & n200 ;
  assign n202 = ~x19 & n138 ;
  assign n203 = ( x15 & x18 ) | ( x15 & n202 ) | ( x18 & n202 ) ;
  assign n204 = ~x15 & n203 ;
  assign n205 = ( x21 & n182 ) | ( x21 & ~n204 ) | ( n182 & ~n204 ) ;
  assign n206 = n204 & n205 ;
  assign n207 = ( x28 & n49 ) | ( x28 & n206 ) | ( n49 & n206 ) ;
  assign n208 = ~x28 & n207 ;
  assign n209 = n201 | n208 ;
  assign n210 = n186 | n209 ;
  assign n211 = n193 | n210 ;
  assign n225 = x0 & x10 ;
  assign n226 = ( x11 & x18 ) | ( x11 & n225 ) | ( x18 & n225 ) ;
  assign n227 = ~x18 & n226 ;
  assign n228 = x21 & n227 ;
  assign n229 = ( x19 & x20 ) | ( x19 & n228 ) | ( x20 & n228 ) ;
  assign n230 = ~x19 & n229 ;
  assign n231 = ( x29 & n221 ) | ( x29 & n230 ) | ( n221 & n230 ) ;
  assign n232 = ~x29 & n231 ;
  assign n233 = x0 & ~x18 ;
  assign n234 = ( x11 & ~x19 ) | ( x11 & n233 ) | ( ~x19 & n233 ) ;
  assign n235 = ~x11 & n234 ;
  assign n236 = ( x21 & n190 ) | ( x21 & ~n235 ) | ( n190 & ~n235 ) ;
  assign n237 = n235 & n236 ;
  assign n238 = n49 & n237 ;
  assign n239 = n232 | n238 ;
  assign n240 = n211 | n239 ;
  assign n241 = ( ~n179 & n224 ) | ( ~n179 & n240 ) | ( n224 & n240 ) ;
  assign n242 = n179 | n241 ;
  assign n301 = ~x21 & x22 ;
  assign n302 = ( x20 & n103 ) | ( x20 & n301 ) | ( n103 & n301 ) ;
  assign n303 = ~x20 & n302 ;
  assign n304 = ~x30 & n303 ;
  assign n305 = x29 & n304 ;
  assign n319 = x0 & x20 ;
  assign n320 = ( x18 & x19 ) | ( x18 & n319 ) | ( x19 & n319 ) ;
  assign n321 = ~x18 & n320 ;
  assign n322 = n301 & n321 ;
  assign n323 = x28 & n322 ;
  assign n324 = ( x29 & x30 ) | ( x29 & n323 ) | ( x30 & n323 ) ;
  assign n325 = ~x30 & n324 ;
  assign n313 = n46 & n138 ;
  assign n314 = ( x21 & n182 ) | ( x21 & n313 ) | ( n182 & n313 ) ;
  assign n315 = ~x21 & n314 ;
  assign n316 = ~x30 & n315 ;
  assign n317 = ( x28 & x29 ) | ( x28 & n316 ) | ( x29 & n316 ) ;
  assign n318 = ~x28 & n317 ;
  assign n326 = x0 & x17 ;
  assign n327 = ( x18 & x19 ) | ( x18 & n326 ) | ( x19 & n326 ) ;
  assign n328 = ~x19 & n327 ;
  assign n329 = ( x21 & n190 ) | ( x21 & n328 ) | ( n190 & n328 ) ;
  assign n330 = ~x21 & n329 ;
  assign n331 = ~x30 & n330 ;
  assign n332 = ( x28 & x29 ) | ( x28 & n331 ) | ( x29 & n331 ) ;
  assign n333 = ~x28 & n332 ;
  assign n334 = ( x17 & x18 ) | ( x17 & n96 ) | ( x18 & n96 ) ;
  assign n335 = ~x17 & n334 ;
  assign n336 = ( x21 & n190 ) | ( x21 & n335 ) | ( n190 & n335 ) ;
  assign n337 = ~x21 & n336 ;
  assign n338 = ~x30 & n337 ;
  assign n339 = ( x28 & x29 ) | ( x28 & n338 ) | ( x29 & n338 ) ;
  assign n340 = ~x28 & n339 ;
  assign n341 = n333 | n340 ;
  assign n342 = n318 | n341 ;
  assign n343 = n325 | n342 ;
  assign n306 = ( ~x0 & x11 ) | ( ~x0 & n243 ) | ( x11 & n243 ) ;
  assign n307 = x0 & n306 ;
  assign n308 = ( x20 & n246 ) | ( x20 & n307 ) | ( n246 & n307 ) ;
  assign n309 = ~x20 & n308 ;
  assign n310 = x25 & n309 ;
  assign n311 = ( x29 & x30 ) | ( x29 & n310 ) | ( x30 & n310 ) ;
  assign n312 = ~x30 & n311 ;
  assign n344 = ( x11 & x18 ) | ( x11 & n96 ) | ( x18 & n96 ) ;
  assign n345 = ~x11 & n344 ;
  assign n346 = ( x21 & n190 ) | ( x21 & n345 ) | ( n190 & n345 ) ;
  assign n347 = ~x21 & n346 ;
  assign n348 = ( x29 & n111 ) | ( x29 & n347 ) | ( n111 & n347 ) ;
  assign n349 = ~x29 & n348 ;
  assign n350 = x0 & x11 ;
  assign n351 = ( x18 & x19 ) | ( x18 & n350 ) | ( x19 & n350 ) ;
  assign n352 = ~x19 & n351 ;
  assign n353 = ( x21 & n190 ) | ( x21 & n352 ) | ( n190 & n352 ) ;
  assign n354 = ~x21 & n353 ;
  assign n355 = ( x29 & n111 ) | ( x29 & n354 ) | ( n111 & n354 ) ;
  assign n356 = ~x29 & n355 ;
  assign n357 = n349 | n356 ;
  assign n358 = n312 | n357 ;
  assign n359 = ( ~n305 & n343 ) | ( ~n305 & n358 ) | ( n343 & n358 ) ;
  assign n360 = n305 | n359 ;
  assign n361 = n242 | n360 ;
  assign n362 = n300 | n361 ;
  assign n363 = n201 | n232 ;
  assign n364 = n223 | n363 ;
  assign n365 = n251 | n364 ;
  assign n366 = ( ~n157 & n312 ) | ( ~n157 & n365 ) | ( n312 & n365 ) ;
  assign n367 = n157 | n366 ;
  assign n368 = n186 | n224 ;
  assign n369 = n238 | n368 ;
  assign n370 = n173 | n209 ;
  assign n371 = ( ~n165 & n369 ) | ( ~n165 & n370 ) | ( n369 & n370 ) ;
  assign n372 = n165 | n371 ;
  assign n373 = n124 | n356 ;
  assign n374 = ( ~n305 & n325 ) | ( ~n305 & n373 ) | ( n325 & n373 ) ;
  assign n375 = n305 | n374 ;
  assign n376 = n296 | n375 ;
  assign n377 = ( n251 & ~n281 ) | ( n251 & n376 ) | ( ~n281 & n376 ) ;
  assign n378 = n281 | n377 ;
  assign n379 = n372 | n378 ;
  assign n380 = n137 | n273 ;
  assign n381 = n132 | n380 ;
  assign n397 = ~x19 & x21 ;
  assign n398 = ( x18 & ~x20 ) | ( x18 & n397 ) | ( ~x20 & n397 ) ;
  assign n399 = ~x18 & n398 ;
  assign n400 = x22 & x29 ;
  assign n401 = ( x28 & n399 ) | ( x28 & n400 ) | ( n399 & n400 ) ;
  assign n402 = ~x28 & n401 ;
  assign n403 = x30 & n402 ;
  assign n382 = x18 | x20 ;
  assign n383 = ( ~x9 & x19 ) | ( ~x9 & n382 ) | ( x19 & n382 ) ;
  assign n384 = x9 | n383 ;
  assign n385 = x21 & ~n384 ;
  assign n386 = ( x22 & x28 ) | ( x22 & n385 ) | ( x28 & n385 ) ;
  assign n387 = ~x28 & n386 ;
  assign n388 = ~x30 & n387 ;
  assign n389 = x29 & n388 ;
  assign n390 = ~x38 & n389 ;
  assign n391 = ~x39 & n390 ;
  assign n392 = ~x41 & n391 ;
  assign n393 = ( x40 & ~x42 ) | ( x40 & n392 ) | ( ~x42 & n392 ) ;
  assign n394 = ~x40 & n393 ;
  assign n395 = ~x43 & x44 ;
  assign n396 = n394 & n395 ;
  assign n406 = x39 & x42 ;
  assign n407 = ( x41 & n390 ) | ( x41 & n406 ) | ( n390 & n406 ) ;
  assign n408 = ~x41 & n407 ;
  assign n404 = ~x41 & x42 ;
  assign n405 = n391 & n404 ;
  assign n409 = x39 & ~x42 ;
  assign n410 = ( x41 & n390 ) | ( x41 & n409 ) | ( n390 & n409 ) ;
  assign n411 = ~x41 & n410 ;
  assign n412 = n405 | n411 ;
  assign n413 = n408 | n412 ;
  assign n414 = n396 | n413 ;
  assign n415 = n403 | n414 ;
  assign n444 = ( x17 & x19 ) | ( x17 & n141 ) | ( x19 & n141 ) ;
  assign n445 = ~x19 & n444 ;
  assign n446 = n252 & n445 ;
  assign n447 = ~x28 & n446 ;
  assign n448 = ~x30 & n447 ;
  assign n449 = x29 & n448 ;
  assign n457 = ( x17 & x18 ) | ( x17 & n90 ) | ( x18 & n90 ) ;
  assign n458 = ~x17 & n457 ;
  assign n459 = ~x28 & n458 ;
  assign n460 = ( x21 & x26 ) | ( x21 & n459 ) | ( x26 & n459 ) ;
  assign n461 = ~x21 & n460 ;
  assign n462 = x30 & n461 ;
  assign n463 = x29 & n462 ;
  assign n450 = x18 & ~x21 ;
  assign n451 = ( x19 & x20 ) | ( x19 & n450 ) | ( x20 & n450 ) ;
  assign n452 = ~x19 & n451 ;
  assign n453 = x26 & x29 ;
  assign n454 = ( x28 & ~n452 ) | ( x28 & n453 ) | ( ~n452 & n453 ) ;
  assign n455 = n452 & n454 ;
  assign n456 = ~x30 & n455 ;
  assign n464 = ~x21 & n46 ;
  assign n465 = x20 & n464 ;
  assign n470 = ~x28 & n465 ;
  assign n471 = x22 & n470 ;
  assign n472 = x30 & n471 ;
  assign n473 = x29 & n472 ;
  assign n466 = x28 & n465 ;
  assign n467 = x22 & n466 ;
  assign n468 = x30 & n467 ;
  assign n469 = x29 & n468 ;
  assign n474 = x1 & ~x20 ;
  assign n475 = ( x18 & x19 ) | ( x18 & n474 ) | ( x19 & n474 ) ;
  assign n476 = ~x18 & n475 ;
  assign n477 = ~x21 & n476 ;
  assign n478 = x23 & n477 ;
  assign n479 = ( x29 & x30 ) | ( x29 & n478 ) | ( x30 & n478 ) ;
  assign n480 = ~x30 & n479 ;
  assign n481 = n469 | n480 ;
  assign n482 = n473 | n481 ;
  assign n483 = n456 | n482 ;
  assign n484 = ( ~n449 & n463 ) | ( ~n449 & n483 ) | ( n463 & n483 ) ;
  assign n485 = n449 | n484 ;
  assign n416 = x41 & n390 ;
  assign n427 = x38 & n389 ;
  assign n417 = x9 & ~x19 ;
  assign n418 = ( x18 & ~x20 ) | ( x18 & n417 ) | ( ~x20 & n417 ) ;
  assign n419 = ~x18 & n418 ;
  assign n420 = x21 & n419 ;
  assign n421 = ( x22 & x28 ) | ( x22 & n420 ) | ( x28 & n420 ) ;
  assign n422 = ~x28 & n421 ;
  assign n423 = n49 & n422 ;
  assign n424 = ~x33 & x39 ;
  assign n425 = ( x31 & n423 ) | ( x31 & n424 ) | ( n423 & n424 ) ;
  assign n426 = ~x31 & n425 ;
  assign n429 = x18 & x19 ;
  assign n430 = ( x20 & x21 ) | ( x20 & n429 ) | ( x21 & n429 ) ;
  assign n431 = ~x21 & n430 ;
  assign n432 = x29 & n431 ;
  assign n433 = ( x27 & x28 ) | ( x27 & n432 ) | ( x28 & n432 ) ;
  assign n434 = ~x27 & n433 ;
  assign n435 = x30 & n434 ;
  assign n428 = n49 & n387 ;
  assign n436 = x27 & x30 ;
  assign n437 = ( x29 & n431 ) | ( x29 & n436 ) | ( n431 & n436 ) ;
  assign n438 = ~x29 & n437 ;
  assign n439 = n428 | n438 ;
  assign n440 = n435 | n439 ;
  assign n441 = n426 | n440 ;
  assign n442 = ( ~n416 & n427 ) | ( ~n416 & n441 ) | ( n427 & n441 ) ;
  assign n443 = n416 | n442 ;
  assign n492 = ~x29 & n431 ;
  assign n493 = ( x27 & x28 ) | ( x27 & n492 ) | ( x28 & n492 ) ;
  assign n494 = ~x27 & n493 ;
  assign n495 = ~x30 & n494 ;
  assign n486 = ( x18 & x20 ) | ( x18 & n246 ) | ( x20 & n246 ) ;
  assign n487 = ~x20 & n486 ;
  assign n488 = x28 & n487 ;
  assign n489 = x26 & n488 ;
  assign n490 = ~x30 & n489 ;
  assign n491 = x29 & n490 ;
  assign n500 = ( x29 & n212 ) | ( x29 & ~n487 ) | ( n212 & ~n487 ) ;
  assign n501 = n487 & n500 ;
  assign n496 = ~x28 & n487 ;
  assign n497 = x26 & n496 ;
  assign n498 = x30 & n497 ;
  assign n499 = x29 & n498 ;
  assign n502 = ( x29 & n221 ) | ( x29 & ~n487 ) | ( n221 & ~n487 ) ;
  assign n503 = n487 & n502 ;
  assign n504 = n499 | n503 ;
  assign n505 = n501 | n504 ;
  assign n506 = n491 | n505 ;
  assign n507 = n495 | n506 ;
  assign n508 = n443 | n507 ;
  assign n509 = ( ~n415 & n485 ) | ( ~n415 & n508 ) | ( n485 & n508 ) ;
  assign n510 = n415 | n509 ;
  assign n540 = ( ~x18 & x20 ) | ( ~x18 & n53 ) | ( x20 & n53 ) ;
  assign n541 = x18 & n540 ;
  assign n542 = ~x30 & n541 ;
  assign n543 = x29 & n542 ;
  assign n526 = x25 & x29 ;
  assign n544 = ( x11 & x19 ) | ( x11 & n141 ) | ( x19 & n141 ) ;
  assign n545 = ~x19 & n544 ;
  assign n546 = x21 & n545 ;
  assign n549 = ( x28 & n526 ) | ( x28 & n546 ) | ( n526 & n546 ) ;
  assign n550 = ~x28 & n549 ;
  assign n523 = ( x11 & x18 ) | ( x11 & n90 ) | ( x18 & n90 ) ;
  assign n524 = ~x11 & n523 ;
  assign n525 = x21 & n524 ;
  assign n551 = ( x28 & n453 ) | ( x28 & n525 ) | ( n453 & n525 ) ;
  assign n552 = ~x28 & n551 ;
  assign n553 = x30 & ~n552 ;
  assign n554 = ( n550 & n552 ) | ( n550 & ~n553 ) | ( n552 & ~n553 ) ;
  assign n547 = ( x28 & n453 ) | ( x28 & n546 ) | ( n453 & n546 ) ;
  assign n548 = ~x28 & n547 ;
  assign n555 = x22 & n477 ;
  assign n556 = ( x29 & x30 ) | ( x29 & n555 ) | ( x30 & n555 ) ;
  assign n557 = ~x30 & n556 ;
  assign n558 = ( x18 & ~x21 ) | ( x18 & n90 ) | ( ~x21 & n90 ) ;
  assign n559 = ~x18 & n558 ;
  assign n563 = x30 & n559 ;
  assign n564 = ( x28 & x29 ) | ( x28 & n563 ) | ( x29 & n563 ) ;
  assign n565 = ~x28 & n564 ;
  assign n560 = x28 & n559 ;
  assign n561 = ( x29 & x30 ) | ( x29 & n560 ) | ( x30 & n560 ) ;
  assign n562 = ~x30 & n561 ;
  assign n566 = x19 | x21 ;
  assign n567 = ( ~x18 & x20 ) | ( ~x18 & n566 ) | ( x20 & n566 ) ;
  assign n568 = x18 | n567 ;
  assign n569 = x30 & ~n568 ;
  assign n570 = ( x28 & x29 ) | ( x28 & n569 ) | ( x29 & n569 ) ;
  assign n571 = ~x28 & n570 ;
  assign n572 = x28 & ~n568 ;
  assign n573 = ( x29 & x30 ) | ( x29 & n572 ) | ( x30 & n572 ) ;
  assign n574 = ~x30 & n573 ;
  assign n575 = n571 | n574 ;
  assign n576 = n562 | n575 ;
  assign n577 = ( ~n557 & n565 ) | ( ~n557 & n576 ) | ( n565 & n576 ) ;
  assign n578 = n557 | n577 ;
  assign n579 = n548 | n578 ;
  assign n580 = ( ~n543 & n554 ) | ( ~n543 & n579 ) | ( n554 & n579 ) ;
  assign n581 = n543 | n580 ;
  assign n511 = x20 & n47 ;
  assign n512 = ( x28 & n400 ) | ( x28 & n511 ) | ( n400 & n511 ) ;
  assign n513 = ~x28 & n512 ;
  assign n514 = ~x30 & n513 ;
  assign n518 = ( x18 & x19 ) | ( x18 & n59 ) | ( x19 & n59 ) ;
  assign n519 = ~x19 & n518 ;
  assign n520 = ~x30 & n519 ;
  assign n521 = ( x28 & x29 ) | ( x28 & n520 ) | ( x29 & n520 ) ;
  assign n522 = ~x28 & n521 ;
  assign n515 = x28 & n47 ;
  assign n516 = ( x29 & x30 ) | ( x29 & n515 ) | ( x30 & n515 ) ;
  assign n517 = ~x30 & n516 ;
  assign n527 = ( x28 & n525 ) | ( x28 & n526 ) | ( n525 & n526 ) ;
  assign n528 = ~x28 & n527 ;
  assign n529 = ~x30 & n528 ;
  assign n530 = x18 & x21 ;
  assign n531 = ( x19 & x20 ) | ( x19 & n530 ) | ( x20 & n530 ) ;
  assign n532 = ~x19 & n531 ;
  assign n533 = ( x28 & n400 ) | ( x28 & n532 ) | ( n400 & n532 ) ;
  assign n534 = ~x28 & n533 ;
  assign n535 = ~x30 & n534 ;
  assign n536 = n529 | n535 ;
  assign n537 = n517 | n536 ;
  assign n538 = ( ~n514 & n522 ) | ( ~n514 & n537 ) | ( n522 & n537 ) ;
  assign n539 = n514 | n538 ;
  assign n582 = x21 & n476 ;
  assign n583 = ( x23 & x28 ) | ( x23 & n582 ) | ( x28 & n582 ) ;
  assign n584 = ~x28 & n583 ;
  assign n585 = n49 & n584 ;
  assign n586 = ( x18 & x20 ) | ( x18 & n397 ) | ( x20 & n397 ) ;
  assign n587 = ~x18 & n586 ;
  assign n591 = ~x30 & n587 ;
  assign n592 = ( x26 & x29 ) | ( x26 & n591 ) | ( x29 & n591 ) ;
  assign n593 = ~x26 & n592 ;
  assign n594 = x26 & n587 ;
  assign n595 = ( x29 & x30 ) | ( x29 & n594 ) | ( x30 & n594 ) ;
  assign n596 = ~x30 & n595 ;
  assign n597 = n593 | n596 ;
  assign n588 = x26 & x30 ;
  assign n589 = ( x29 & ~n587 ) | ( x29 & n588 ) | ( ~n587 & n588 ) ;
  assign n590 = n587 & n589 ;
  assign n598 = ( x22 & x28 ) | ( x22 & n582 ) | ( x28 & n582 ) ;
  assign n599 = ~x28 & n598 ;
  assign n600 = n49 & n599 ;
  assign n601 = x24 & n587 ;
  assign n602 = ( x29 & x30 ) | ( x29 & n601 ) | ( x30 & n601 ) ;
  assign n603 = ~x30 & n602 ;
  assign n604 = n600 | n603 ;
  assign n605 = n590 | n604 ;
  assign n606 = ( ~n585 & n597 ) | ( ~n585 & n605 ) | ( n597 & n605 ) ;
  assign n607 = n585 | n606 ;
  assign n608 = n539 | n607 ;
  assign n609 = ( ~n510 & n581 ) | ( ~n510 & n608 ) | ( n581 & n608 ) ;
  assign n610 = n510 | n609 ;
  assign n611 = ~x44 & n394 ;
  assign n612 = x43 & n611 ;
  assign n613 = ( x3 & x19 ) | ( x3 & n141 ) | ( x19 & n141 ) ;
  assign n614 = ~x3 & n613 ;
  assign n615 = ~x29 & n614 ;
  assign n616 = ( x21 & x27 ) | ( x21 & n615 ) | ( x27 & n615 ) ;
  assign n617 = ~x21 & n616 ;
  assign n618 = ~x30 & n617 ;
  assign n619 = n495 | n618 ;
  assign n620 = x28 & ~x30 ;
  assign n621 = ( x29 & n446 ) | ( x29 & n620 ) | ( n446 & n620 ) ;
  assign n622 = ~x29 & n621 ;
  assign n623 = ~x29 & n489 ;
  assign n624 = ~x30 & n623 ;
  assign n625 = n499 | n624 ;
  assign n626 = n473 | n625 ;
  assign n627 = ( ~n449 & n622 ) | ( ~n449 & n626 ) | ( n622 & n626 ) ;
  assign n628 = n449 | n627 ;
  assign n629 = n438 | n628 ;
  assign n630 = ( ~n612 & n619 ) | ( ~n612 & n629 ) | ( n619 & n629 ) ;
  assign n631 = n612 | n630 ;
  assign n672 = n543 | n571 ;
  assign n673 = n574 | n672 ;
  assign n674 = n562 | n673 ;
  assign n675 = n565 | n674 ;
  assign n632 = x30 & n513 ;
  assign n633 = ( x29 & ~n47 ) | ( x29 & n111 ) | ( ~n47 & n111 ) ;
  assign n634 = n47 & n633 ;
  assign n635 = n514 | n634 ;
  assign n636 = n517 | n635 ;
  assign n637 = x30 & n519 ;
  assign n638 = ( x28 & x29 ) | ( x28 & n637 ) | ( x29 & n637 ) ;
  assign n639 = ~x28 & n638 ;
  assign n640 = n528 | n534 ;
  assign n641 = n639 | n640 ;
  assign n642 = n522 | n641 ;
  assign n643 = ( ~n632 & n636 ) | ( ~n632 & n642 ) | ( n636 & n642 ) ;
  assign n644 = n632 | n643 ;
  assign n663 = n590 | n603 ;
  assign n651 = x23 & n46 ;
  assign n652 = ( x20 & x21 ) | ( x20 & n651 ) | ( x21 & n651 ) ;
  assign n653 = ~x20 & n652 ;
  assign n654 = ~x30 & n653 ;
  assign n655 = ( x28 & x29 ) | ( x28 & n654 ) | ( x29 & n654 ) ;
  assign n656 = ~x28 & n655 ;
  assign n645 = x22 & n46 ;
  assign n646 = ( x20 & x21 ) | ( x20 & n645 ) | ( x21 & n645 ) ;
  assign n647 = ~x20 & n646 ;
  assign n648 = ~x30 & n647 ;
  assign n649 = ( x28 & x29 ) | ( x28 & n648 ) | ( x29 & n648 ) ;
  assign n650 = ~x28 & n649 ;
  assign n657 = ( x29 & n56 ) | ( x29 & ~n587 ) | ( n56 & ~n587 ) ;
  assign n658 = n587 & n657 ;
  assign n659 = n600 | n658 ;
  assign n660 = n650 | n659 ;
  assign n661 = ( ~n585 & n656 ) | ( ~n585 & n660 ) | ( n656 & n660 ) ;
  assign n662 = n585 | n661 ;
  assign n664 = x30 & n587 ;
  assign n665 = ( x26 & x29 ) | ( x26 & n664 ) | ( x29 & n664 ) ;
  assign n666 = ~x26 & n665 ;
  assign n667 = n593 | n666 ;
  assign n668 = n596 | n667 ;
  assign n669 = n662 | n668 ;
  assign n670 = ( ~n644 & n663 ) | ( ~n644 & n669 ) | ( n663 & n669 ) ;
  assign n671 = n644 | n670 ;
  assign n676 = ~x30 & n550 ;
  assign n677 = n548 | n552 ;
  assign n678 = ( n550 & ~n676 ) | ( n550 & n677 ) | ( ~n676 & n677 ) ;
  assign n679 = n671 | n678 ;
  assign n680 = ( ~n631 & n675 ) | ( ~n631 & n679 ) | ( n675 & n679 ) ;
  assign n681 = n631 | n680 ;
  assign n688 = n435 | n618 ;
  assign n682 = n456 | n503 ;
  assign n683 = ( ~n499 & n501 ) | ( ~n499 & n682 ) | ( n501 & n682 ) ;
  assign n684 = n499 | n683 ;
  assign n685 = n491 | n624 ;
  assign n686 = n495 | n685 ;
  assign n687 = n684 | n686 ;
  assign n689 = ~x43 & n394 ;
  assign n690 = ~x44 & n689 ;
  assign n691 = n396 | n428 ;
  assign n692 = n690 | n691 ;
  assign n693 = n687 | n692 ;
  assign n694 = ( ~n438 & n688 ) | ( ~n438 & n693 ) | ( n688 & n693 ) ;
  assign n695 = n438 | n694 ;
  assign n730 = n463 | n482 ;
  assign n731 = ( ~n449 & n622 ) | ( ~n449 & n730 ) | ( n622 & n730 ) ;
  assign n732 = n449 | n731 ;
  assign n696 = x30 & n550 ;
  assign n699 = x30 & n528 ;
  assign n700 = n676 | n699 ;
  assign n697 = x30 & n534 ;
  assign n698 = n529 | n697 ;
  assign n701 = n535 | n639 ;
  assign n702 = n698 | n701 ;
  assign n703 = ( ~n696 & n700 ) | ( ~n696 & n702 ) | ( n700 & n702 ) ;
  assign n704 = n696 | n703 ;
  assign n718 = n517 | n656 ;
  assign n719 = n634 | n718 ;
  assign n720 = n632 | n719 ;
  assign n721 = ( ~n514 & n522 ) | ( ~n514 & n720 ) | ( n522 & n720 ) ;
  assign n722 = n514 | n721 ;
  assign n705 = x30 & n548 ;
  assign n710 = ( x19 & x20 ) | ( x19 & n243 ) | ( x20 & n243 ) ;
  assign n711 = ~x20 & n710 ;
  assign n712 = ( x25 & n105 ) | ( x25 & ~n711 ) | ( n105 & ~n711 ) ;
  assign n713 = n711 & n712 ;
  assign n706 = ( x18 & x20 ) | ( x18 & n53 ) | ( x20 & n53 ) ;
  assign n707 = ~x20 & n706 ;
  assign n708 = x30 & n707 ;
  assign n709 = x26 & n708 ;
  assign n714 = ( n548 & n552 ) | ( n548 & ~n553 ) | ( n552 & ~n553 ) ;
  assign n715 = n709 | n714 ;
  assign n716 = ( ~n705 & n713 ) | ( ~n705 & n715 ) | ( n713 & n715 ) ;
  assign n717 = n705 | n716 ;
  assign n723 = x29 & n587 ;
  assign n724 = n603 | n723 ;
  assign n725 = ( ~n650 & n658 ) | ( ~n650 & n724 ) | ( n658 & n724 ) ;
  assign n726 = n650 | n725 ;
  assign n727 = n717 | n726 ;
  assign n728 = ( ~n704 & n722 ) | ( ~n704 & n727 ) | ( n722 & n727 ) ;
  assign n729 = n704 | n728 ;
  assign n733 = x30 & n541 ;
  assign n734 = x29 & n733 ;
  assign n735 = n543 | n575 ;
  assign n736 = n734 | n735 ;
  assign n737 = n562 | n736 ;
  assign n738 = ( ~n557 & n565 ) | ( ~n557 & n737 ) | ( n565 & n737 ) ;
  assign n739 = n557 | n738 ;
  assign n740 = n729 | n739 ;
  assign n741 = ( ~n695 & n732 ) | ( ~n695 & n740 ) | ( n732 & n740 ) ;
  assign n742 = n695 | n741 ;
  assign n812 = ( x29 & n212 ) | ( x29 & n487 ) | ( n212 & n487 ) ;
  assign n813 = ~x29 & n812 ;
  assign n818 = n456 | n463 ;
  assign n814 = n49 & n447 ;
  assign n815 = n49 & n461 ;
  assign n816 = n814 | n815 ;
  assign n817 = n622 | n816 ;
  assign n819 = n49 & n497 ;
  assign n820 = ~x29 & n711 ;
  assign n821 = ( x21 & x25 ) | ( x21 & n820 ) | ( x25 & n820 ) ;
  assign n822 = ~x21 & n821 ;
  assign n823 = x30 & n822 ;
  assign n824 = n503 | n823 ;
  assign n825 = n501 | n824 ;
  assign n826 = n624 | n825 ;
  assign n827 = n819 | n826 ;
  assign n828 = n817 | n827 ;
  assign n829 = ( ~n813 & n818 ) | ( ~n813 & n828 ) | ( n818 & n828 ) ;
  assign n830 = n813 | n829 ;
  assign n780 = x3 & x20 ;
  assign n781 = ( x18 & x19 ) | ( x18 & n780 ) | ( x19 & n780 ) ;
  assign n782 = ~x18 & n781 ;
  assign n783 = x28 & n782 ;
  assign n784 = ( x21 & x22 ) | ( x21 & n783 ) | ( x22 & n783 ) ;
  assign n785 = ~x21 & n784 ;
  assign n786 = n49 & n785 ;
  assign n773 = ~x3 & x19 ;
  assign n774 = ( x2 & ~x18 ) | ( x2 & n773 ) | ( ~x18 & n773 ) ;
  assign n775 = ~x2 & n774 ;
  assign n776 = ( x21 & n182 ) | ( x21 & n775 ) | ( n182 & n775 ) ;
  assign n777 = ~x21 & n776 ;
  assign n778 = ( x29 & n111 ) | ( x29 & n777 ) | ( n111 & n777 ) ;
  assign n779 = ~x29 & n778 ;
  assign n787 = x30 & n452 ;
  assign n788 = x22 & n787 ;
  assign n789 = x23 & n787 ;
  assign n790 = n788 | n789 ;
  assign n791 = n779 | n790 ;
  assign n792 = ( ~n469 & n786 ) | ( ~n469 & n791 ) | ( n786 & n791 ) ;
  assign n793 = n469 | n792 ;
  assign n757 = n676 | n713 ;
  assign n758 = n585 | n757 ;
  assign n747 = ~x20 & n46 ;
  assign n748 = ~x21 & n747 ;
  assign n749 = ( x29 & n212 ) | ( x29 & n748 ) | ( n212 & n748 ) ;
  assign n750 = ~x29 & n749 ;
  assign n743 = x23 & ~x29 ;
  assign n744 = ( x28 & n559 ) | ( x28 & n743 ) | ( n559 & n743 ) ;
  assign n745 = ~x28 & n744 ;
  assign n746 = x30 & n745 ;
  assign n751 = ( x28 & n49 ) | ( x28 & ~n568 ) | ( n49 & ~n568 ) ;
  assign n752 = ~x28 & n751 ;
  assign n753 = n734 | n752 ;
  assign n754 = n709 | n753 ;
  assign n755 = n746 | n754 ;
  assign n756 = n750 | n755 ;
  assign n759 = x14 & ~x28 ;
  assign n760 = ( x27 & ~x29 ) | ( x27 & n759 ) | ( ~x29 & n759 ) ;
  assign n761 = ~x27 & n760 ;
  assign n762 = ~x30 & n761 ;
  assign n763 = x13 & ~x27 ;
  assign n764 = ( x14 & x21 ) | ( x14 & n763 ) | ( x21 & n763 ) ;
  assign n765 = ~x14 & n764 ;
  assign n766 = ~x29 & n765 ;
  assign n767 = ( x28 & ~x30 ) | ( x28 & n766 ) | ( ~x30 & n766 ) ;
  assign n768 = ~x28 & n767 ;
  assign n769 = n762 | n768 ;
  assign n770 = n756 | n769 ;
  assign n771 = ( ~n600 & n758 ) | ( ~n600 & n770 ) | ( n758 & n770 ) ;
  assign n772 = n600 | n771 ;
  assign n794 = x26 & ~x29 ;
  assign n795 = ( x28 & n465 ) | ( x28 & n794 ) | ( n465 & n794 ) ;
  assign n796 = ~x28 & n795 ;
  assign n797 = x30 & n796 ;
  assign n799 = ( x28 & n465 ) | ( x28 & n743 ) | ( n465 & n743 ) ;
  assign n800 = ~x28 & n799 ;
  assign n801 = x30 & n800 ;
  assign n798 = n49 & n471 ;
  assign n802 = x23 & x30 ;
  assign n803 = ( x29 & n748 ) | ( x29 & n802 ) | ( n748 & n802 ) ;
  assign n804 = ~x29 & n803 ;
  assign n805 = n480 | n804 ;
  assign n806 = n557 | n805 ;
  assign n807 = n798 | n806 ;
  assign n808 = ( ~n797 & n801 ) | ( ~n797 & n807 ) | ( n801 & n807 ) ;
  assign n809 = n797 | n808 ;
  assign n810 = n772 | n809 ;
  assign n811 = n793 | n810 ;
  assign n831 = ~x27 & n431 ;
  assign n832 = ~x28 & n831 ;
  assign n833 = n49 & n832 ;
  assign n834 = n435 | n833 ;
  assign n835 = n491 | n834 ;
  assign n836 = n426 | n835 ;
  assign n837 = n618 | n836 ;
  assign n838 = n811 | n837 ;
  assign n839 = ( ~n415 & n830 ) | ( ~n415 & n838 ) | ( n830 & n838 ) ;
  assign n840 = n415 | n839 ;
  assign n841 = x40 & ~x42 ;
  assign n842 = ( x41 & n391 ) | ( x41 & n841 ) | ( n391 & n841 ) ;
  assign n843 = ~x41 & n842 ;
  assign n844 = n403 | n843 ;
  assign n845 = n411 | n844 ;
  assign n860 = x33 & n423 ;
  assign n861 = n426 | n618 ;
  assign n862 = ( ~n416 & n860 ) | ( ~n416 & n861 ) | ( n860 & n861 ) ;
  assign n863 = n416 | n862 ;
  assign n847 = n557 | n709 ;
  assign n848 = ( ~n480 & n786 ) | ( ~n480 & n847 ) | ( n786 & n847 ) ;
  assign n849 = n480 | n848 ;
  assign n846 = n469 | n779 ;
  assign n850 = x30 & n552 ;
  assign n851 = n585 | n590 ;
  assign n852 = ( ~n632 & n634 ) | ( ~n632 & n851 ) | ( n634 & n851 ) ;
  assign n853 = n632 | n852 ;
  assign n854 = n850 | n853 ;
  assign n855 = ( n676 & ~n705 ) | ( n676 & n854 ) | ( ~n705 & n854 ) ;
  assign n856 = n705 | n855 ;
  assign n857 = n846 | n856 ;
  assign n858 = ( ~n622 & n849 ) | ( ~n622 & n857 ) | ( n849 & n857 ) ;
  assign n859 = n622 | n858 ;
  assign n864 = n501 | n818 ;
  assign n865 = n503 | n864 ;
  assign n866 = n435 | n865 ;
  assign n867 = n685 | n866 ;
  assign n868 = n859 | n867 ;
  assign n869 = ( ~n845 & n863 ) | ( ~n845 & n868 ) | ( n863 & n868 ) ;
  assign n870 = n845 | n869 ;
  assign n873 = x23 & n399 ;
  assign n874 = ( x29 & x30 ) | ( x29 & n873 ) | ( x30 & n873 ) ;
  assign n875 = ~x30 & n874 ;
  assign n876 = x31 & n875 ;
  assign n877 = ( x32 & n875 ) | ( x32 & n876 ) | ( n875 & n876 ) ;
  assign n871 = ( x29 & n399 ) | ( x29 & n802 ) | ( n399 & n802 ) ;
  assign n872 = ~x29 & n871 ;
  assign n878 = ~x32 & n875 ;
  assign n879 = ( x31 & ~x33 ) | ( x31 & n878 ) | ( ~x33 & n878 ) ;
  assign n880 = ~x31 & n879 ;
  assign n883 = x34 & n880 ;
  assign n884 = ( x35 & n880 ) | ( x35 & n883 ) | ( n880 & n883 ) ;
  assign n881 = ~x34 & n880 ;
  assign n882 = ~x35 & n881 ;
  assign n885 = ( ~x36 & n882 ) | ( ~x36 & n884 ) | ( n882 & n884 ) ;
  assign n886 = x37 & ~n885 ;
  assign n887 = ( x37 & n884 ) | ( x37 & ~n886 ) | ( n884 & ~n886 ) ;
  assign n888 = n872 | n887 ;
  assign n889 = ( ~n612 & n877 ) | ( ~n612 & n888 ) | ( n877 & n888 ) ;
  assign n890 = n612 | n889 ;
  assign n892 = x27 & x29 ;
  assign n893 = ( x28 & n431 ) | ( x28 & n892 ) | ( n431 & n892 ) ;
  assign n894 = ~x28 & n893 ;
  assign n895 = ~x30 & n894 ;
  assign n896 = ( x28 & n212 ) | ( x28 & ~n399 ) | ( n212 & ~n399 ) ;
  assign n897 = n399 & n896 ;
  assign n898 = n895 | n897 ;
  assign n891 = n273 | n438 ;
  assign n899 = ( ~x4 & x19 ) | ( ~x4 & n141 ) | ( x19 & n141 ) ;
  assign n900 = x4 & n899 ;
  assign n901 = ~x27 & x28 ;
  assign n902 = ( x21 & n900 ) | ( x21 & n901 ) | ( n900 & n901 ) ;
  assign n903 = ~x21 & n902 ;
  assign n904 = ~x30 & n903 ;
  assign n905 = x29 & n904 ;
  assign n906 = ( ~x5 & x19 ) | ( ~x5 & n141 ) | ( x19 & n141 ) ;
  assign n907 = x5 & n906 ;
  assign n908 = ~x27 & n907 ;
  assign n909 = ( x21 & ~x28 ) | ( x21 & n908 ) | ( ~x28 & n908 ) ;
  assign n910 = ~x21 & n909 ;
  assign n911 = x30 & n910 ;
  assign n912 = x29 & n911 ;
  assign n913 = n495 | n912 ;
  assign n914 = ( ~n435 & n905 ) | ( ~n435 & n913 ) | ( n905 & n913 ) ;
  assign n915 = n435 | n914 ;
  assign n916 = n891 | n915 ;
  assign n917 = ( ~n890 & n898 ) | ( ~n890 & n916 ) | ( n898 & n916 ) ;
  assign n918 = n890 | n917 ;
  assign n967 = ~x30 & n548 ;
  assign n969 = x3 & ~x18 ;
  assign n970 = ~x19 & n969 ;
  assign n971 = ~x21 & n970 ;
  assign n972 = ( x20 & ~x28 ) | ( x20 & n971 ) | ( ~x28 & n971 ) ;
  assign n973 = ~x20 & n972 ;
  assign n974 = ~x30 & n973 ;
  assign n975 = x29 & n974 ;
  assign n968 = ~x30 & n552 ;
  assign n976 = n543 | n968 ;
  assign n977 = ( ~n967 & n975 ) | ( ~n967 & n976 ) | ( n975 & n976 ) ;
  assign n978 = n967 | n977 ;
  assign n946 = n124 | n562 ;
  assign n947 = n750 | n946 ;
  assign n944 = ( x29 & n56 ) | ( x29 & n559 ) | ( n56 & n559 ) ;
  assign n945 = ~x29 & n944 ;
  assign n948 = x6 & ~x19 ;
  assign n949 = ( x3 & x18 ) | ( x3 & n948 ) | ( x18 & n948 ) ;
  assign n950 = ~x18 & n949 ;
  assign n951 = x20 & x28 ;
  assign n952 = ( x21 & n950 ) | ( x21 & n951 ) | ( n950 & n951 ) ;
  assign n953 = ~x21 & n952 ;
  assign n954 = n49 & n953 ;
  assign n955 = ~x3 & x6 ;
  assign n956 = ( x2 & ~x18 ) | ( x2 & n955 ) | ( ~x18 & n955 ) ;
  assign n957 = ~x2 & n956 ;
  assign n958 = ~x21 & n957 ;
  assign n959 = ( x19 & x20 ) | ( x19 & n958 ) | ( x20 & n958 ) ;
  assign n960 = ~x19 & n959 ;
  assign n961 = ( x29 & n111 ) | ( x29 & n960 ) | ( n111 & n960 ) ;
  assign n962 = ~x29 & n961 ;
  assign n963 = n954 | n962 ;
  assign n964 = n945 | n963 ;
  assign n965 = ( ~n565 & n947 ) | ( ~n565 & n964 ) | ( n947 & n964 ) ;
  assign n966 = n565 | n965 ;
  assign n979 = x5 & ~x18 ;
  assign n980 = ( x3 & ~x19 ) | ( x3 & n979 ) | ( ~x19 & n979 ) ;
  assign n981 = ~x3 & n980 ;
  assign n982 = ~x21 & n981 ;
  assign n983 = ( x20 & ~x28 ) | ( x20 & n982 ) | ( ~x28 & n982 ) ;
  assign n984 = ~x20 & n983 ;
  assign n985 = ~x30 & n984 ;
  assign n986 = x29 & n985 ;
  assign n987 = n574 | n986 ;
  assign n988 = ( ~n132 & n571 ) | ( ~n132 & n987 ) | ( n571 & n987 ) ;
  assign n989 = n132 | n988 ;
  assign n990 = n966 | n989 ;
  assign n991 = n978 | n990 ;
  assign n922 = ( x2 & x3 ) | ( x2 & n46 ) | ( x3 & n46 ) ;
  assign n923 = ~x3 & n922 ;
  assign n924 = ( x21 & n182 ) | ( x21 & n923 ) | ( n182 & n923 ) ;
  assign n925 = ~x21 & n924 ;
  assign n926 = ( x29 & n111 ) | ( x29 & n925 ) | ( n111 & n925 ) ;
  assign n927 = ~x29 & n926 ;
  assign n928 = n469 | n927 ;
  assign n929 = ( ~n449 & n814 ) | ( ~n449 & n928 ) | ( n814 & n928 ) ;
  assign n930 = n449 | n929 ;
  assign n919 = n499 | n865 ;
  assign n920 = ( ~n491 & n819 ) | ( ~n491 & n919 ) | ( n819 & n919 ) ;
  assign n921 = n491 | n920 ;
  assign n931 = x5 & x20 ;
  assign n932 = ( x18 & x19 ) | ( x18 & n931 ) | ( x19 & n931 ) ;
  assign n933 = ~x18 & n932 ;
  assign n934 = ~x28 & n933 ;
  assign n935 = ( x21 & x22 ) | ( x21 & n934 ) | ( x22 & n934 ) ;
  assign n936 = ~x21 & n935 ;
  assign n937 = ~x30 & n936 ;
  assign n938 = x29 & n937 ;
  assign n939 = n480 | n938 ;
  assign n940 = ( ~n473 & n557 ) | ( ~n473 & n939 ) | ( n557 & n939 ) ;
  assign n941 = n473 | n940 ;
  assign n942 = n921 | n941 ;
  assign n943 = n930 | n942 ;
  assign n997 = n517 | n585 ;
  assign n998 = n769 | n997 ;
  assign n999 = ( n597 & ~n604 ) | ( n597 & n998 ) | ( ~n604 & n998 ) ;
  assign n1000 = n604 | n999 ;
  assign n992 = ( x29 & n519 ) | ( x29 & n620 ) | ( n519 & n620 ) ;
  assign n993 = ~x29 & n992 ;
  assign n994 = n101 | n993 ;
  assign n995 = ( ~n514 & n522 ) | ( ~n514 & n994 ) | ( n522 & n994 ) ;
  assign n996 = n514 | n995 ;
  assign n1001 = n536 | n996 ;
  assign n1002 = ( ~n676 & n1000 ) | ( ~n676 & n1001 ) | ( n1000 & n1001 ) ;
  assign n1003 = n676 | n1002 ;
  assign n1004 = n943 | n1003 ;
  assign n1005 = ( ~n918 & n991 ) | ( ~n918 & n1004 ) | ( n991 & n1004 ) ;
  assign n1006 = n918 | n1005 ;
  assign n1009 = n403 | n408 ;
  assign n1007 = n405 | n416 ;
  assign n1008 = n411 | n1007 ;
  assign n1010 = n273 | n688 ;
  assign n1011 = n895 | n1010 ;
  assign n1012 = n427 | n1011 ;
  assign n1013 = ( ~n426 & n428 ) | ( ~n426 & n1012 ) | ( n428 & n1012 ) ;
  assign n1014 = n426 | n1013 ;
  assign n1015 = n1008 | n1014 ;
  assign n1016 = ( ~n396 & n1009 ) | ( ~n396 & n1015 ) | ( n1009 & n1015 ) ;
  assign n1017 = n396 | n1016 ;
  assign n1045 = n813 | n864 ;
  assign n1046 = n823 | n1045 ;
  assign n1047 = ( n503 & ~n819 ) | ( n503 & n1046 ) | ( ~n819 & n1046 ) ;
  assign n1048 = n819 | n1047 ;
  assign n1018 = n779 | n927 ;
  assign n1019 = n469 | n938 ;
  assign n1020 = n786 | n1019 ;
  assign n1021 = n797 | n801 ;
  assign n1022 = n557 | n1021 ;
  assign n1023 = ( ~n480 & n1020 ) | ( ~n480 & n1022 ) | ( n1020 & n1022 ) ;
  assign n1024 = n480 | n1023 ;
  assign n1025 = n817 | n1024 ;
  assign n1026 = ( ~n788 & n1018 ) | ( ~n788 & n1025 ) | ( n1018 & n1025 ) ;
  assign n1027 = n788 | n1026 ;
  assign n1033 = n124 | n963 ;
  assign n1028 = n967 | n975 ;
  assign n1029 = n968 | n1028 ;
  assign n1030 = n596 | n1029 ;
  assign n1031 = ( ~n676 & n769 ) | ( ~n676 & n1030 ) | ( n769 & n1030 ) ;
  assign n1032 = n676 | n1031 ;
  assign n1034 = ( x29 & n212 ) | ( x29 & n559 ) | ( n212 & n559 ) ;
  assign n1035 = ~x29 & n1034 ;
  assign n1036 = x24 & n559 ;
  assign n1037 = ( x29 & x30 ) | ( x29 & n1036 ) | ( x30 & n1036 ) ;
  assign n1038 = ~x30 & n1037 ;
  assign n1039 = n986 | n1038 ;
  assign n1040 = ( ~n132 & n1035 ) | ( ~n132 & n1039 ) | ( n1035 & n1039 ) ;
  assign n1041 = n132 | n1040 ;
  assign n1042 = n1032 | n1041 ;
  assign n1043 = ( ~n1027 & n1033 ) | ( ~n1027 & n1042 ) | ( n1033 & n1042 ) ;
  assign n1044 = n1027 | n1043 ;
  assign n1049 = n905 | n913 ;
  assign n1050 = ~x30 & n832 ;
  assign n1051 = x29 & n1050 ;
  assign n1052 = n833 | n1051 ;
  assign n1053 = n685 | n1052 ;
  assign n1054 = n1049 | n1053 ;
  assign n1055 = n1044 | n1054 ;
  assign n1056 = ( ~n1017 & n1048 ) | ( ~n1017 & n1055 ) | ( n1048 & n1055 ) ;
  assign n1057 = n1017 | n1056 ;
  assign n1058 = x36 & n882 ;
  assign n1059 = ( x37 & n882 ) | ( x37 & n1058 ) | ( n882 & n1058 ) ;
  assign n1060 = n843 | n897 ;
  assign n1061 = ( ~n690 & n860 ) | ( ~n690 & n1060 ) | ( n860 & n1060 ) ;
  assign n1062 = n690 | n1061 ;
  assign n1063 = n872 | n1062 ;
  assign n1064 = ( ~n612 & n1059 ) | ( ~n612 & n1063 ) | ( n1059 & n1063 ) ;
  assign n1065 = n612 | n1064 ;
  assign n1092 = n685 | n819 ;
  assign n1093 = ( ~n499 & n503 ) | ( ~n499 & n1092 ) | ( n503 & n1092 ) ;
  assign n1094 = n499 | n1093 ;
  assign n1095 = n438 | n895 ;
  assign n1096 = n1051 | n1095 ;
  assign n1097 = ( ~n435 & n1094 ) | ( ~n435 & n1096 ) | ( n1094 & n1096 ) ;
  assign n1098 = n435 | n1097 ;
  assign n1066 = ( x29 & n111 ) | ( x29 & n519 ) | ( n111 & n519 ) ;
  assign n1067 = ~x29 & n1066 ;
  assign n1068 = n639 | n698 ;
  assign n1069 = ( ~n535 & n1067 ) | ( ~n535 & n1068 ) | ( n1067 & n1068 ) ;
  assign n1070 = n535 | n1069 ;
  assign n1071 = n696 | n700 ;
  assign n1072 = ( ~n850 & n1070 ) | ( ~n850 & n1071 ) | ( n1070 & n1071 ) ;
  assign n1073 = n850 | n1072 ;
  assign n1085 = ( x22 & x30 ) | ( x22 & ~n707 ) | ( x30 & ~n707 ) ;
  assign n1086 = ( n705 & n707 ) | ( n705 & n1085 ) | ( n707 & n1085 ) ;
  assign n1087 = n709 | n1086 ;
  assign n1088 = n713 | n1087 ;
  assign n1074 = n659 | n663 ;
  assign n1077 = ( ~n585 & n650 ) | ( ~n585 & n718 ) | ( n650 & n718 ) ;
  assign n1078 = n585 | n1077 ;
  assign n1075 = n513 | n634 ;
  assign n1076 = n522 | n1075 ;
  assign n1079 = n596 | n769 ;
  assign n1080 = ( ~n593 & n666 ) | ( ~n593 & n1079 ) | ( n666 & n1079 ) ;
  assign n1081 = n593 | n1080 ;
  assign n1082 = n1076 | n1081 ;
  assign n1083 = ( ~n1074 & n1078 ) | ( ~n1074 & n1082 ) | ( n1078 & n1082 ) ;
  assign n1084 = n1074 | n1083 ;
  assign n1089 = n736 | n1084 ;
  assign n1090 = ( ~n1073 & n1088 ) | ( ~n1073 & n1089 ) | ( n1088 & n1089 ) ;
  assign n1091 = n1073 | n1090 ;
  assign n1105 = n473 | n786 ;
  assign n1099 = n463 | n501 ;
  assign n1100 = ( ~n456 & n622 ) | ( ~n456 & n1099 ) | ( n622 & n1099 ) ;
  assign n1101 = n456 | n1100 ;
  assign n1102 = n790 | n814 ;
  assign n1103 = ( ~n449 & n1101 ) | ( ~n449 & n1102 ) | ( n1101 & n1102 ) ;
  assign n1104 = n449 | n1103 ;
  assign n1106 = n562 | n945 ;
  assign n1107 = n565 | n1106 ;
  assign n1108 = n801 | n1107 ;
  assign n1109 = n750 | n1108 ;
  assign n1110 = n1104 | n1109 ;
  assign n1111 = ( ~n846 & n1105 ) | ( ~n846 & n1110 ) | ( n1105 & n1110 ) ;
  assign n1112 = n846 | n1111 ;
  assign n1113 = n1091 | n1112 ;
  assign n1114 = ( ~n1065 & n1098 ) | ( ~n1065 & n1113 ) | ( n1098 & n1113 ) ;
  assign n1115 = n1065 | n1114 ;
  assign n1116 = n571 | n752 ;
  assign n1117 = n574 | n1116 ;
  assign n1118 = n536 | n543 ;
  assign n1119 = n1117 | n1118 ;
  assign n1124 = n746 | n945 ;
  assign n1125 = n562 | n1124 ;
  assign n1126 = ( n565 & ~n750 ) | ( n565 & n1125 ) | ( ~n750 & n1125 ) ;
  assign n1127 = n750 | n1126 ;
  assign n1120 = n514 | n517 ;
  assign n1121 = n101 | n1120 ;
  assign n1122 = n522 | n1121 ;
  assign n1123 = n1067 | n1122 ;
  assign n1128 = n593 | n604 ;
  assign n1129 = ( ~n585 & n769 ) | ( ~n585 & n1128 ) | ( n769 & n1128 ) ;
  assign n1130 = n585 | n1129 ;
  assign n1131 = n1123 | n1130 ;
  assign n1132 = ( ~n1119 & n1127 ) | ( ~n1119 & n1131 ) | ( n1127 & n1131 ) ;
  assign n1133 = n1119 | n1132 ;
  assign n1144 = x18 & ~x20 ;
  assign n1145 = ( x10 & x19 ) | ( x10 & n1144 ) | ( x19 & n1144 ) ;
  assign n1146 = ~x19 & n1145 ;
  assign n1147 = x30 & n1146 ;
  assign n1148 = ( x21 & x25 ) | ( x21 & n1147 ) | ( x25 & n1147 ) ;
  assign n1149 = ~x21 & n1148 ;
  assign n1150 = n473 | n1149 ;
  assign n1151 = n788 | n1150 ;
  assign n1152 = n449 | n1151 ;
  assign n1153 = n815 | n1152 ;
  assign n1134 = n499 | n813 ;
  assign n1135 = n823 | n1134 ;
  assign n1136 = n833 | n1135 ;
  assign n1137 = ( n438 & ~n618 ) | ( n438 & n1136 ) | ( ~n618 & n1136 ) ;
  assign n1138 = n618 | n1137 ;
  assign n1139 = ( ~x34 & x35 ) | ( ~x34 & n895 ) | ( x35 & n895 ) ;
  assign n1140 = n880 | n895 ;
  assign n1141 = ( x34 & n1139 ) | ( x34 & n1140 ) | ( n1139 & n1140 ) ;
  assign n1142 = n1059 | n1141 ;
  assign n1143 = n1138 | n1142 ;
  assign n1154 = n809 | n1143 ;
  assign n1155 = ( ~n1133 & n1153 ) | ( ~n1133 & n1154 ) | ( n1153 & n1154 ) ;
  assign n1156 = n1133 | n1155 ;
  assign n1163 = n438 | n625 ;
  assign n1164 = ( n619 & ~n833 ) | ( n619 & n1163 ) | ( ~n833 & n1163 ) ;
  assign n1165 = n833 | n1164 ;
  assign n1157 = ~x34 & x35 ;
  assign n1158 = n880 & n1157 ;
  assign n1159 = ~x32 & x33 ;
  assign n1160 = ~x31 & n875 ;
  assign n1161 = ( x32 & n1159 ) | ( x32 & n1160 ) | ( n1159 & n1160 ) ;
  assign n1162 = n1158 | n1161 ;
  assign n1166 = n898 | n1162 ;
  assign n1167 = ( ~n612 & n1165 ) | ( ~n612 & n1166 ) | ( n1165 & n1166 ) ;
  assign n1168 = n612 | n1167 ;
  assign n1190 = n449 | n815 ;
  assign n1191 = n622 | n1190 ;
  assign n1192 = n823 | n1191 ;
  assign n1193 = ( n813 & ~n819 ) | ( n813 & n1192 ) | ( ~n819 & n1192 ) ;
  assign n1194 = n819 | n1193 ;
  assign n1178 = n565 | n746 ;
  assign n1179 = n562 | n1178 ;
  assign n1180 = n804 | n1179 ;
  assign n1181 = ( ~n480 & n750 ) | ( ~n480 & n1180 ) | ( n750 & n1180 ) ;
  assign n1182 = n480 | n1181 ;
  assign n1172 = n101 | n522 ;
  assign n1169 = n597 | n604 ;
  assign n1170 = ( ~n514 & n997 ) | ( ~n514 & n1169 ) | ( n997 & n1169 ) ;
  assign n1171 = n514 | n1170 ;
  assign n1173 = n529 | n967 ;
  assign n1174 = n968 | n1173 ;
  assign n1175 = n1171 | n1174 ;
  assign n1176 = ( ~n535 & n1172 ) | ( ~n535 & n1175 ) | ( n1172 & n1175 ) ;
  assign n1177 = n535 | n1176 ;
  assign n1183 = n574 | n1035 ;
  assign n1184 = n543 | n752 ;
  assign n1185 = n1038 | n1184 ;
  assign n1186 = ( ~n571 & n1183 ) | ( ~n571 & n1185 ) | ( n1183 & n1185 ) ;
  assign n1187 = n571 | n1186 ;
  assign n1188 = n1177 | n1187 ;
  assign n1189 = n1182 | n1188 ;
  assign n1195 = n789 | n814 ;
  assign n1196 = n779 | n1195 ;
  assign n1197 = n801 | n1196 ;
  assign n1198 = ( ~n798 & n1105 ) | ( ~n798 & n1197 ) | ( n1105 & n1197 ) ;
  assign n1199 = n798 | n1198 ;
  assign n1200 = n1189 | n1199 ;
  assign n1201 = ( ~n1168 & n1194 ) | ( ~n1168 & n1200 ) | ( n1194 & n1200 ) ;
  assign n1202 = n1168 | n1201 ;
  assign n1203 = n612 | n872 ;
  assign n1204 = n690 | n1203 ;
  assign n1205 = n396 | n843 ;
  assign n1206 = n897 | n1205 ;
  assign n1207 = ( ~n403 & n1204 ) | ( ~n403 & n1206 ) | ( n1204 & n1206 ) ;
  assign n1208 = n403 | n1207 ;
  assign n1212 = ( x31 & n875 ) | ( x31 & n1159 ) | ( n875 & n1159 ) ;
  assign n1213 = ~x31 & n1212 ;
  assign n1214 = x34 | n1213 ;
  assign n1215 = ( n880 & n1213 ) | ( n880 & n1214 ) | ( n1213 & n1214 ) ;
  assign n1209 = ( ~x36 & x37 ) | ( ~x36 & n1158 ) | ( x37 & n1158 ) ;
  assign n1210 = n882 | n1158 ;
  assign n1211 = ( x36 & n1209 ) | ( x36 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1216 = n877 | n1211 ;
  assign n1217 = ( ~n1208 & n1215 ) | ( ~n1208 & n1216 ) | ( n1215 & n1216 ) ;
  assign n1218 = n1208 | n1217 ;
  assign n1219 = n426 | n860 ;
  assign n1220 = ( ~n416 & n427 ) | ( ~n416 & n1219 ) | ( n427 & n1219 ) ;
  assign n1221 = n416 | n1220 ;
  assign n1222 = n495 | n688 ;
  assign n1223 = n905 | n1222 ;
  assign n1224 = n891 | n895 ;
  assign n1225 = ( ~n428 & n1223 ) | ( ~n428 & n1224 ) | ( n1223 & n1224 ) ;
  assign n1226 = n428 | n1225 ;
  assign n1227 = n413 | n1226 ;
  assign n1228 = ( ~n1218 & n1221 ) | ( ~n1218 & n1227 ) | ( n1221 & n1227 ) ;
  assign n1229 = n1218 | n1228 ;
  assign n1260 = n639 | n993 ;
  assign n1261 = n535 | n1260 ;
  assign n1262 = n1067 | n1261 ;
  assign n1263 = n632 | n1262 ;
  assign n1264 = ( ~n514 & n1172 ) | ( ~n514 & n1263 ) | ( n1172 & n1263 ) ;
  assign n1265 = n514 | n1264 ;
  assign n1266 = ~x10 & n138 ;
  assign n1267 = ~x15 & n1266 ;
  assign n1268 = ( x19 & n141 ) | ( x19 & n1267 ) | ( n141 & n1267 ) ;
  assign n1269 = ~x19 & n1268 ;
  assign n1270 = x21 & n1269 ;
  assign n1271 = ( x25 & x28 ) | ( x25 & n1270 ) | ( x28 & n1270 ) ;
  assign n1272 = ~x28 & n1271 ;
  assign n1273 = n49 & n1272 ;
  assign n1274 = x5 & ~x19 ;
  assign n1275 = ( x10 & x18 ) | ( x10 & n1274 ) | ( x18 & n1274 ) ;
  assign n1276 = ~x10 & n1275 ;
  assign n1277 = ( x21 & n153 ) | ( x21 & ~n1276 ) | ( n153 & ~n1276 ) ;
  assign n1278 = n1276 & n1277 ;
  assign n1279 = ( x28 & n49 ) | ( x28 & n1278 ) | ( n49 & n1278 ) ;
  assign n1280 = ~x28 & n1279 ;
  assign n1281 = n529 | n1280 ;
  assign n1282 = ( n697 & ~n1273 ) | ( n697 & n1281 ) | ( ~n1273 & n1281 ) ;
  assign n1283 = n1273 | n1282 ;
  assign n1284 = n700 | n1283 ;
  assign n1285 = ( ~n696 & n1265 ) | ( ~n696 & n1284 ) | ( n1265 & n1284 ) ;
  assign n1286 = n696 | n1285 ;
  assign n1287 = ~x10 & x19 ;
  assign n1288 = ~x18 & n1287 ;
  assign n1289 = x21 & n1288 ;
  assign n1290 = ( x25 & x28 ) | ( x25 & n1289 ) | ( x28 & n1289 ) ;
  assign n1291 = ~x28 & n1290 ;
  assign n1292 = n49 & n1291 ;
  assign n1293 = n600 | n1292 ;
  assign n1294 = ( ~n585 & n650 ) | ( ~n585 & n1293 ) | ( n650 & n1293 ) ;
  assign n1295 = n585 | n1294 ;
  assign n1296 = ( x10 & ~x19 ) | ( x10 & n74 ) | ( ~x19 & n74 ) ;
  assign n1297 = ~x10 & n1296 ;
  assign n1298 = x25 & n1297 ;
  assign n1299 = x21 & n1298 ;
  assign n1300 = n666 | n1299 ;
  assign n1301 = n590 | n658 ;
  assign n1302 = ( n596 & ~n603 ) | ( n596 & n1301 ) | ( ~n603 & n1301 ) ;
  assign n1303 = n603 | n1302 ;
  assign n1304 = n762 | n1303 ;
  assign n1305 = ( ~n593 & n1300 ) | ( ~n593 & n1304 ) | ( n1300 & n1304 ) ;
  assign n1306 = n593 | n1305 ;
  assign n1307 = n719 | n1306 ;
  assign n1308 = ( ~n1286 & n1295 ) | ( ~n1286 & n1307 ) | ( n1295 & n1307 ) ;
  assign n1309 = n1286 | n1308 ;
  assign n1230 = ~x10 & n1145 ;
  assign n1231 = ~x29 & n1230 ;
  assign n1232 = ( x21 & x25 ) | ( x21 & n1231 ) | ( x25 & n1231 ) ;
  assign n1233 = ~x21 & n1232 ;
  assign n1234 = x30 & n1233 ;
  assign n1235 = ( x30 & n822 ) | ( x30 & n1234 ) | ( n822 & n1234 ) ;
  assign n1236 = n499 | n685 ;
  assign n1237 = n819 | n1236 ;
  assign n1238 = n912 | n1237 ;
  assign n1239 = n1052 | n1238 ;
  assign n1240 = n1045 | n1239 ;
  assign n1241 = ( ~n503 & n1235 ) | ( ~n503 & n1240 ) | ( n1235 & n1240 ) ;
  assign n1242 = n503 | n1241 ;
  assign n1243 = n797 | n1105 ;
  assign n1244 = n938 | n1243 ;
  assign n1245 = n846 | n1149 ;
  assign n1246 = ( ~n927 & n1244 ) | ( ~n927 & n1245 ) | ( n1244 & n1245 ) ;
  assign n1247 = n927 | n1246 ;
  assign n1248 = x18 & ~x19 ;
  assign n1249 = ( x10 & ~x20 ) | ( x10 & n1248 ) | ( ~x20 & n1248 ) ;
  assign n1250 = ~x10 & n1249 ;
  assign n1251 = x30 & n1250 ;
  assign n1252 = ( x21 & x25 ) | ( x21 & n1251 ) | ( x25 & n1251 ) ;
  assign n1253 = ~x21 & n1252 ;
  assign n1254 = n788 | n1253 ;
  assign n1255 = ( n789 & ~n814 ) | ( n789 & n1254 ) | ( ~n814 & n1254 ) ;
  assign n1256 = n814 | n1255 ;
  assign n1257 = n1247 | n1256 ;
  assign n1258 = ( n1191 & ~n1242 ) | ( n1191 & n1257 ) | ( ~n1242 & n1257 ) ;
  assign n1259 = n1242 | n1258 ;
  assign n1310 = ( n734 & ~n975 ) | ( n734 & n1184 ) | ( ~n975 & n1184 ) ;
  assign n1311 = n975 | n1310 ;
  assign n1312 = n986 | n1311 ;
  assign n1313 = ( ~n132 & n571 ) | ( ~n132 & n1312 ) | ( n571 & n1312 ) ;
  assign n1314 = n132 | n1313 ;
  assign n1325 = n557 | n750 ;
  assign n1326 = ( ~n124 & n804 ) | ( ~n124 & n1325 ) | ( n804 & n1325 ) ;
  assign n1327 = n124 | n1326 ;
  assign n1328 = n801 | n1327 ;
  assign n1329 = ( n480 & ~n798 ) | ( n480 & n1328 ) | ( ~n798 & n1328 ) ;
  assign n1330 = n798 | n1329 ;
  assign n1315 = ( x25 & n105 ) | ( x25 & ~n1230 ) | ( n105 & ~n1230 ) ;
  assign n1316 = n1230 & n1315 ;
  assign n1317 = ( x22 & n707 ) | ( x22 & n713 ) | ( n707 & n713 ) ;
  assign n1318 = x30 & ~n1317 ;
  assign n1319 = ( x30 & n713 ) | ( x30 & ~n1318 ) | ( n713 & ~n1318 ) ;
  assign n1320 = n709 | n1319 ;
  assign n1321 = n1316 | n1320 ;
  assign n1322 = n968 | n1321 ;
  assign n1323 = ( n548 & ~n850 ) | ( n548 & n1322 ) | ( ~n850 & n1322 ) ;
  assign n1324 = n850 | n1323 ;
  assign n1331 = n945 | n1035 ;
  assign n1332 = n746 | n1038 ;
  assign n1333 = n1331 | n1332 ;
  assign n1334 = n962 | n1333 ;
  assign n1335 = ( n565 & ~n954 ) | ( n565 & n1334 ) | ( ~n954 & n1334 ) ;
  assign n1336 = n954 | n1335 ;
  assign n1337 = n1324 | n1336 ;
  assign n1338 = ( ~n1314 & n1330 ) | ( ~n1314 & n1337 ) | ( n1330 & n1337 ) ;
  assign n1339 = n1314 | n1338 ;
  assign n1340 = n1259 | n1339 ;
  assign n1341 = ( ~n1229 & n1309 ) | ( ~n1229 & n1340 ) | ( n1309 & n1340 ) ;
  assign n1342 = n1229 | n1341 ;
  assign n1343 = n596 | n967 ;
  assign n1344 = n968 | n1343 ;
  assign n1345 = n819 | n872 ;
  assign n1346 = n833 | n1345 ;
  assign n1347 = n813 | n1346 ;
  assign n1348 = ( ~n815 & n1235 ) | ( ~n815 & n1347 ) | ( n1235 & n1347 ) ;
  assign n1349 = n815 | n1348 ;
  assign n1350 = ( x19 & ~x21 ) | ( x19 & n1144 ) | ( ~x21 & n1144 ) ;
  assign n1351 = ~x19 & n1350 ;
  assign n1352 = x30 & n1351 ;
  assign n1353 = x22 & n1352 ;
  assign n1354 = n1149 | n1353 ;
  assign n1355 = n1256 | n1354 ;
  assign n1356 = ( ~n1021 & n1349 ) | ( ~n1021 & n1355 ) | ( n1349 & n1355 ) ;
  assign n1357 = n1021 | n1356 ;
  assign n1362 = ( x29 & n559 ) | ( x29 & n588 ) | ( n559 & n588 ) ;
  assign n1363 = ~x29 & n1362 ;
  assign n1364 = n746 | n1363 ;
  assign n1365 = n1331 | n1364 ;
  assign n1366 = n804 | n1365 ;
  assign n1367 = ( n750 & ~n798 ) | ( n750 & n1366 ) | ( ~n798 & n1366 ) ;
  assign n1368 = n798 | n1367 ;
  assign n1358 = x22 & n733 ;
  assign n1359 = n752 | n1358 ;
  assign n1360 = ( ~n1273 & n1316 ) | ( ~n1273 & n1359 ) | ( n1316 & n1359 ) ;
  assign n1361 = n1273 | n1360 ;
  assign n1369 = n1292 | n1299 ;
  assign n1370 = ( n768 & ~n1280 ) | ( n768 & n1369 ) | ( ~n1280 & n1369 ) ;
  assign n1371 = n1280 | n1370 ;
  assign n1372 = n1361 | n1371 ;
  assign n1373 = ( ~n1357 & n1368 ) | ( ~n1357 & n1372 ) | ( n1368 & n1372 ) ;
  assign n1374 = n1357 | n1373 ;
  assign n1375 = n746 | n752 ;
  assign n1376 = ( ~n798 & n833 ) | ( ~n798 & n1375 ) | ( n833 & n1375 ) ;
  assign n1377 = n798 | n1376 ;
  assign n1378 = n986 | n1033 ;
  assign n1379 = ( ~n132 & n975 ) | ( ~n132 & n1378 ) | ( n975 & n1378 ) ;
  assign n1380 = n132 | n1379 ;
  assign n1381 = n912 | n938 ;
  assign n1382 = n927 | n1381 ;
  assign n1383 = n905 | n1382 ;
  assign n1384 = ( ~n273 & n1380 ) | ( ~n273 & n1383 ) | ( n1380 & n1383 ) ;
  assign n1385 = n273 | n1384 ;
  assign n1402 = n650 | n658 ;
  assign n1403 = n1292 | n1402 ;
  assign n1411 = ( x7 & x16 ) | ( x7 & n46 ) | ( x16 & n46 ) ;
  assign n1412 = ~x16 & n1411 ;
  assign n1413 = ( x21 & n182 ) | ( x21 & ~n1412 ) | ( n182 & ~n1412 ) ;
  assign n1414 = n1412 & n1413 ;
  assign n1415 = ( x29 & n620 ) | ( x29 & n1414 ) | ( n620 & n1414 ) ;
  assign n1416 = ~x29 & n1415 ;
  assign n1404 = x16 & x19 ;
  assign n1405 = ( x8 & x18 ) | ( x8 & n1404 ) | ( x18 & n1404 ) ;
  assign n1406 = ~x18 & n1405 ;
  assign n1407 = ( x21 & n182 ) | ( x21 & ~n1406 ) | ( n182 & ~n1406 ) ;
  assign n1408 = n1406 & n1407 ;
  assign n1409 = ( x29 & n620 ) | ( x29 & n1408 ) | ( n620 & n1408 ) ;
  assign n1410 = ~x29 & n1409 ;
  assign n1417 = x21 & n933 ;
  assign n1418 = ( x22 & x28 ) | ( x22 & n1417 ) | ( x28 & n1417 ) ;
  assign n1419 = ~x28 & n1418 ;
  assign n1420 = n49 & n1419 ;
  assign n1421 = n634 | n1420 ;
  assign n1422 = n656 | n1421 ;
  assign n1423 = n1410 | n1422 ;
  assign n1424 = n1416 | n1423 ;
  assign n1425 = n1403 | n1424 ;
  assign n1426 = ( ~n590 & n1300 ) | ( ~n590 & n1425 ) | ( n1300 & n1425 ) ;
  assign n1427 = n590 | n1426 ;
  assign n1386 = n690 | n897 ;
  assign n1387 = ( n875 & ~n1160 ) | ( n875 & n1386 ) | ( ~n1160 & n1386 ) ;
  assign n1390 = n709 | n1316 ;
  assign n1391 = n713 | n1390 ;
  assign n1389 = n734 | n1358 ;
  assign n1392 = n1038 | n1363 ;
  assign n1393 = n1253 | n1392 ;
  assign n1394 = ( ~n1149 & n1353 ) | ( ~n1149 & n1393 ) | ( n1353 & n1393 ) ;
  assign n1395 = n1149 | n1394 ;
  assign n1396 = n1389 | n1395 ;
  assign n1397 = ( ~n1035 & n1391 ) | ( ~n1035 & n1396 ) | ( n1391 & n1396 ) ;
  assign n1398 = n1035 | n1397 ;
  assign n1388 = n882 | n884 ;
  assign n1399 = n1161 | n1388 ;
  assign n1400 = ( ~n1387 & n1398 ) | ( ~n1387 & n1399 ) | ( n1398 & n1399 ) ;
  assign n1401 = n1387 | n1400 ;
  assign n1435 = ( x5 & x19 ) | ( x5 & n141 ) | ( x19 & n141 ) ;
  assign n1436 = ~x19 & n1435 ;
  assign n1437 = x21 & ~x28 ;
  assign n1438 = ( x25 & n1436 ) | ( x25 & n1437 ) | ( n1436 & n1437 ) ;
  assign n1439 = ~x25 & n1438 ;
  assign n1440 = n49 & n1439 ;
  assign n1428 = x5 & x10 ;
  assign n1429 = ( x18 & x19 ) | ( x18 & n1428 ) | ( x19 & n1428 ) ;
  assign n1430 = ~x19 & n1429 ;
  assign n1431 = ( x21 & n153 ) | ( x21 & ~n1430 ) | ( n153 & ~n1430 ) ;
  assign n1432 = n1430 & n1431 ;
  assign n1433 = ( x28 & n49 ) | ( x28 & n1432 ) | ( n49 & n1432 ) ;
  assign n1434 = ~x28 & n1433 ;
  assign n1441 = n1067 | n1434 ;
  assign n1442 = n1440 | n1441 ;
  assign n1448 = x7 & ~x19 ;
  assign n1449 = ( x16 & x18 ) | ( x16 & n1448 ) | ( x18 & n1448 ) ;
  assign n1450 = ~x16 & n1449 ;
  assign n1451 = ( x21 & n951 ) | ( x21 & ~n1450 ) | ( n951 & ~n1450 ) ;
  assign n1452 = n1450 & n1451 ;
  assign n1443 = x8 & x16 ;
  assign n1444 = ( x18 & x19 ) | ( x18 & n1443 ) | ( x19 & n1443 ) ;
  assign n1445 = ~x19 & n1444 ;
  assign n1446 = ( x21 & n951 ) | ( x21 & ~n1445 ) | ( n951 & ~n1445 ) ;
  assign n1447 = n1445 & n1446 ;
  assign n1453 = n1086 | n1447 ;
  assign n1454 = ( ~n696 & n1452 ) | ( ~n696 & n1453 ) | ( n1452 & n1453 ) ;
  assign n1455 = n696 | n1454 ;
  assign n1456 = n1280 | n1455 ;
  assign n1457 = ( ~n1273 & n1442 ) | ( ~n1273 & n1456 ) | ( n1442 & n1456 ) ;
  assign n1458 = n1273 | n1457 ;
  assign n1459 = n1401 | n1458 ;
  assign n1460 = n1427 | n1459 ;
  assign n1470 = n257 | n265 ;
  assign n1471 = n273 | n1470 ;
  assign n1472 = n333 | n1471 ;
  assign n1473 = ( n124 & ~n318 ) | ( n124 & n1472 ) | ( ~n318 & n1472 ) ;
  assign n1474 = n318 | n1473 ;
  assign n1461 = n193 | n238 ;
  assign n1462 = n232 | n1461 ;
  assign n1463 = ( ~n95 & n224 ) | ( ~n95 & n1462 ) | ( n224 & n1462 ) ;
  assign n1464 = n95 | n1463 ;
  assign n1465 = n113 | n186 ;
  assign n1466 = n101 | n1465 ;
  assign n1467 = n209 | n1466 ;
  assign n1468 = ( ~n157 & n1464 ) | ( ~n157 & n1467 ) | ( n1464 & n1467 ) ;
  assign n1469 = n157 | n1468 ;
  assign n1475 = n132 | n173 ;
  assign n1476 = n137 | n1475 ;
  assign n1477 = n165 | n1476 ;
  assign n1478 = ( n107 & ~n147 ) | ( n107 & n1477 ) | ( ~n147 & n1477 ) ;
  assign n1479 = n147 | n1478 ;
  assign n1480 = n1469 | n1479 ;
  assign n1481 = n1474 | n1480 ;
  assign n1482 = n305 | n325 ;
  assign n1483 = n340 | n1482 ;
  assign n1484 = n251 | n312 ;
  assign n1485 = n281 | n1484 ;
  assign n1486 = n1483 | n1485 ;
  assign n1487 = n325 | n349 ;
  assign n1488 = n356 | n1487 ;
  assign n1489 = n281 | n297 ;
  assign n1490 = n1488 | n1489 ;
  assign n1491 = ~x13 & x21 ;
  assign n1492 = ( x12 & ~x14 ) | ( x12 & n1491 ) | ( ~x14 & n1491 ) ;
  assign n1493 = ~x12 & n1492 ;
  assign n1494 = ~x28 & n1493 ;
  assign n1495 = ( x27 & ~x29 ) | ( x27 & n1494 ) | ( ~x29 & n1494 ) ;
  assign n1496 = ~x27 & n1495 ;
  assign n1497 = ~x30 & n1496 ;
  assign n1498 = n891 | n905 ;
  assign n1499 = ( ~n435 & n912 ) | ( ~n435 & n1498 ) | ( n912 & n1498 ) ;
  assign n1500 = n435 | n1499 ;
  assign n1503 = n405 | n427 ;
  assign n1504 = n416 | n1503 ;
  assign n1501 = n396 | n845 ;
  assign n1502 = n612 | n1501 ;
  assign n1505 = x31 & n423 ;
  assign n1506 = ( ~x33 & n423 ) | ( ~x33 & n1505 ) | ( n423 & n1505 ) ;
  assign n1507 = n1502 | n1506 ;
  assign n1508 = n1504 | n1507 ;
  assign n1522 = n66 | n87 ;
  assign n1523 = n517 | n1522 ;
  assign n1524 = ( n113 & ~n632 ) | ( n113 & n1523 ) | ( ~n632 & n1523 ) ;
  assign n1525 = n632 | n1524 ;
  assign n1520 = n571 | n850 ;
  assign n1521 = n699 | n1520 ;
  assign n1526 = n1260 | n1521 ;
  assign n1527 = ( ~n697 & n1525 ) | ( ~n697 & n1526 ) | ( n1525 & n1526 ) ;
  assign n1528 = n697 | n1527 ;
  assign n1509 = n349 | n622 ;
  assign n1510 = n356 | n1509 ;
  assign n1511 = x30 & n494 ;
  assign n1512 = n265 | n495 ;
  assign n1513 = n296 | n1512 ;
  assign n1514 = n281 | n1513 ;
  assign n1515 = ( ~n860 & n1511 ) | ( ~n860 & n1514 ) | ( n1511 & n1514 ) ;
  assign n1516 = n860 | n1515 ;
  assign n1517 = n625 | n1516 ;
  assign n1518 = ( ~n290 & n1510 ) | ( ~n290 & n1517 ) | ( n1510 & n1517 ) ;
  assign n1519 = n290 | n1518 ;
  assign n1529 = ( x29 & n559 ) | ( x29 & n620 ) | ( n559 & n620 ) ;
  assign n1530 = ~x29 & n1529 ;
  assign n1531 = ( x29 & ~n568 ) | ( x29 & n620 ) | ( ~n568 & n620 ) ;
  assign n1532 = ~x29 & n1531 ;
  assign n1533 = n132 | n1532 ;
  assign n1534 = n565 | n1533 ;
  assign n1535 = n124 | n1534 ;
  assign n1536 = ( ~n473 & n1530 ) | ( ~n473 & n1535 ) | ( n1530 & n1535 ) ;
  assign n1537 = n473 | n1536 ;
  assign n1538 = ~x29 & n467 ;
  assign n1539 = ~x30 & n1538 ;
  assign n1540 = n786 | n1539 ;
  assign n1541 = n325 | n1540 ;
  assign n1542 = n779 | n1541 ;
  assign n1543 = ( ~n449 & n1537 ) | ( ~n449 & n1542 ) | ( n1537 & n1542 ) ;
  assign n1544 = n449 | n1543 ;
  assign n1545 = n1519 | n1544 ;
  assign n1546 = ( ~n1508 & n1528 ) | ( ~n1508 & n1545 ) | ( n1528 & n1545 ) ;
  assign n1547 = n1508 | n1546 ;
  assign n1548 = x3 | x18 ;
  assign n1549 = ( ~x2 & x6 ) | ( ~x2 & n1548 ) | ( x6 & n1548 ) ;
  assign n1550 = x2 | n1549 ;
  assign n1551 = x21 | n1550 ;
  assign n1552 = ( x19 & x20 ) | ( x19 & ~n1551 ) | ( x20 & ~n1551 ) ;
  assign n1553 = ~x19 & n1552 ;
  assign n1554 = ( x29 & n111 ) | ( x29 & n1553 ) | ( n111 & n1553 ) ;
  assign n1555 = ~x29 & n1554 ;
  assign n1556 = n124 | n1555 ;
  assign n1557 = n750 | n1556 ;
  assign n1558 = n469 | n786 ;
  assign n1559 = ( ~n318 & n325 ) | ( ~n318 & n1558 ) | ( n325 & n1558 ) ;
  assign n1560 = n318 | n1559 ;
  assign n1561 = n804 | n1560 ;
  assign n1562 = ( ~n798 & n1557 ) | ( ~n798 & n1561 ) | ( n1557 & n1561 ) ;
  assign n1563 = n798 | n1562 ;
  assign n1564 = n341 | n779 ;
  assign n1565 = ( ~n814 & n815 ) | ( ~n814 & n1564 ) | ( n815 & n1564 ) ;
  assign n1566 = n814 | n1565 ;
  assign n1567 = n305 | n813 ;
  assign n1568 = n1566 | n1567 ;
  assign n1569 = ( n357 & ~n1563 ) | ( n357 & n1568 ) | ( ~n1563 & n1568 ) ;
  assign n1570 = n1563 | n1569 ;
  assign n1574 = n257 | n819 ;
  assign n1575 = n312 | n1574 ;
  assign n1576 = ( ~n251 & n823 ) | ( ~n251 & n1575 ) | ( n823 & n1575 ) ;
  assign n1577 = n251 | n1576 ;
  assign n1578 = n1052 | n1577 ;
  assign n1579 = n297 | n1578 ;
  assign n1571 = n428 | n872 ;
  assign n1572 = ( ~n408 & n438 ) | ( ~n408 & n1571 ) | ( n438 & n1571 ) ;
  assign n1573 = n408 | n1572 ;
  assign n1580 = n905 | n1511 ;
  assign n1581 = n912 | n1580 ;
  assign n1582 = n281 | n1581 ;
  assign n1583 = n618 | n1582 ;
  assign n1584 = n1573 | n1583 ;
  assign n1585 = ( ~n1570 & n1579 ) | ( ~n1570 & n1584 ) | ( n1579 & n1584 ) ;
  assign n1586 = n1570 | n1585 ;
  assign n1595 = n214 | n593 ;
  assign n1596 = n193 | n604 ;
  assign n1597 = ( ~n95 & n596 ) | ( ~n95 & n1596 ) | ( n596 & n1596 ) ;
  assign n1598 = n95 | n1597 ;
  assign n1599 = n239 | n1598 ;
  assign n1600 = ( ~n223 & n1595 ) | ( ~n223 & n1599 ) | ( n1595 & n1599 ) ;
  assign n1601 = n223 | n1600 ;
  assign n1606 = n208 | n535 ;
  assign n1602 = n186 | n514 ;
  assign n1603 = n517 | n1602 ;
  assign n1604 = ( n113 & ~n585 ) | ( n113 & n1603 ) | ( ~n585 & n1603 ) ;
  assign n1605 = n585 | n1604 ;
  assign n1607 = n1172 | n1605 ;
  assign n1608 = ( ~n1601 & n1606 ) | ( ~n1601 & n1607 ) | ( n1606 & n1607 ) ;
  assign n1609 = n1601 | n1608 ;
  assign n1587 = n107 | n967 ;
  assign n1588 = ( ~n147 & n968 ) | ( ~n147 & n1587 ) | ( n968 & n1587 ) ;
  assign n1589 = n147 | n1588 ;
  assign n1590 = n157 | n529 ;
  assign n1591 = n201 | n1590 ;
  assign n1592 = n676 | n1591 ;
  assign n1593 = ( ~n165 & n1589 ) | ( ~n165 & n1592 ) | ( n1589 & n1592 ) ;
  assign n1594 = n165 | n1593 ;
  assign n1610 = ( x6 & ~x19 ) | ( x6 & n969 ) | ( ~x19 & n969 ) ;
  assign n1611 = ~x6 & n1610 ;
  assign n1612 = ( x21 & n951 ) | ( x21 & n1611 ) | ( n951 & n1611 ) ;
  assign n1613 = ~x21 & n1612 ;
  assign n1614 = n49 & n1613 ;
  assign n1615 = x3 | x19 ;
  assign n1616 = ( ~x2 & x18 ) | ( ~x2 & n1615 ) | ( x18 & n1615 ) ;
  assign n1617 = x2 | n1616 ;
  assign n1618 = x20 | n1617 ;
  assign n1619 = x21 | n1618 ;
  assign n1620 = ( x29 & n111 ) | ( x29 & ~n1619 ) | ( n111 & ~n1619 ) ;
  assign n1621 = ~x29 & n1620 ;
  assign n1622 = n173 | n1184 ;
  assign n1623 = ( ~n132 & n1621 ) | ( ~n132 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1624 = n132 | n1623 ;
  assign n1625 = n1614 | n1624 ;
  assign n1626 = ( ~n137 & n1124 ) | ( ~n137 & n1625 ) | ( n1124 & n1625 ) ;
  assign n1627 = n137 | n1626 ;
  assign n1628 = n1594 | n1627 ;
  assign n1629 = ( ~n1586 & n1609 ) | ( ~n1586 & n1628 ) | ( n1609 & n1628 ) ;
  assign n1630 = n1586 | n1629 ;
  assign n1631 = n495 | n1051 ;
  assign n1632 = n624 | n1631 ;
  assign n1633 = n273 | n618 ;
  assign n1634 = n281 | n1633 ;
  assign n1635 = n408 | n1634 ;
  assign n1636 = ( ~n843 & n860 ) | ( ~n843 & n1635 ) | ( n860 & n1635 ) ;
  assign n1637 = n843 | n1636 ;
  assign n1638 = n1484 | n1637 ;
  assign n1639 = ( ~n257 & n1632 ) | ( ~n257 & n1638 ) | ( n1632 & n1638 ) ;
  assign n1640 = n257 | n1639 ;
  assign n1661 = ( x14 & ~x20 ) | ( x14 & n1248 ) | ( ~x20 & n1248 ) ;
  assign n1662 = ~x14 & n1661 ;
  assign n1663 = ~x27 & n1662 ;
  assign n1664 = ( x21 & ~x28 ) | ( x21 & n1663 ) | ( ~x28 & n1663 ) ;
  assign n1665 = ~x21 & n1664 ;
  assign n1666 = ~x29 & n1665 ;
  assign n1667 = ~x30 & n1666 ;
  assign n1653 = ( x14 & ~x19 ) | ( x14 & n74 ) | ( ~x19 & n74 ) ;
  assign n1654 = ~x14 & n1653 ;
  assign n1655 = ~x23 & n1654 ;
  assign n1656 = ( x21 & ~x27 ) | ( x21 & n1655 ) | ( ~x27 & n1655 ) ;
  assign n1657 = ~x21 & n1656 ;
  assign n1658 = ~x29 & n1657 ;
  assign n1659 = ( x28 & ~x30 ) | ( x28 & n1658 ) | ( ~x30 & n1658 ) ;
  assign n1660 = ~x28 & n1659 ;
  assign n1668 = x13 & ~x21 ;
  assign n1669 = ( x14 & ~x27 ) | ( x14 & n1668 ) | ( ~x27 & n1668 ) ;
  assign n1670 = ~x14 & n1669 ;
  assign n1671 = ~x29 & n1670 ;
  assign n1672 = ( x28 & ~x30 ) | ( x28 & n1671 ) | ( ~x30 & n1671 ) ;
  assign n1673 = ~x28 & n1672 ;
  assign n1674 = n1660 | n1673 ;
  assign n1675 = ( ~n1497 & n1667 ) | ( ~n1497 & n1674 ) | ( n1667 & n1674 ) ;
  assign n1676 = n1497 | n1675 ;
  assign n1677 = ( x5 & x15 ) | ( x5 & n46 ) | ( x15 & n46 ) ;
  assign n1678 = ~x5 & n1677 ;
  assign n1679 = ( x21 & n182 ) | ( x21 & ~n1678 ) | ( n182 & ~n1678 ) ;
  assign n1680 = n1678 & n1679 ;
  assign n1681 = ( x28 & n49 ) | ( x28 & n1680 ) | ( n49 & n1680 ) ;
  assign n1682 = ~x28 & n1681 ;
  assign n1683 = ( ~n514 & n1523 ) | ( ~n514 & n1682 ) | ( n1523 & n1682 ) ;
  assign n1684 = n514 | n1683 ;
  assign n1685 = n1676 | n1684 ;
  assign n1686 = ( n597 & ~n603 ) | ( n597 & n1685 ) | ( ~n603 & n1685 ) ;
  assign n1687 = n603 | n1686 ;
  assign n1643 = n340 | n622 ;
  assign n1641 = n325 | n1539 ;
  assign n1642 = n333 | n1641 ;
  assign n1644 = n173 | n1532 ;
  assign n1645 = ( n543 & ~n967 ) | ( n543 & n1644 ) | ( ~n967 & n1644 ) ;
  assign n1646 = n967 | n1645 ;
  assign n1647 = n137 | n1646 ;
  assign n1648 = ( ~n318 & n1530 ) | ( ~n318 & n1647 ) | ( n1530 & n1647 ) ;
  assign n1649 = n318 | n1648 ;
  assign n1650 = n1642 | n1649 ;
  assign n1651 = ( ~n305 & n1643 ) | ( ~n305 & n1650 ) | ( n1643 & n1650 ) ;
  assign n1652 = n305 | n1651 ;
  assign n1700 = x15 & ~x19 ;
  assign n1701 = ( x5 & x18 ) | ( x5 & n1700 ) | ( x18 & n1700 ) ;
  assign n1702 = ~x5 & n1701 ;
  assign n1703 = x20 & n1702 ;
  assign n1704 = ( x21 & x28 ) | ( x21 & n1703 ) | ( x28 & n1703 ) ;
  assign n1705 = ~x28 & n1704 ;
  assign n1706 = n49 & n1705 ;
  assign n1713 = ~x16 & x19 ;
  assign n1714 = ( x7 & ~x18 ) | ( x7 & n1713 ) | ( ~x18 & n1713 ) ;
  assign n1715 = ~x7 & n1714 ;
  assign n1716 = ( x21 & n182 ) | ( x21 & ~n1715 ) | ( n182 & ~n1715 ) ;
  assign n1717 = n1715 & n1716 ;
  assign n1718 = ( x29 & n620 ) | ( x29 & n1717 ) | ( n620 & n1717 ) ;
  assign n1719 = ~x29 & n1718 ;
  assign n1707 = ( x8 & x16 ) | ( x8 & n46 ) | ( x16 & n46 ) ;
  assign n1708 = ~x8 & n1707 ;
  assign n1709 = ( x21 & n182 ) | ( x21 & ~n1708 ) | ( n182 & ~n1708 ) ;
  assign n1710 = n1708 & n1709 ;
  assign n1711 = ( x29 & n620 ) | ( x29 & n1710 ) | ( n620 & n1710 ) ;
  assign n1712 = ~x29 & n1711 ;
  assign n1720 = n522 | n1712 ;
  assign n1721 = n1719 | n1720 ;
  assign n1722 = n1706 | n1721 ;
  assign n1723 = ( ~n535 & n993 ) | ( ~n535 & n1722 ) | ( n993 & n1722 ) ;
  assign n1724 = n535 | n1723 ;
  assign n1688 = ~x16 & x18 ;
  assign n1689 = ( x7 & ~x19 ) | ( x7 & n1688 ) | ( ~x19 & n1688 ) ;
  assign n1690 = ~x7 & n1689 ;
  assign n1691 = ( x21 & n951 ) | ( x21 & ~n1690 ) | ( n951 & ~n1690 ) ;
  assign n1692 = n1690 & n1691 ;
  assign n1693 = x16 & ~x19 ;
  assign n1694 = ( x8 & x18 ) | ( x8 & n1693 ) | ( x18 & n1693 ) ;
  assign n1695 = ~x8 & n1694 ;
  assign n1696 = ( x21 & n951 ) | ( x21 & ~n1695 ) | ( n951 & ~n1695 ) ;
  assign n1697 = n1695 & n1696 ;
  assign n1698 = n529 | n1697 ;
  assign n1699 = n1692 | n1698 ;
  assign n1725 = n700 | n1699 ;
  assign n1726 = ( ~n968 & n1724 ) | ( ~n968 & n1725 ) | ( n1724 & n1725 ) ;
  assign n1727 = n968 | n1726 ;
  assign n1728 = n1652 | n1727 ;
  assign n1729 = ( ~n1640 & n1687 ) | ( ~n1640 & n1728 ) | ( n1687 & n1728 ) ;
  assign n1730 = n1640 | n1729 ;
  assign n1731 = n1204 | n1388 ;
  assign n1732 = ( n877 & ~n1213 ) | ( n877 & n1731 ) | ( ~n1213 & n1731 ) ;
  assign n1733 = n1213 | n1732 ;
  assign n1741 = n281 | n1511 ;
  assign n1742 = n905 | n1741 ;
  assign n1743 = ( x33 & n423 ) | ( x33 & n1505 ) | ( n423 & n1505 ) ;
  assign n1744 = n428 | n1095 ;
  assign n1745 = n1743 | n1744 ;
  assign n1746 = n688 | n1745 ;
  assign n1747 = ( ~n273 & n1742 ) | ( ~n273 & n1746 ) | ( n1742 & n1746 ) ;
  assign n1748 = n273 | n1747 ;
  assign n1734 = ~x31 & n423 ;
  assign n1735 = ~x33 & n1734 ;
  assign n1736 = n427 | n1735 ;
  assign n1737 = n1008 | n1736 ;
  assign n1738 = n1205 | n1737 ;
  assign n1739 = ( ~n897 & n1009 ) | ( ~n897 & n1738 ) | ( n1009 & n1738 ) ;
  assign n1740 = n897 | n1739 ;
  assign n1749 = n290 | n624 ;
  assign n1750 = n296 | n1749 ;
  assign n1751 = n491 | n1051 ;
  assign n1752 = n833 | n1751 ;
  assign n1753 = n495 | n1752 ;
  assign n1754 = ( ~n265 & n912 ) | ( ~n265 & n1753 ) | ( n912 & n1753 ) ;
  assign n1755 = n265 | n1754 ;
  assign n1756 = n1574 | n1755 ;
  assign n1757 = ( ~n499 & n1750 ) | ( ~n499 & n1756 ) | ( n1750 & n1756 ) ;
  assign n1758 = n499 | n1757 ;
  assign n1759 = n1740 | n1758 ;
  assign n1760 = ( ~n1733 & n1748 ) | ( ~n1733 & n1759 ) | ( n1748 & n1759 ) ;
  assign n1761 = n1733 | n1760 ;
  assign n1809 = n1033 | n1614 ;
  assign n1810 = ( n1530 & ~n1555 ) | ( n1530 & n1809 ) | ( ~n1555 & n1809 ) ;
  assign n1811 = n1555 | n1810 ;
  assign n1804 = n318 | n1539 ;
  assign n1805 = n473 | n1804 ;
  assign n1801 = n325 | n1018 ;
  assign n1802 = ( ~n469 & n786 ) | ( ~n469 & n1801 ) | ( n786 & n1801 ) ;
  assign n1803 = n469 | n1802 ;
  assign n1806 = n1021 | n1803 ;
  assign n1807 = ( ~n938 & n1805 ) | ( ~n938 & n1806 ) | ( n1805 & n1806 ) ;
  assign n1808 = n938 | n1807 ;
  assign n1812 = n557 | n562 ;
  assign n1813 = n750 | n1812 ;
  assign n1814 = n480 | n1813 ;
  assign n1815 = ( ~n798 & n804 ) | ( ~n798 & n1814 ) | ( n804 & n1814 ) ;
  assign n1816 = n798 | n1815 ;
  assign n1817 = n1808 | n1816 ;
  assign n1818 = n1811 | n1817 ;
  assign n1826 = n501 | n1567 ;
  assign n1827 = ( n357 & ~n456 ) | ( n357 & n1826 ) | ( ~n456 & n1826 ) ;
  assign n1828 = n456 | n1827 ;
  assign n1819 = n790 | n1253 ;
  assign n1820 = ( ~n814 & n1354 ) | ( ~n814 & n1819 ) | ( n1354 & n1819 ) ;
  assign n1821 = n814 | n1820 ;
  assign n1822 = n333 | n1190 ;
  assign n1823 = n1821 | n1822 ;
  assign n1824 = ( ~n463 & n1643 ) | ( ~n463 & n1823 ) | ( n1643 & n1823 ) ;
  assign n1825 = n463 | n1824 ;
  assign n1829 = n312 | n1235 ;
  assign n1830 = ( ~n251 & n503 ) | ( ~n251 & n1829 ) | ( n503 & n1829 ) ;
  assign n1831 = n251 | n1830 ;
  assign n1832 = n1825 | n1831 ;
  assign n1833 = ( ~n1818 & n1828 ) | ( ~n1818 & n1832 ) | ( n1828 & n1832 ) ;
  assign n1834 = n1818 | n1833 ;
  assign n1762 = n165 | n696 ;
  assign n1763 = n968 | n1762 ;
  assign n1764 = n676 | n1763 ;
  assign n1765 = ( ~n157 & n699 ) | ( ~n157 & n1764 ) | ( n699 & n1764 ) ;
  assign n1766 = n157 | n1765 ;
  assign n1772 = n967 | n1086 ;
  assign n1773 = ( ~n147 & n850 ) | ( ~n147 & n1772 ) | ( n850 & n1772 ) ;
  assign n1774 = n147 | n1773 ;
  assign n1767 = n201 | n1697 ;
  assign n1768 = n529 | n1767 ;
  assign n1769 = n1447 | n1768 ;
  assign n1770 = ( ~n1273 & n1452 ) | ( ~n1273 & n1769 ) | ( n1452 & n1769 ) ;
  assign n1771 = n1273 | n1770 ;
  assign n1775 = n697 | n1692 ;
  assign n1776 = n1706 | n1775 ;
  assign n1777 = n1434 | n1776 ;
  assign n1778 = ( ~n1280 & n1440 ) | ( ~n1280 & n1777 ) | ( n1440 & n1777 ) ;
  assign n1779 = n1280 | n1778 ;
  assign n1780 = n1771 | n1779 ;
  assign n1781 = ( ~n1766 & n1774 ) | ( ~n1766 & n1780 ) | ( n1774 & n1780 ) ;
  assign n1782 = n1766 | n1781 ;
  assign n1790 = n752 | n975 ;
  assign n1791 = n734 | n1790 ;
  assign n1792 = n986 | n1791 ;
  assign n1793 = ( ~n173 & n571 ) | ( ~n173 & n1792 ) | ( n571 & n1792 ) ;
  assign n1794 = n173 | n1793 ;
  assign n1783 = n1533 | n1621 ;
  assign n1784 = n746 | n1392 ;
  assign n1785 = ( ~n137 & n565 ) | ( ~n137 & n1784 ) | ( n565 & n1784 ) ;
  assign n1786 = n137 | n1785 ;
  assign n1787 = n1783 | n1786 ;
  assign n1788 = ( ~n945 & n1183 ) | ( ~n945 & n1787 ) | ( n1183 & n1787 ) ;
  assign n1789 = n945 | n1788 ;
  assign n1795 = n543 | n1391 ;
  assign n1796 = ( ~n107 & n1358 ) | ( ~n107 & n1795 ) | ( n1358 & n1795 ) ;
  assign n1797 = n107 | n1796 ;
  assign n1798 = n1789 | n1797 ;
  assign n1799 = ( ~n1782 & n1794 ) | ( ~n1782 & n1798 ) | ( n1794 & n1798 ) ;
  assign n1800 = n1782 | n1799 ;
  assign n1835 = n1172 | n1416 ;
  assign n1836 = n1712 | n1835 ;
  assign n1837 = ( ~n1410 & n1719 ) | ( ~n1410 & n1836 ) | ( n1719 & n1836 ) ;
  assign n1838 = n1410 | n1837 ;
  assign n1839 = n1606 | n1838 ;
  assign n1840 = ( ~n1067 & n1260 ) | ( ~n1067 & n1839 ) | ( n1260 & n1839 ) ;
  assign n1841 = n1067 | n1840 ;
  assign n1852 = n66 | n658 ;
  assign n1853 = n73 | n1852 ;
  assign n1854 = n95 | n590 ;
  assign n1855 = n603 | n1854 ;
  assign n1856 = n596 | n1461 ;
  assign n1857 = n1855 | n1856 ;
  assign n1858 = n600 | n1857 ;
  assign n1859 = ( ~n51 & n1853 ) | ( ~n51 & n1858 ) | ( n1853 & n1858 ) ;
  assign n1860 = n51 | n1859 ;
  assign n1842 = n585 | n1292 ;
  assign n1843 = n650 | n1842 ;
  assign n1844 = n656 | n1843 ;
  assign n1845 = ( n113 & ~n517 ) | ( n113 & n1844 ) | ( ~n517 & n1844 ) ;
  assign n1846 = n517 | n1845 ;
  assign n1847 = n634 | n1682 ;
  assign n1848 = n1420 | n1847 ;
  assign n1849 = n1846 | n1848 ;
  assign n1850 = ( ~n632 & n1602 ) | ( ~n632 & n1849 ) | ( n1602 & n1849 ) ;
  assign n1851 = n632 | n1850 ;
  assign n1861 = n223 | n1299 ;
  assign n1862 = n232 | n1861 ;
  assign n1863 = x26 & n105 ;
  assign n1864 = ( x19 & n141 ) | ( x19 & ~n1863 ) | ( n141 & ~n1863 ) ;
  assign n1865 = n1863 & n1864 ;
  assign n1866 = n1660 | n1865 ;
  assign n1867 = n762 | n1866 ;
  assign n1868 = n1667 | n1867 ;
  assign n1869 = ( ~n1497 & n1673 ) | ( ~n1497 & n1868 ) | ( n1673 & n1868 ) ;
  assign n1870 = n1497 | n1869 ;
  assign n1871 = n1595 | n1870 ;
  assign n1872 = ( ~n666 & n1862 ) | ( ~n666 & n1871 ) | ( n1862 & n1871 ) ;
  assign n1873 = n666 | n1872 ;
  assign n1874 = n1851 | n1873 ;
  assign n1875 = ( ~n1841 & n1860 ) | ( ~n1841 & n1874 ) | ( n1860 & n1874 ) ;
  assign n1876 = n1841 | n1875 ;
  assign n1877 = n1800 | n1876 ;
  assign n1878 = ( ~n1761 & n1834 ) | ( ~n1761 & n1877 ) | ( n1834 & n1877 ) ;
  assign n1879 = n1761 | n1878 ;
  assign n1880 = x21 & n49 ;
  assign n1881 = ( x18 & n90 ) | ( x18 & n1880 ) | ( n90 & n1880 ) ;
  assign n1882 = ~x18 & n1881 ;
  assign n1883 = ~x21 & x29 ;
  assign n1884 = ~x30 & n1883 ;
  assign n1885 = x18 & n1884 ;
  assign n1886 = ( x19 & x20 ) | ( x19 & n1885 ) | ( x20 & n1885 ) ;
  assign n1887 = ~x20 & n1886 ;
  assign n1888 = n1882 | n1887 ;
  assign n1889 = x25 & n1888 ;
  assign n1890 = ( x22 & n1888 ) | ( x22 & n1889 ) | ( n1888 & n1889 ) ;
  assign n1939 = ~x19 & x28 ;
  assign n1942 = x11 & x30 ;
  assign n1943 = ( x26 & ~n1939 ) | ( x26 & n1942 ) | ( ~n1939 & n1942 ) ;
  assign n1944 = n1939 & n1943 ;
  assign n1945 = ( x3 & x19 ) | ( x3 & n1944 ) | ( x19 & n1944 ) ;
  assign n1946 = x27 & ~n1945 ;
  assign n1947 = ( x27 & n1944 ) | ( x27 & ~n1946 ) | ( n1944 & ~n1946 ) ;
  assign n1948 = x18 & ~n1947 ;
  assign n1940 = ~x3 & x30 ;
  assign n1941 = x2 & n1940 ;
  assign n1949 = n1939 & n1941 ;
  assign n1950 = x18 | n1949 ;
  assign n1951 = ~n1948 & n1950 ;
  assign n1952 = ~x29 & n1951 ;
  assign n1925 = x22 & x28 ;
  assign n1926 = ( ~x5 & x22 ) | ( ~x5 & n1925 ) | ( x22 & n1925 ) ;
  assign n1927 = x19 & ~n1926 ;
  assign n1928 = x23 & ~x28 ;
  assign n1929 = x19 | n1928 ;
  assign n1930 = ~n1927 & n1929 ;
  assign n1931 = ( x18 & ~x30 ) | ( x18 & n1930 ) | ( ~x30 & n1930 ) ;
  assign n1919 = x4 | x27 ;
  assign n1920 = x19 & ~x28 ;
  assign n1921 = x19 & ~n1920 ;
  assign n1922 = ~n1919 & n1921 ;
  assign n1923 = ( x26 & ~n1920 ) | ( x26 & n1921 ) | ( ~n1920 & n1921 ) ;
  assign n1924 = ( ~x28 & n1922 ) | ( ~x28 & n1923 ) | ( n1922 & n1923 ) ;
  assign n1932 = ( x18 & x30 ) | ( x18 & ~n1924 ) | ( x30 & ~n1924 ) ;
  assign n1933 = n1931 & ~n1932 ;
  assign n1934 = ~x5 & x30 ;
  assign n1935 = ~x27 & n1934 ;
  assign n1936 = x18 & n1935 ;
  assign n1937 = ( x19 & x28 ) | ( x19 & n1936 ) | ( x28 & n1936 ) ;
  assign n1938 = ~x28 & n1937 ;
  assign n1953 = n1933 | n1938 ;
  assign n1954 = x29 & n1953 ;
  assign n1955 = n1952 | n1954 ;
  assign n1956 = x20 & n1955 ;
  assign n1904 = ( ~x26 & x28 ) | ( ~x26 & x29 ) | ( x28 & x29 ) ;
  assign n1905 = ( x29 & x30 ) | ( x29 & ~n1904 ) | ( x30 & ~n1904 ) ;
  assign n1906 = ( ~x28 & x30 ) | ( ~x28 & n1904 ) | ( x30 & n1904 ) ;
  assign n1907 = n1905 & ~n1906 ;
  assign n1915 = x19 & ~n46 ;
  assign n1916 = n1907 & n1915 ;
  assign n1910 = ~x28 & x29 ;
  assign n1911 = ( x5 & ~x30 ) | ( x5 & n1910 ) | ( ~x30 & n1910 ) ;
  assign n1912 = ~x5 & n1911 ;
  assign n1908 = ( x2 & x28 ) | ( x2 & n49 ) | ( x28 & n49 ) ;
  assign n1909 = ~x2 & n1908 ;
  assign n1913 = ~x3 & n1909 ;
  assign n1914 = ( ~x3 & n1912 ) | ( ~x3 & n1913 ) | ( n1912 & n1913 ) ;
  assign n1917 = ( ~n46 & n1914 ) | ( ~n46 & n1915 ) | ( n1914 & n1915 ) ;
  assign n1918 = ( ~x18 & n1916 ) | ( ~x18 & n1917 ) | ( n1916 & n1917 ) ;
  assign n1957 = x20 | n1918 ;
  assign n1958 = ( ~x20 & n1956 ) | ( ~x20 & n1957 ) | ( n1956 & n1957 ) ;
  assign n1959 = x21 | n1958 ;
  assign n1891 = x5 | x28 ;
  assign n1892 = x15 | n1891 ;
  assign n1893 = ( x20 & x22 ) | ( x20 & x28 ) | ( x22 & x28 ) ;
  assign n1894 = n1892 | n1893 ;
  assign n1895 = ( x28 & ~n1892 ) | ( x28 & n1894 ) | ( ~n1892 & n1894 ) ;
  assign n1896 = x19 & ~n1895 ;
  assign n1897 = x19 | n190 ;
  assign n1898 = ~n1896 & n1897 ;
  assign n1901 = ( x18 & ~x30 ) | ( x18 & n1898 ) | ( ~x30 & n1898 ) ;
  assign n1899 = ( x19 & n141 ) | ( x19 & ~n1892 ) | ( n141 & ~n1892 ) ;
  assign n1900 = ~x19 & n1899 ;
  assign n1902 = x30 & n1900 ;
  assign n1903 = ( n1898 & ~n1901 ) | ( n1898 & n1902 ) | ( ~n1901 & n1902 ) ;
  assign n1960 = ~x29 & n1903 ;
  assign n1961 = x21 & ~n1960 ;
  assign n1962 = n1959 & ~n1961 ;
  assign n1966 = ~x22 & x23 ;
  assign n1963 = x28 | x29 ;
  assign n1964 = x30 & n1963 ;
  assign n1965 = ( n105 & n1883 ) | ( n105 & ~n1964 ) | ( n1883 & ~n1964 ) ;
  assign n1967 = ~x20 & n1965 ;
  assign n1968 = ( x22 & n1966 ) | ( x22 & n1967 ) | ( n1966 & n1967 ) ;
  assign n1969 = ( x1 & n46 ) | ( x1 & n1968 ) | ( n46 & n1968 ) ;
  assign n1970 = ~x1 & n1969 ;
  assign n1971 = n63 | n1970 ;
  assign n1972 = ( ~n58 & n80 ) | ( ~n58 & n1971 ) | ( n80 & n1971 ) ;
  assign n1973 = n58 | n1972 ;
  assign n1974 = ( ~n1890 & n1962 ) | ( ~n1890 & n1973 ) | ( n1962 & n1973 ) ;
  assign n1975 = x0 & ~n1973 ;
  assign n1976 = ( n1890 & n1974 ) | ( n1890 & ~n1975 ) | ( n1974 & ~n1975 ) ;
  assign n1977 = n865 | n905 ;
  assign n1978 = ( n438 & ~n491 ) | ( n438 & n1977 ) | ( ~n491 & n1977 ) ;
  assign n1979 = n491 | n1978 ;
  assign n1980 = n522 | n529 ;
  assign n1981 = ( n535 & ~n676 ) | ( n535 & n1980 ) | ( ~n676 & n1980 ) ;
  assign n1982 = n676 | n1981 ;
  assign n1983 = n968 | n1982 ;
  assign n1984 = ( n543 & ~n967 ) | ( n543 & n1983 ) | ( ~n967 & n1983 ) ;
  assign n1985 = n967 | n1984 ;
  assign n1986 = n562 | n574 ;
  assign n1987 = ( ~n557 & n565 ) | ( ~n557 & n1986 ) | ( n565 & n1986 ) ;
  assign n1988 = n557 | n1987 ;
  assign n1989 = n927 | n1988 ;
  assign n1990 = ( ~n480 & n938 ) | ( ~n480 & n1989 ) | ( n938 & n1989 ) ;
  assign n1991 = n480 | n1990 ;
  assign n1992 = n1985 | n1991 ;
  assign n1993 = ( n1171 & ~n1979 ) | ( n1171 & n1992 ) | ( ~n1979 & n1992 ) ;
  assign n1994 = n1979 | n1993 ;
  assign n1995 = n1420 | n1440 ;
  assign n1996 = ( ~n975 & n1434 ) | ( ~n975 & n1995 ) | ( n1434 & n1995 ) ;
  assign n1997 = n975 | n1996 ;
  assign n1998 = n912 | n1997 ;
  assign n1999 = ( n938 & ~n986 ) | ( n938 & n1998 ) | ( ~n986 & n1998 ) ;
  assign n2000 = n986 | n1999 ;
  assign y0 = n85 ;
  assign y1 = n86 ;
  assign y2 = 1'b0 ;
  assign y3 = n87 ;
  assign y4 = n89 ;
  assign y5 = n116 ;
  assign y6 = n362 ;
  assign y7 = n367 ;
  assign y8 = n379 ;
  assign y9 = n381 ;
  assign y10 = n610 ;
  assign y11 = n681 ;
  assign y12 = n742 ;
  assign y13 = n840 ;
  assign y14 = n870 ;
  assign y15 = n1006 ;
  assign y16 = n1057 ;
  assign y17 = n1115 ;
  assign y18 = n1156 ;
  assign y19 = n1202 ;
  assign y20 = n463 ;
  assign y21 = n456 ;
  assign y22 = n1342 ;
  assign y23 = n1344 ;
  assign y24 = n1035 ;
  assign y25 = n1374 ;
  assign y26 = n1377 ;
  assign y27 = n1385 ;
  assign y28 = n1460 ;
  assign y29 = n1481 ;
  assign y30 = n1486 ;
  assign y31 = n1490 ;
  assign y32 = n1497 ;
  assign y33 = n1500 ;
  assign y34 = n1547 ;
  assign y35 = n1630 ;
  assign y36 = n1730 ;
  assign y37 = n1879 ;
  assign y38 = n1976 ;
  assign y39 = n1994 ;
  assign y40 = n2000 ;
  assign y41 = n186 ;
  assign y42 = 1'b0 ;
  assign y43 = n1331 ;
  assign y44 = n1035 ;
endmodule
