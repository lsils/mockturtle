module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 ;
  wire n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 ;
  assign n208 = x1 | x20 ;
  assign n209 = x107 & x163 ;
  assign n210 = ( ~x73 & x151 ) | ( ~x73 & n209 ) | ( x151 & n209 ) ;
  assign n211 = x73 & n210 ;
  assign n212 = x133 & x153 ;
  assign n213 = ( ~x75 & x141 ) | ( ~x75 & n212 ) | ( x141 & n212 ) ;
  assign n214 = x75 & n213 ;
  assign n215 = x106 & x109 ;
  assign n216 = ( ~x105 & x108 ) | ( ~x105 & n215 ) | ( x108 & n215 ) ;
  assign n217 = x105 & n216 ;
  assign n218 = x95 & x122 ;
  assign n219 = ( ~x85 & x111 ) | ( ~x85 & n218 ) | ( x111 & n218 ) ;
  assign n220 = x85 & n219 ;
  assign n221 = ~x1 & x165 ;
  assign n222 = ~x1 & x67 ;
  assign n223 = x66 & n222 ;
  assign n224 = x0 & x86 ;
  assign n225 = x5 & ~x152 ;
  assign n226 = ~x5 & x12 ;
  assign n227 = ( x5 & ~n225 ) | ( x5 & n226 ) | ( ~n225 & n226 ) ;
  assign n228 = ( x5 & x186 ) | ( x5 & n227 ) | ( x186 & n227 ) ;
  assign n229 = n227 & ~n228 ;
  assign n230 = ( x186 & ~n228 ) | ( x186 & n229 ) | ( ~n228 & n229 ) ;
  assign n231 = ~x205 & n230 ;
  assign n232 = x205 | n230 ;
  assign n233 = ( ~n230 & n231 ) | ( ~n230 & n232 ) | ( n231 & n232 ) ;
  assign n234 = x5 & ~x83 ;
  assign n235 = ~x5 & x69 ;
  assign n236 = ( x5 & ~n234 ) | ( x5 & n235 ) | ( ~n234 & n235 ) ;
  assign n237 = x177 | n236 ;
  assign n238 = ~x177 & n236 ;
  assign n239 = ( ~n236 & n237 ) | ( ~n236 & n238 ) | ( n237 & n238 ) ;
  assign n240 = x2 & x3 ;
  assign n241 = x80 & ~n240 ;
  assign n242 = ( x5 & n240 ) | ( x5 & ~n241 ) | ( n240 & ~n241 ) ;
  assign n243 = x180 | n242 ;
  assign n244 = ~x180 & n242 ;
  assign n245 = ( ~n242 & n243 ) | ( ~n242 & n244 ) | ( n243 & n244 ) ;
  assign n246 = x5 & ~x74 ;
  assign n247 = ~x5 & x72 ;
  assign n248 = ( x5 & ~n246 ) | ( x5 & n247 ) | ( ~n246 & n247 ) ;
  assign n249 = x176 | n248 ;
  assign n250 = ~x176 & n248 ;
  assign n251 = ( ~n248 & n249 ) | ( ~n248 & n250 ) | ( n249 & n250 ) ;
  assign n252 = x5 & ~x81 ;
  assign n253 = ~x5 & x68 ;
  assign n254 = ( x5 & ~n252 ) | ( x5 & n253 ) | ( ~n252 & n253 ) ;
  assign n255 = x179 | n254 ;
  assign n256 = ~x179 & n254 ;
  assign n257 = ( ~n254 & n255 ) | ( ~n254 & n256 ) | ( n255 & n256 ) ;
  assign n258 = x5 & ~x82 ;
  assign n259 = x5 | x71 ;
  assign n260 = ( x178 & n258 ) | ( x178 & ~n259 ) | ( n258 & ~n259 ) ;
  assign n261 = ( ~x178 & n259 ) | ( ~x178 & n260 ) | ( n259 & n260 ) ;
  assign n262 = ( ~n258 & n260 ) | ( ~n258 & n261 ) | ( n260 & n261 ) ;
  assign n263 = n257 | n262 ;
  assign n264 = ( n245 & n251 ) | ( n245 & n263 ) | ( n251 & n263 ) ;
  assign n265 = n245 & ~n264 ;
  assign n266 = ~n239 & n265 ;
  assign n267 = x76 & ~n240 ;
  assign n268 = ( x5 & n240 ) | ( x5 & ~n267 ) | ( n240 & ~n267 ) ;
  assign n269 = x184 | n268 ;
  assign n270 = ~x184 & n268 ;
  assign n271 = ( ~n268 & n269 ) | ( ~n268 & n270 ) | ( n269 & n270 ) ;
  assign n272 = x77 & ~n240 ;
  assign n273 = ( x5 & n240 ) | ( x5 & ~n272 ) | ( n240 & ~n272 ) ;
  assign n274 = x183 | n273 ;
  assign n275 = ~x183 & n273 ;
  assign n276 = ( ~n273 & n274 ) | ( ~n273 & n275 ) | ( n274 & n275 ) ;
  assign n277 = x78 & ~n240 ;
  assign n278 = ( x5 & n240 ) | ( x5 & ~n277 ) | ( n240 & ~n277 ) ;
  assign n279 = x182 | n278 ;
  assign n280 = ~x182 & n278 ;
  assign n281 = ( ~n278 & n279 ) | ( ~n278 & n280 ) | ( n279 & n280 ) ;
  assign n282 = x79 & ~n240 ;
  assign n283 = ( x5 & n240 ) | ( x5 & ~n282 ) | ( n240 & ~n282 ) ;
  assign n284 = x181 | n283 ;
  assign n285 = ~x181 & n283 ;
  assign n286 = ( ~n283 & n284 ) | ( ~n283 & n285 ) | ( n284 & n285 ) ;
  assign n287 = n281 & n286 ;
  assign n288 = ( ~n271 & n276 ) | ( ~n271 & n287 ) | ( n276 & n287 ) ;
  assign n289 = n271 & n288 ;
  assign n290 = n266 & n289 ;
  assign n291 = x5 & ~x158 ;
  assign n292 = ~x5 & x52 ;
  assign n293 = ( x5 & ~n291 ) | ( x5 & n292 ) | ( ~n291 & n292 ) ;
  assign n294 = x190 | n293 ;
  assign n295 = ~x190 & n293 ;
  assign n296 = ( ~n293 & n294 ) | ( ~n293 & n295 ) | ( n294 & n295 ) ;
  assign n297 = x5 & ~x161 ;
  assign n298 = ~x5 & x8 ;
  assign n299 = ( x5 & ~n297 ) | ( x5 & n298 ) | ( ~n297 & n298 ) ;
  assign n300 = x187 | n299 ;
  assign n301 = ~x187 & n299 ;
  assign n302 = ( ~n299 & n300 ) | ( ~n299 & n301 ) | ( n300 & n301 ) ;
  assign n303 = x5 & ~x160 ;
  assign n304 = ~x5 & x7 ;
  assign n305 = ( x5 & ~n303 ) | ( x5 & n304 ) | ( ~n303 & n304 ) ;
  assign n306 = x188 | n305 ;
  assign n307 = ~x188 & n305 ;
  assign n308 = ( ~n305 & n306 ) | ( ~n305 & n307 ) | ( n306 & n307 ) ;
  assign n309 = ~x186 & n227 ;
  assign n310 = ~x5 & n309 ;
  assign n311 = ~n308 & n310 ;
  assign n312 = ( n296 & ~n302 ) | ( n296 & n311 ) | ( ~n302 & n311 ) ;
  assign n313 = ~n296 & n312 ;
  assign n314 = x187 | n308 ;
  assign n315 = ( n296 & n299 ) | ( n296 & ~n314 ) | ( n299 & ~n314 ) ;
  assign n316 = ~n296 & n315 ;
  assign n317 = x5 & ~x159 ;
  assign n318 = ~x5 & x6 ;
  assign n319 = ( x5 & ~n317 ) | ( x5 & n318 ) | ( ~n317 & n318 ) ;
  assign n320 = ~x189 & n319 ;
  assign n321 = ( ~x190 & n293 ) | ( ~x190 & n320 ) | ( n293 & n320 ) ;
  assign n322 = x189 | n319 ;
  assign n323 = ( ~n319 & n320 ) | ( ~n319 & n322 ) | ( n320 & n322 ) ;
  assign n324 = ( n296 & ~n321 ) | ( n296 & n323 ) | ( ~n321 & n323 ) ;
  assign n325 = n307 & n324 ;
  assign n326 = ( n307 & n321 ) | ( n307 & ~n325 ) | ( n321 & ~n325 ) ;
  assign n327 = ( ~n313 & n316 ) | ( ~n313 & n326 ) | ( n316 & n326 ) ;
  assign n328 = n323 & ~n326 ;
  assign n329 = ( n313 & n327 ) | ( n313 & ~n328 ) | ( n327 & ~n328 ) ;
  assign n330 = x5 & ~x154 ;
  assign n331 = ~x5 & x51 ;
  assign n332 = ( x5 & ~n330 ) | ( x5 & n331 ) | ( ~n330 & n331 ) ;
  assign n333 = x194 | n332 ;
  assign n334 = ~x194 & n332 ;
  assign n335 = ( ~n332 & n333 ) | ( ~n332 & n334 ) | ( n333 & n334 ) ;
  assign n336 = x5 & ~x156 ;
  assign n337 = ~x5 & x64 ;
  assign n338 = ( x5 & ~n336 ) | ( x5 & n337 ) | ( ~n336 & n337 ) ;
  assign n339 = x192 | n338 ;
  assign n340 = ~x192 & n338 ;
  assign n341 = ( ~n338 & n339 ) | ( ~n338 & n340 ) | ( n339 & n340 ) ;
  assign n342 = x5 & ~x155 ;
  assign n343 = ~x5 & x63 ;
  assign n344 = ( x5 & ~n342 ) | ( x5 & n343 ) | ( ~n342 & n343 ) ;
  assign n345 = x193 | n344 ;
  assign n346 = ~x193 & n344 ;
  assign n347 = ( ~n344 & n345 ) | ( ~n344 & n346 ) | ( n345 & n346 ) ;
  assign n348 = x5 & ~x157 ;
  assign n349 = ~x5 & x65 ;
  assign n350 = ( x5 & ~n348 ) | ( x5 & n349 ) | ( ~n348 & n349 ) ;
  assign n351 = x191 | n350 ;
  assign n352 = ~x191 & n350 ;
  assign n353 = ( ~n350 & n351 ) | ( ~n350 & n352 ) | ( n351 & n352 ) ;
  assign n354 = n347 | n353 ;
  assign n355 = ( ~n335 & n341 ) | ( ~n335 & n354 ) | ( n341 & n354 ) ;
  assign n356 = n335 | n355 ;
  assign n357 = x5 & ~x149 ;
  assign n358 = ~x5 & x50 ;
  assign n359 = ( x5 & ~n357 ) | ( x5 & n358 ) | ( ~n357 & n358 ) ;
  assign n360 = x197 | n359 ;
  assign n361 = ~x197 & n359 ;
  assign n362 = ( ~n359 & n360 ) | ( ~n359 & n361 ) | ( n360 & n361 ) ;
  assign n363 = x5 & ~x146 ;
  assign n364 = ~x5 & x14 ;
  assign n365 = ( x5 & ~n363 ) | ( x5 & n364 ) | ( ~n363 & n364 ) ;
  assign n366 = x200 | n365 ;
  assign n367 = ~x200 & n365 ;
  assign n368 = ( ~n365 & n366 ) | ( ~n365 & n367 ) | ( n366 & n367 ) ;
  assign n369 = x5 & ~x140 ;
  assign n370 = ~x5 & x61 ;
  assign n371 = ( x5 & ~n369 ) | ( x5 & n370 ) | ( ~n369 & n370 ) ;
  assign n372 = x196 | n371 ;
  assign n373 = ~x196 & n371 ;
  assign n374 = ( ~n371 & n372 ) | ( ~n371 & n373 ) | ( n372 & n373 ) ;
  assign n375 = x5 & ~x147 ;
  assign n376 = ~x5 & x62 ;
  assign n377 = ( x5 & ~n375 ) | ( x5 & n376 ) | ( ~n375 & n376 ) ;
  assign n378 = x199 | n377 ;
  assign n379 = ~x199 & n377 ;
  assign n380 = ( ~n377 & n378 ) | ( ~n377 & n379 ) | ( n378 & n379 ) ;
  assign n381 = x5 & ~x148 ;
  assign n382 = x5 | x49 ;
  assign n383 = ( x198 & n381 ) | ( x198 & ~n382 ) | ( n381 & ~n382 ) ;
  assign n384 = ( ~x198 & n382 ) | ( ~x198 & n383 ) | ( n382 & n383 ) ;
  assign n385 = ( ~n381 & n383 ) | ( ~n381 & n384 ) | ( n383 & n384 ) ;
  assign n386 = n380 | n385 ;
  assign n387 = ( ~n368 & n374 ) | ( ~n368 & n386 ) | ( n374 & n386 ) ;
  assign n388 = n368 | n387 ;
  assign n389 = n362 | n388 ;
  assign n390 = x5 & ~x142 ;
  assign n391 = ~x5 & x29 ;
  assign n392 = ( x5 & ~n390 ) | ( x5 & n391 ) | ( ~n390 & n391 ) ;
  assign n393 = x204 | n392 ;
  assign n394 = ~x204 & n392 ;
  assign n395 = ( ~n392 & n393 ) | ( ~n392 & n394 ) | ( n393 & n394 ) ;
  assign n396 = x5 & ~x143 ;
  assign n397 = ~x5 & x15 ;
  assign n398 = ( x5 & ~n396 ) | ( x5 & n397 ) | ( ~n396 & n397 ) ;
  assign n399 = x203 | n398 ;
  assign n400 = ~x203 & n398 ;
  assign n401 = ( ~n398 & n399 ) | ( ~n398 & n400 ) | ( n399 & n400 ) ;
  assign n402 = x5 & ~x144 ;
  assign n403 = ~x5 & x9 ;
  assign n404 = ( x5 & ~n402 ) | ( x5 & n403 ) | ( ~n402 & n403 ) ;
  assign n405 = x202 | n404 ;
  assign n406 = ~x202 & n404 ;
  assign n407 = ( ~n404 & n405 ) | ( ~n404 & n406 ) | ( n405 & n406 ) ;
  assign n408 = x5 & ~x145 ;
  assign n409 = ~x5 & x10 ;
  assign n410 = ( x5 & ~n408 ) | ( x5 & n409 ) | ( ~n408 & n409 ) ;
  assign n411 = x201 | n410 ;
  assign n412 = ~x201 & n410 ;
  assign n413 = ( ~n410 & n411 ) | ( ~n410 & n412 ) | ( n411 & n412 ) ;
  assign n414 = n407 | n413 ;
  assign n415 = ( ~n395 & n401 ) | ( ~n395 & n414 ) | ( n401 & n414 ) ;
  assign n416 = n395 | n415 ;
  assign n417 = n389 | n416 ;
  assign n418 = ( n329 & n356 ) | ( n329 & n417 ) | ( n356 & n417 ) ;
  assign n419 = ( n335 & n340 ) | ( n335 & ~n347 ) | ( n340 & ~n347 ) ;
  assign n420 = ~n335 & n352 ;
  assign n421 = ~n341 & n420 ;
  assign n422 = ~n347 & n421 ;
  assign n423 = ( ~n335 & n419 ) | ( ~n335 & n422 ) | ( n419 & n422 ) ;
  assign n424 = ( ~x194 & n332 ) | ( ~x194 & n346 ) | ( n332 & n346 ) ;
  assign n425 = n423 | n424 ;
  assign n426 = ~n417 & n425 ;
  assign n427 = ( n329 & ~n418 ) | ( n329 & n426 ) | ( ~n418 & n426 ) ;
  assign n428 = n290 & n427 ;
  assign n429 = n308 | n323 ;
  assign n430 = ( ~n230 & n296 ) | ( ~n230 & n429 ) | ( n296 & n429 ) ;
  assign n431 = n230 | n430 ;
  assign n432 = n302 | n431 ;
  assign n433 = x205 & ~n432 ;
  assign n434 = ( ~n356 & n417 ) | ( ~n356 & n433 ) | ( n417 & n433 ) ;
  assign n435 = ~n417 & n434 ;
  assign n436 = n290 & n435 ;
  assign n437 = ~n368 & n373 ;
  assign n438 = ( n362 & ~n385 ) | ( n362 & n437 ) | ( ~n385 & n437 ) ;
  assign n439 = ~n362 & n438 ;
  assign n440 = ( n361 & n368 ) | ( n361 & ~n385 ) | ( n368 & ~n385 ) ;
  assign n441 = ~n368 & n440 ;
  assign n442 = ( x5 & x49 ) | ( x5 & ~x198 ) | ( x49 & ~x198 ) ;
  assign n443 = ( x5 & ~x148 ) | ( x5 & x198 ) | ( ~x148 & x198 ) ;
  assign n444 = n442 & ~n443 ;
  assign n445 = ( ~x200 & n365 ) | ( ~x200 & n379 ) | ( n365 & n379 ) ;
  assign n446 = ( n368 & n380 ) | ( n368 & ~n445 ) | ( n380 & ~n445 ) ;
  assign n447 = n444 & n446 ;
  assign n448 = ( n444 & n445 ) | ( n444 & ~n447 ) | ( n445 & ~n447 ) ;
  assign n449 = ( ~n439 & n441 ) | ( ~n439 & n448 ) | ( n441 & n448 ) ;
  assign n450 = n380 & ~n448 ;
  assign n451 = ( n439 & n449 ) | ( n439 & ~n450 ) | ( n449 & ~n450 ) ;
  assign n452 = ( n395 & ~n401 ) | ( n395 & n406 ) | ( ~n401 & n406 ) ;
  assign n453 = ~n395 & n412 ;
  assign n454 = ~n407 & n453 ;
  assign n455 = ~n401 & n454 ;
  assign n456 = ( ~n395 & n452 ) | ( ~n395 & n455 ) | ( n452 & n455 ) ;
  assign n457 = ( ~x204 & n392 ) | ( ~x204 & n400 ) | ( n392 & n400 ) ;
  assign n458 = n456 | n457 ;
  assign n459 = n416 & ~n458 ;
  assign n460 = ( n451 & n458 ) | ( n451 & ~n459 ) | ( n458 & ~n459 ) ;
  assign n461 = n290 & n460 ;
  assign n462 = ~n239 & n250 ;
  assign n463 = ( n245 & n262 ) | ( n245 & ~n462 ) | ( n262 & ~n462 ) ;
  assign n464 = n245 & ~n463 ;
  assign n465 = ( ~n238 & n245 ) | ( ~n238 & n262 ) | ( n245 & n262 ) ;
  assign n466 = n245 & ~n465 ;
  assign n467 = ( x5 & x71 ) | ( x5 & ~x178 ) | ( x71 & ~x178 ) ;
  assign n468 = ( x5 & ~x82 ) | ( x5 & x178 ) | ( ~x82 & x178 ) ;
  assign n469 = n467 & ~n468 ;
  assign n470 = ( x180 & n242 ) | ( x180 & ~n256 ) | ( n242 & ~n256 ) ;
  assign n471 = ( ~n245 & n257 ) | ( ~n245 & n470 ) | ( n257 & n470 ) ;
  assign n472 = n469 & n471 ;
  assign n473 = ( ~n469 & n470 ) | ( ~n469 & n472 ) | ( n470 & n472 ) ;
  assign n474 = ( n464 & ~n466 ) | ( n464 & n473 ) | ( ~n466 & n473 ) ;
  assign n475 = n257 & n473 ;
  assign n476 = ( ~n464 & n474 ) | ( ~n464 & n475 ) | ( n474 & n475 ) ;
  assign n477 = ( n271 & ~n276 ) | ( n271 & n279 ) | ( ~n276 & n279 ) ;
  assign n478 = n281 & ~n283 ;
  assign n479 = ( x181 & n271 ) | ( x181 & ~n478 ) | ( n271 & ~n478 ) ;
  assign n480 = n271 & ~n479 ;
  assign n481 = n276 & n480 ;
  assign n482 = ( n271 & ~n477 ) | ( n271 & n481 ) | ( ~n477 & n481 ) ;
  assign n483 = ( x184 & n268 ) | ( x184 & n274 ) | ( n268 & n274 ) ;
  assign n484 = ~n482 & n483 ;
  assign n485 = ~n289 & n484 ;
  assign n486 = ( n476 & n484 ) | ( n476 & n485 ) | ( n484 & n485 ) ;
  assign n487 = x139 & ~n240 ;
  assign n488 = ( x5 & n240 ) | ( x5 & ~n487 ) | ( n240 & ~n487 ) ;
  assign n489 = x169 | n488 ;
  assign n490 = ~x169 & n488 ;
  assign n491 = ( ~n488 & n489 ) | ( ~n488 & n490 ) | ( n489 & n490 ) ;
  assign n492 = x138 & ~n240 ;
  assign n493 = ( x5 & n240 ) | ( x5 & ~n492 ) | ( n240 & ~n492 ) ;
  assign n494 = ~x53 & n493 ;
  assign n495 = x53 | n493 ;
  assign n496 = ( ~n493 & n494 ) | ( ~n493 & n495 ) | ( n494 & n495 ) ;
  assign n497 = x136 & ~n240 ;
  assign n498 = ( x5 & n240 ) | ( x5 & ~n497 ) | ( n240 & ~n497 ) ;
  assign n499 = x171 | n498 ;
  assign n500 = ~x171 & n498 ;
  assign n501 = ( ~n498 & n499 ) | ( ~n498 & n500 ) | ( n499 & n500 ) ;
  assign n502 = x132 & ~n240 ;
  assign n503 = ( x5 & n240 ) | ( x5 & ~n502 ) | ( n240 & ~n502 ) ;
  assign n504 = x168 | n503 ;
  assign n505 = n501 & ~n504 ;
  assign n506 = ( ~n491 & n496 ) | ( ~n491 & n505 ) | ( n496 & n505 ) ;
  assign n507 = n491 & n506 ;
  assign n508 = ~n488 & n496 ;
  assign n509 = ( x169 & n501 ) | ( x169 & ~n508 ) | ( n501 & ~n508 ) ;
  assign n510 = n501 & ~n509 ;
  assign n511 = x5 & x138 ;
  assign n512 = x53 | n240 ;
  assign n513 = ( x5 & ~n511 ) | ( x5 & n512 ) | ( ~n511 & n512 ) ;
  assign n514 = x137 & ~n240 ;
  assign n515 = ( x5 & n240 ) | ( x5 & ~n514 ) | ( n240 & ~n514 ) ;
  assign n516 = x170 | n515 ;
  assign n517 = ( x171 & n498 ) | ( x171 & n516 ) | ( n498 & n516 ) ;
  assign n518 = ~x170 & n515 ;
  assign n519 = ( ~n515 & n516 ) | ( ~n515 & n518 ) | ( n516 & n518 ) ;
  assign n520 = ( n501 & ~n517 ) | ( n501 & n519 ) | ( ~n517 & n519 ) ;
  assign n521 = n513 | n520 ;
  assign n522 = ( n513 & n517 ) | ( n513 & ~n521 ) | ( n517 & ~n521 ) ;
  assign n523 = ( n507 & ~n510 ) | ( n507 & n522 ) | ( ~n510 & n522 ) ;
  assign n524 = ~n519 & n522 ;
  assign n525 = ( ~n507 & n523 ) | ( ~n507 & n524 ) | ( n523 & n524 ) ;
  assign n526 = ( ~x11 & x172 ) | ( ~x11 & x173 ) | ( x172 & x173 ) ;
  assign n527 = x206 & ~n526 ;
  assign n528 = ( x11 & ~x206 ) | ( x11 & n527 ) | ( ~x206 & n527 ) ;
  assign n529 = x172 & x206 ;
  assign n530 = ~x11 & n529 ;
  assign n531 = x11 | n529 ;
  assign n532 = ( ~n529 & n530 ) | ( ~n529 & n531 ) | ( n530 & n531 ) ;
  assign n533 = x173 & ~x206 ;
  assign n534 = ( x11 & x173 ) | ( x11 & n533 ) | ( x173 & n533 ) ;
  assign n535 = ( x11 & ~x173 ) | ( x11 & n533 ) | ( ~x173 & n533 ) ;
  assign n536 = ( x173 & ~n534 ) | ( x173 & n535 ) | ( ~n534 & n535 ) ;
  assign n537 = ( ~n528 & n532 ) | ( ~n528 & n536 ) | ( n532 & n536 ) ;
  assign n538 = ~n525 & n537 ;
  assign n539 = ( n525 & ~n528 ) | ( n525 & n538 ) | ( ~n528 & n538 ) ;
  assign n540 = ( n461 & n486 ) | ( n461 & n539 ) | ( n486 & n539 ) ;
  assign n541 = ~x168 & n503 ;
  assign n542 = ( ~n503 & n504 ) | ( ~n503 & n541 ) | ( n504 & n541 ) ;
  assign n543 = n496 & n519 ;
  assign n544 = ( ~n501 & n542 ) | ( ~n501 & n543 ) | ( n542 & n543 ) ;
  assign n545 = n501 & n544 ;
  assign n546 = n491 & n545 ;
  assign n547 = ~n532 & n546 ;
  assign n548 = ~n536 & n547 ;
  assign n549 = n539 & ~n548 ;
  assign n550 = ( ~n461 & n540 ) | ( ~n461 & n549 ) | ( n540 & n549 ) ;
  assign n551 = ( n428 & ~n436 ) | ( n428 & n550 ) | ( ~n436 & n550 ) ;
  assign n552 = ~n548 & n550 ;
  assign n553 = ( ~n428 & n551 ) | ( ~n428 & n552 ) | ( n551 & n552 ) ;
  assign n554 = x100 & ~n240 ;
  assign n555 = ( x5 & n240 ) | ( x5 & ~n554 ) | ( n240 & ~n554 ) ;
  assign n556 = x5 & ~x180 ;
  assign n557 = x5 | x27 ;
  assign n558 = ( ~x5 & n556 ) | ( ~x5 & n557 ) | ( n556 & n557 ) ;
  assign n559 = ~n555 & n558 ;
  assign n560 = n555 & n558 ;
  assign n561 = ( n555 & n559 ) | ( n555 & ~n560 ) | ( n559 & ~n560 ) ;
  assign n562 = x5 & x178 ;
  assign n563 = x5 & ~x102 ;
  assign n564 = ~x5 & x71 ;
  assign n565 = ( x5 & ~n563 ) | ( x5 & n564 ) | ( ~n563 & n564 ) ;
  assign n566 = x5 | x43 ;
  assign n567 = ( ~n562 & n565 ) | ( ~n562 & n566 ) | ( n565 & n566 ) ;
  assign n568 = ( n565 & n566 ) | ( n565 & ~n567 ) | ( n566 & ~n567 ) ;
  assign n569 = ( n562 & n567 ) | ( n562 & ~n568 ) | ( n567 & ~n568 ) ;
  assign n570 = x5 & ~x177 ;
  assign n571 = x5 | x42 ;
  assign n572 = ( ~x5 & n570 ) | ( ~x5 & n571 ) | ( n570 & n571 ) ;
  assign n573 = x5 & ~x103 ;
  assign n574 = ( x5 & n235 ) | ( x5 & ~n573 ) | ( n235 & ~n573 ) ;
  assign n575 = ( ~n569 & n572 ) | ( ~n569 & n574 ) | ( n572 & n574 ) ;
  assign n576 = x5 & ~x176 ;
  assign n577 = x5 | x28 ;
  assign n578 = ( ~x5 & n576 ) | ( ~x5 & n577 ) | ( n576 & n577 ) ;
  assign n579 = x5 & ~x94 ;
  assign n580 = ( x5 & n247 ) | ( x5 & ~n579 ) | ( n247 & ~n579 ) ;
  assign n581 = ~n578 & n580 ;
  assign n582 = n578 & n580 ;
  assign n583 = ( n578 & n581 ) | ( n578 & ~n582 ) | ( n581 & ~n582 ) ;
  assign n584 = ( n572 & n574 ) | ( n572 & n583 ) | ( n574 & n583 ) ;
  assign n585 = ~n575 & n584 ;
  assign n586 = x5 & x179 ;
  assign n587 = x5 & ~x101 ;
  assign n588 = ( x5 & n253 ) | ( x5 & ~n587 ) | ( n253 & ~n587 ) ;
  assign n589 = x5 | x44 ;
  assign n590 = ( ~n586 & n588 ) | ( ~n586 & n589 ) | ( n588 & n589 ) ;
  assign n591 = ( n588 & n589 ) | ( n588 & ~n590 ) | ( n589 & ~n590 ) ;
  assign n592 = ( n586 & n590 ) | ( n586 & ~n591 ) | ( n590 & ~n591 ) ;
  assign n593 = x97 & ~n240 ;
  assign n594 = ( x5 & n240 ) | ( x5 & ~n593 ) | ( n240 & ~n593 ) ;
  assign n595 = x5 & ~x183 ;
  assign n596 = x5 | x54 ;
  assign n597 = ( ~x5 & n595 ) | ( ~x5 & n596 ) | ( n595 & n596 ) ;
  assign n598 = ~n594 & n597 ;
  assign n599 = n594 & n597 ;
  assign n600 = ( n594 & n598 ) | ( n594 & ~n599 ) | ( n598 & ~n599 ) ;
  assign n601 = x96 & ~n240 ;
  assign n602 = ( x5 & n240 ) | ( x5 & ~n601 ) | ( n240 & ~n601 ) ;
  assign n603 = x5 & ~x184 ;
  assign n604 = x5 | x55 ;
  assign n605 = ( ~x5 & n603 ) | ( ~x5 & n604 ) | ( n603 & n604 ) ;
  assign n606 = ~n602 & n605 ;
  assign n607 = n602 & n605 ;
  assign n608 = ( n602 & n606 ) | ( n602 & ~n607 ) | ( n606 & ~n607 ) ;
  assign n609 = x5 & ~x181 ;
  assign n610 = x5 | x26 ;
  assign n611 = ( ~x5 & n609 ) | ( ~x5 & n610 ) | ( n609 & n610 ) ;
  assign n612 = x98 & ~n240 ;
  assign n613 = ( x5 & n240 ) | ( x5 & ~n612 ) | ( n240 & ~n612 ) ;
  assign n614 = x5 & ~x182 ;
  assign n615 = x5 | x45 ;
  assign n616 = ( ~x5 & n614 ) | ( ~x5 & n615 ) | ( n614 & n615 ) ;
  assign n617 = ~n613 & n616 ;
  assign n618 = n613 & n616 ;
  assign n619 = ( n613 & n617 ) | ( n613 & ~n618 ) | ( n617 & ~n618 ) ;
  assign n620 = x99 & ~n240 ;
  assign n621 = ( x5 & n240 ) | ( x5 & ~n620 ) | ( n240 & ~n620 ) ;
  assign n622 = ( ~n611 & n619 ) | ( ~n611 & n621 ) | ( n619 & n621 ) ;
  assign n623 = n621 & ~n622 ;
  assign n624 = ( n611 & n622 ) | ( n611 & ~n623 ) | ( n622 & ~n623 ) ;
  assign n625 = n608 | n624 ;
  assign n626 = n600 | n625 ;
  assign n627 = n592 & ~n626 ;
  assign n628 = ( n561 & n585 ) | ( n561 & n627 ) | ( n585 & n627 ) ;
  assign n629 = ~n561 & n628 ;
  assign n630 = x5 & ~x190 ;
  assign n631 = x5 | x32 ;
  assign n632 = ( ~x5 & n630 ) | ( ~x5 & n631 ) | ( n630 & n631 ) ;
  assign n633 = x5 & ~x127 ;
  assign n634 = ( x5 & n292 ) | ( x5 & ~n633 ) | ( n292 & ~n633 ) ;
  assign n635 = ~n632 & n634 ;
  assign n636 = n632 & n634 ;
  assign n637 = ( n632 & n635 ) | ( n632 & ~n636 ) | ( n635 & ~n636 ) ;
  assign n638 = x5 & ~x187 ;
  assign n639 = x5 | x33 ;
  assign n640 = ( ~x5 & n638 ) | ( ~x5 & n639 ) | ( n638 & n639 ) ;
  assign n641 = x5 & ~x188 ;
  assign n642 = x5 | x35 ;
  assign n643 = ( ~x5 & n641 ) | ( ~x5 & n642 ) | ( n641 & n642 ) ;
  assign n644 = x5 & ~x129 ;
  assign n645 = ( x5 & n304 ) | ( x5 & ~n644 ) | ( n304 & ~n644 ) ;
  assign n646 = ~n643 & n645 ;
  assign n647 = n643 & n645 ;
  assign n648 = ( n643 & n646 ) | ( n643 & ~n647 ) | ( n646 & ~n647 ) ;
  assign n649 = x5 & ~x130 ;
  assign n650 = ( x5 & n298 ) | ( x5 & ~n649 ) | ( n298 & ~n649 ) ;
  assign n651 = n648 & n650 ;
  assign n652 = ( ~n637 & n640 ) | ( ~n637 & n651 ) | ( n640 & n651 ) ;
  assign n653 = n637 & n652 ;
  assign n654 = ~n640 & n650 ;
  assign n655 = n640 & n650 ;
  assign n656 = ( n640 & n654 ) | ( n640 & ~n655 ) | ( n654 & ~n655 ) ;
  assign n657 = x5 & ~x121 ;
  assign n658 = ( x5 & n226 ) | ( x5 & ~n657 ) | ( n226 & ~n657 ) ;
  assign n659 = x31 & n658 ;
  assign n660 = ~x5 & n659 ;
  assign n661 = n648 & n660 ;
  assign n662 = ( ~n637 & n656 ) | ( ~n637 & n661 ) | ( n656 & n661 ) ;
  assign n663 = n637 & n662 ;
  assign n664 = x5 & ~x189 ;
  assign n665 = x5 | x34 ;
  assign n666 = ( ~x5 & n664 ) | ( ~x5 & n665 ) | ( n664 & n665 ) ;
  assign n667 = x5 & ~x128 ;
  assign n668 = ( x5 & n318 ) | ( x5 & ~n667 ) | ( n318 & ~n667 ) ;
  assign n669 = ~n666 & n668 ;
  assign n670 = n666 & n668 ;
  assign n671 = ( n666 & n669 ) | ( n666 & ~n670 ) | ( n669 & ~n670 ) ;
  assign n672 = n637 & n645 ;
  assign n673 = ( n643 & ~n671 ) | ( n643 & n672 ) | ( ~n671 & n672 ) ;
  assign n674 = n671 & n673 ;
  assign n675 = ( n632 & n634 ) | ( n632 & n670 ) | ( n634 & n670 ) ;
  assign n676 = n674 | n675 ;
  assign n677 = ( ~n653 & n663 ) | ( ~n653 & n676 ) | ( n663 & n676 ) ;
  assign n678 = n671 | n676 ;
  assign n679 = ( n653 & n677 ) | ( n653 & n678 ) | ( n677 & n678 ) ;
  assign n680 = x5 & ~x193 ;
  assign n681 = x5 | x18 ;
  assign n682 = ( ~x5 & n680 ) | ( ~x5 & n681 ) | ( n680 & n681 ) ;
  assign n683 = x5 & ~x124 ;
  assign n684 = ( x5 & n343 ) | ( x5 & ~n683 ) | ( n343 & ~n683 ) ;
  assign n685 = ~n682 & n684 ;
  assign n686 = n682 & n684 ;
  assign n687 = ( n682 & n685 ) | ( n682 & ~n686 ) | ( n685 & ~n686 ) ;
  assign n688 = x5 & ~x194 ;
  assign n689 = x5 | x19 ;
  assign n690 = ( ~x5 & n688 ) | ( ~x5 & n689 ) | ( n688 & n689 ) ;
  assign n691 = x5 & ~x123 ;
  assign n692 = ( x5 & n331 ) | ( x5 & ~n691 ) | ( n331 & ~n691 ) ;
  assign n693 = ~n690 & n692 ;
  assign n694 = n690 & n692 ;
  assign n695 = ( n690 & n693 ) | ( n690 & ~n694 ) | ( n693 & ~n694 ) ;
  assign n696 = x5 & ~x126 ;
  assign n697 = ( x5 & n349 ) | ( x5 & ~n696 ) | ( n349 & ~n696 ) ;
  assign n698 = x5 & ~x192 ;
  assign n699 = x5 | x17 ;
  assign n700 = ( ~x5 & n698 ) | ( ~x5 & n699 ) | ( n698 & n699 ) ;
  assign n701 = x5 & ~x125 ;
  assign n702 = ( x5 & n337 ) | ( x5 & ~n701 ) | ( n337 & ~n701 ) ;
  assign n703 = ~n700 & n702 ;
  assign n704 = n700 & n702 ;
  assign n705 = ( n700 & n703 ) | ( n700 & ~n704 ) | ( n703 & ~n704 ) ;
  assign n706 = x5 & ~x191 ;
  assign n707 = x5 | x16 ;
  assign n708 = ( ~x5 & n706 ) | ( ~x5 & n707 ) | ( n706 & n707 ) ;
  assign n709 = ( n697 & n705 ) | ( n697 & n708 ) | ( n705 & n708 ) ;
  assign n710 = ~n708 & n709 ;
  assign n711 = ( ~n697 & n709 ) | ( ~n697 & n710 ) | ( n709 & n710 ) ;
  assign n712 = n695 & n711 ;
  assign n713 = n687 & n712 ;
  assign n714 = x5 & ~x203 ;
  assign n715 = x5 | x24 ;
  assign n716 = ( ~x5 & n714 ) | ( ~x5 & n715 ) | ( n714 & n715 ) ;
  assign n717 = x5 & ~x113 ;
  assign n718 = ( x5 & n397 ) | ( x5 & ~n717 ) | ( n397 & ~n717 ) ;
  assign n719 = ~n716 & n718 ;
  assign n720 = n716 & n718 ;
  assign n721 = ( n716 & n719 ) | ( n716 & ~n720 ) | ( n719 & ~n720 ) ;
  assign n722 = x5 & ~x204 ;
  assign n723 = x5 | x25 ;
  assign n724 = ( ~x5 & n722 ) | ( ~x5 & n723 ) | ( n722 & n723 ) ;
  assign n725 = x5 & ~x112 ;
  assign n726 = ( x5 & n391 ) | ( x5 & ~n725 ) | ( n391 & ~n725 ) ;
  assign n727 = ~n724 & n726 ;
  assign n728 = n724 & n726 ;
  assign n729 = ( n724 & n727 ) | ( n724 & ~n728 ) | ( n727 & ~n728 ) ;
  assign n730 = x5 & ~x115 ;
  assign n731 = ( x5 & n409 ) | ( x5 & ~n730 ) | ( n409 & ~n730 ) ;
  assign n732 = x5 & ~x202 ;
  assign n733 = x5 | x23 ;
  assign n734 = ( ~x5 & n732 ) | ( ~x5 & n733 ) | ( n732 & n733 ) ;
  assign n735 = x5 & ~x114 ;
  assign n736 = ( x5 & n403 ) | ( x5 & ~n735 ) | ( n403 & ~n735 ) ;
  assign n737 = ~n734 & n736 ;
  assign n738 = n734 & n736 ;
  assign n739 = ( n734 & n737 ) | ( n734 & ~n738 ) | ( n737 & ~n738 ) ;
  assign n740 = x5 & ~x201 ;
  assign n741 = x5 | x38 ;
  assign n742 = ( ~x5 & n740 ) | ( ~x5 & n741 ) | ( n740 & n741 ) ;
  assign n743 = ( n731 & n739 ) | ( n731 & n742 ) | ( n739 & n742 ) ;
  assign n744 = ~n742 & n743 ;
  assign n745 = ( ~n731 & n743 ) | ( ~n731 & n744 ) | ( n743 & n744 ) ;
  assign n746 = n729 & n745 ;
  assign n747 = n721 & n746 ;
  assign n748 = x5 & ~x200 ;
  assign n749 = x5 | x39 ;
  assign n750 = ( ~x5 & n748 ) | ( ~x5 & n749 ) | ( n748 & n749 ) ;
  assign n751 = x5 & ~x116 ;
  assign n752 = ( x5 & n364 ) | ( x5 & ~n751 ) | ( n364 & ~n751 ) ;
  assign n753 = ~n750 & n752 ;
  assign n754 = n750 & n752 ;
  assign n755 = ( n750 & n753 ) | ( n750 & ~n754 ) | ( n753 & ~n754 ) ;
  assign n756 = x5 & x198 ;
  assign n757 = x5 & ~x118 ;
  assign n758 = ~x5 & x49 ;
  assign n759 = ( x5 & ~n757 ) | ( x5 & n758 ) | ( ~n757 & n758 ) ;
  assign n760 = x5 | x22 ;
  assign n761 = ( ~n756 & n759 ) | ( ~n756 & n760 ) | ( n759 & n760 ) ;
  assign n762 = ( n759 & n760 ) | ( n759 & ~n761 ) | ( n760 & ~n761 ) ;
  assign n763 = ( n756 & n761 ) | ( n756 & ~n762 ) | ( n761 & ~n762 ) ;
  assign n764 = x5 & x199 ;
  assign n765 = x5 & ~x117 ;
  assign n766 = ( x5 & n376 ) | ( x5 & ~n765 ) | ( n376 & ~n765 ) ;
  assign n767 = x5 | x40 ;
  assign n768 = ( ~n764 & n766 ) | ( ~n764 & n767 ) | ( n766 & n767 ) ;
  assign n769 = ( n766 & n767 ) | ( n766 & ~n768 ) | ( n767 & ~n768 ) ;
  assign n770 = ( n764 & n768 ) | ( n764 & ~n769 ) | ( n768 & ~n769 ) ;
  assign n771 = x5 & ~x197 ;
  assign n772 = x5 | x37 ;
  assign n773 = ( ~x5 & n771 ) | ( ~x5 & n772 ) | ( n771 & n772 ) ;
  assign n774 = x5 & ~x119 ;
  assign n775 = ( x5 & n358 ) | ( x5 & ~n774 ) | ( n358 & ~n774 ) ;
  assign n776 = x5 & ~x196 ;
  assign n777 = x5 | x36 ;
  assign n778 = ( ~x5 & n776 ) | ( ~x5 & n777 ) | ( n776 & n777 ) ;
  assign n779 = x5 & ~x110 ;
  assign n780 = ( x5 & n370 ) | ( x5 & ~n779 ) | ( n370 & ~n779 ) ;
  assign n781 = n778 | n780 ;
  assign n782 = ( n773 & n775 ) | ( n773 & n781 ) | ( n775 & n781 ) ;
  assign n783 = n778 & n780 ;
  assign n784 = ( n773 & n775 ) | ( n773 & n783 ) | ( n775 & n783 ) ;
  assign n785 = n782 & ~n784 ;
  assign n786 = n770 & n785 ;
  assign n787 = ( ~n755 & n763 ) | ( ~n755 & n786 ) | ( n763 & n786 ) ;
  assign n788 = n755 & n787 ;
  assign n789 = n747 & n788 ;
  assign n790 = ( ~n679 & n713 ) | ( ~n679 & n789 ) | ( n713 & n789 ) ;
  assign n791 = n697 & n705 ;
  assign n792 = ( ~n695 & n708 ) | ( ~n695 & n791 ) | ( n708 & n791 ) ;
  assign n793 = n695 & n792 ;
  assign n794 = ~n687 & n793 ;
  assign n795 = n687 & n702 ;
  assign n796 = ( ~n695 & n700 ) | ( ~n695 & n795 ) | ( n700 & n795 ) ;
  assign n797 = n695 & n796 ;
  assign n798 = ( n686 & n690 ) | ( n686 & n692 ) | ( n690 & n692 ) ;
  assign n799 = n797 | n798 ;
  assign n800 = ( n793 & ~n794 ) | ( n793 & n799 ) | ( ~n794 & n799 ) ;
  assign n801 = n789 & n800 ;
  assign n802 = ( n679 & n790 ) | ( n679 & n801 ) | ( n790 & n801 ) ;
  assign n803 = n629 & n802 ;
  assign n804 = ~x31 & n658 ;
  assign n805 = ( x5 & x31 ) | ( x5 & ~n658 ) | ( x31 & ~n658 ) ;
  assign n806 = ( n656 & n804 ) | ( n656 & n805 ) | ( n804 & n805 ) ;
  assign n807 = n637 & n806 ;
  assign n808 = ( n648 & ~n671 ) | ( n648 & n807 ) | ( ~n671 & n807 ) ;
  assign n809 = n671 & n808 ;
  assign n810 = x48 & n713 ;
  assign n811 = ( ~n789 & n809 ) | ( ~n789 & n810 ) | ( n809 & n810 ) ;
  assign n812 = n789 & n811 ;
  assign n813 = n629 & n812 ;
  assign n814 = n763 & n775 ;
  assign n815 = ( ~n755 & n773 ) | ( ~n755 & n814 ) | ( n773 & n814 ) ;
  assign n816 = n755 & n815 ;
  assign n817 = ( ~n755 & n773 ) | ( ~n755 & n775 ) | ( n773 & n775 ) ;
  assign n818 = ( n763 & n773 ) | ( n763 & n775 ) | ( n773 & n775 ) ;
  assign n819 = ~n817 & n818 ;
  assign n820 = n778 & n819 ;
  assign n821 = n780 & n820 ;
  assign n822 = ( x5 & x22 ) | ( x5 & n759 ) | ( x22 & n759 ) ;
  assign n823 = ( x5 & x198 ) | ( x5 & ~n759 ) | ( x198 & ~n759 ) ;
  assign n824 = n822 & ~n823 ;
  assign n825 = n755 & n824 ;
  assign n826 = n770 & n825 ;
  assign n827 = ( x5 & x40 ) | ( x5 & n766 ) | ( x40 & n766 ) ;
  assign n828 = ( x5 & x199 ) | ( x5 & ~n766 ) | ( x199 & ~n766 ) ;
  assign n829 = n827 & ~n828 ;
  assign n830 = ( n750 & n752 ) | ( n750 & n829 ) | ( n752 & n829 ) ;
  assign n831 = n826 | n830 ;
  assign n832 = ( ~n816 & n821 ) | ( ~n816 & n831 ) | ( n821 & n831 ) ;
  assign n833 = n770 | n831 ;
  assign n834 = ( n816 & n832 ) | ( n816 & n833 ) | ( n832 & n833 ) ;
  assign n835 = ( n629 & n747 ) | ( n629 & ~n834 ) | ( n747 & ~n834 ) ;
  assign n836 = n731 & n739 ;
  assign n837 = ( ~n729 & n742 ) | ( ~n729 & n836 ) | ( n742 & n836 ) ;
  assign n838 = n729 & n837 ;
  assign n839 = ~n721 & n838 ;
  assign n840 = n721 & n736 ;
  assign n841 = ( ~n729 & n734 ) | ( ~n729 & n840 ) | ( n734 & n840 ) ;
  assign n842 = n729 & n841 ;
  assign n843 = ( n720 & n724 ) | ( n720 & n726 ) | ( n724 & n726 ) ;
  assign n844 = n842 | n843 ;
  assign n845 = ( n838 & ~n839 ) | ( n838 & n844 ) | ( ~n839 & n844 ) ;
  assign n846 = n629 & n845 ;
  assign n847 = ( n834 & n835 ) | ( n834 & n846 ) | ( n835 & n846 ) ;
  assign n848 = n569 & n574 ;
  assign n849 = ( n561 & n572 ) | ( n561 & n848 ) | ( n572 & n848 ) ;
  assign n850 = ~n561 & n849 ;
  assign n851 = ( n561 & n572 ) | ( n561 & n574 ) | ( n572 & n574 ) ;
  assign n852 = ( n569 & n572 ) | ( n569 & n574 ) | ( n572 & n574 ) ;
  assign n853 = ~n851 & n852 ;
  assign n854 = n578 & n853 ;
  assign n855 = n580 & n854 ;
  assign n856 = ( x5 & x43 ) | ( x5 & n565 ) | ( x43 & n565 ) ;
  assign n857 = ( x5 & x178 ) | ( x5 & ~n565 ) | ( x178 & ~n565 ) ;
  assign n858 = n856 & ~n857 ;
  assign n859 = ( x5 & x44 ) | ( x5 & n588 ) | ( x44 & n588 ) ;
  assign n860 = ( x5 & x179 ) | ( x5 & ~n588 ) | ( x179 & ~n588 ) ;
  assign n861 = n859 & ~n860 ;
  assign n862 = ( ~n555 & n558 ) | ( ~n555 & n861 ) | ( n558 & n861 ) ;
  assign n863 = ( ~n561 & n592 ) | ( ~n561 & n862 ) | ( n592 & n862 ) ;
  assign n864 = n858 & ~n863 ;
  assign n865 = ( n858 & n862 ) | ( n858 & ~n864 ) | ( n862 & ~n864 ) ;
  assign n866 = ( ~n850 & n855 ) | ( ~n850 & n865 ) | ( n855 & n865 ) ;
  assign n867 = n592 | n865 ;
  assign n868 = ( n850 & n866 ) | ( n850 & n867 ) | ( n866 & n867 ) ;
  assign n869 = n626 & n868 ;
  assign n870 = ( ~n600 & n608 ) | ( ~n600 & n617 ) | ( n608 & n617 ) ;
  assign n871 = n619 | n621 ;
  assign n872 = ( n608 & n611 ) | ( n608 & ~n871 ) | ( n611 & ~n871 ) ;
  assign n873 = ~n608 & n872 ;
  assign n874 = ~n600 & n873 ;
  assign n875 = ( ~n608 & n870 ) | ( ~n608 & n874 ) | ( n870 & n874 ) ;
  assign n876 = ( n598 & ~n602 ) | ( n598 & n605 ) | ( ~n602 & n605 ) ;
  assign n877 = n875 | n876 ;
  assign n878 = ( n868 & ~n869 ) | ( n868 & n877 ) | ( ~n869 & n877 ) ;
  assign n879 = ~x166 & x206 ;
  assign n880 = ~x174 & x206 ;
  assign n881 = x89 & ~n240 ;
  assign n882 = ( x5 & n240 ) | ( x5 & ~n881 ) | ( n240 & ~n881 ) ;
  assign n883 = x5 & ~x171 ;
  assign n884 = x5 | x47 ;
  assign n885 = ( ~x5 & n883 ) | ( ~x5 & n884 ) | ( n883 & n884 ) ;
  assign n886 = ~n882 & n885 ;
  assign n887 = n882 & n885 ;
  assign n888 = ( n882 & n886 ) | ( n882 & ~n887 ) | ( n886 & ~n887 ) ;
  assign n889 = x5 & ~x169 ;
  assign n890 = x5 | x56 ;
  assign n891 = ( ~x5 & n889 ) | ( ~x5 & n890 ) | ( n889 & n890 ) ;
  assign n892 = x5 & x53 ;
  assign n893 = x91 & ~n240 ;
  assign n894 = ( x5 & n240 ) | ( x5 & ~n893 ) | ( n240 & ~n893 ) ;
  assign n895 = x5 | x46 ;
  assign n896 = ( ~n892 & n894 ) | ( ~n892 & n895 ) | ( n894 & n895 ) ;
  assign n897 = ( n894 & n895 ) | ( n894 & ~n896 ) | ( n895 & ~n896 ) ;
  assign n898 = ( n892 & n896 ) | ( n892 & ~n897 ) | ( n896 & ~n897 ) ;
  assign n899 = x92 & ~n240 ;
  assign n900 = ( x5 & n240 ) | ( x5 & ~n899 ) | ( n240 & ~n899 ) ;
  assign n901 = n898 | n900 ;
  assign n902 = ( n888 & n891 ) | ( n888 & ~n901 ) | ( n891 & ~n901 ) ;
  assign n903 = ~n888 & n902 ;
  assign n904 = x5 & ~x168 ;
  assign n905 = x5 | x58 ;
  assign n906 = ( ~x5 & n904 ) | ( ~x5 & n905 ) | ( n904 & n905 ) ;
  assign n907 = ( n888 & n891 ) | ( n888 & ~n900 ) | ( n891 & ~n900 ) ;
  assign n908 = ( ~n891 & n898 ) | ( ~n891 & n900 ) | ( n898 & n900 ) ;
  assign n909 = n907 | n908 ;
  assign n910 = n240 | n909 ;
  assign n911 = n906 & ~n910 ;
  assign n912 = ( x5 & x53 ) | ( x5 & n894 ) | ( x53 & n894 ) ;
  assign n913 = ( x5 & x46 ) | ( x5 & ~n894 ) | ( x46 & ~n894 ) ;
  assign n914 = ~n912 & n913 ;
  assign n915 = x90 & ~n240 ;
  assign n916 = ( x5 & n240 ) | ( x5 & ~n915 ) | ( n240 & ~n915 ) ;
  assign n917 = x5 & ~x170 ;
  assign n918 = x5 | x57 ;
  assign n919 = ( ~x5 & n917 ) | ( ~x5 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ~n916 & n919 ;
  assign n921 = ( ~n882 & n885 ) | ( ~n882 & n920 ) | ( n885 & n920 ) ;
  assign n922 = n916 & n919 ;
  assign n923 = ( n916 & n920 ) | ( n916 & ~n922 ) | ( n920 & ~n922 ) ;
  assign n924 = ( n888 & ~n921 ) | ( n888 & n923 ) | ( ~n921 & n923 ) ;
  assign n925 = n914 & n924 ;
  assign n926 = ( n914 & n921 ) | ( n914 & ~n925 ) | ( n921 & ~n925 ) ;
  assign n927 = ( ~n903 & n911 ) | ( ~n903 & n926 ) | ( n911 & n926 ) ;
  assign n928 = n923 & ~n926 ;
  assign n929 = ( n903 & n927 ) | ( n903 & ~n928 ) | ( n927 & ~n928 ) ;
  assign n930 = ( n879 & n880 ) | ( n879 & ~n929 ) | ( n880 & ~n929 ) ;
  assign n931 = ( ~n880 & n929 ) | ( ~n880 & n930 ) | ( n929 & n930 ) ;
  assign n932 = ( x11 & ~n879 ) | ( x11 & n931 ) | ( ~n879 & n931 ) ;
  assign n933 = ( ~n847 & n878 ) | ( ~n847 & n932 ) | ( n878 & n932 ) ;
  assign n934 = n240 & ~n906 ;
  assign n935 = ( ~n891 & n900 ) | ( ~n891 & n934 ) | ( n900 & n934 ) ;
  assign n936 = ~n240 & n906 ;
  assign n937 = ( n891 & ~n900 ) | ( n891 & n936 ) | ( ~n900 & n936 ) ;
  assign n938 = n935 | n937 ;
  assign n939 = n923 | n938 ;
  assign n940 = ( ~n888 & n898 ) | ( ~n888 & n939 ) | ( n898 & n939 ) ;
  assign n941 = n888 | n940 ;
  assign n942 = ( x11 & ~n880 ) | ( x11 & n941 ) | ( ~n880 & n941 ) ;
  assign n943 = ( ~n879 & n880 ) | ( ~n879 & n942 ) | ( n880 & n942 ) ;
  assign n944 = ( ~x11 & n879 ) | ( ~x11 & n942 ) | ( n879 & n942 ) ;
  assign n945 = n943 | n944 ;
  assign n946 = ~n932 & n945 ;
  assign n947 = ( n847 & n933 ) | ( n847 & ~n946 ) | ( n933 & ~n946 ) ;
  assign n948 = ( ~n803 & n813 ) | ( ~n803 & n947 ) | ( n813 & n947 ) ;
  assign n949 = n945 & ~n947 ;
  assign n950 = ( n803 & n948 ) | ( n803 & ~n949 ) | ( n948 & ~n949 ) ;
  assign n951 = ( ~n362 & n374 ) | ( ~n362 & n386 ) | ( n374 & n386 ) ;
  assign n952 = n362 | n951 ;
  assign n953 = n368 | n952 ;
  assign n954 = n416 | n953 ;
  assign n955 = ( n329 & n356 ) | ( n329 & n954 ) | ( n356 & n954 ) ;
  assign n956 = n425 & ~n954 ;
  assign n957 = ( n329 & ~n955 ) | ( n329 & n956 ) | ( ~n955 & n956 ) ;
  assign n958 = ( ~n239 & n251 ) | ( ~n239 & n263 ) | ( n251 & n263 ) ;
  assign n959 = n239 | n958 ;
  assign n960 = n245 & ~n959 ;
  assign n961 = n289 & n960 ;
  assign n962 = n957 & n961 ;
  assign n963 = n302 | n323 ;
  assign n964 = ( ~n230 & n308 ) | ( ~n230 & n963 ) | ( n308 & n963 ) ;
  assign n965 = n230 | n964 ;
  assign n966 = n296 | n965 ;
  assign n967 = x205 & ~n966 ;
  assign n968 = ( ~n356 & n954 ) | ( ~n356 & n967 ) | ( n954 & n967 ) ;
  assign n969 = ~n954 & n968 ;
  assign n970 = n961 & n969 ;
  assign n971 = n460 & n961 ;
  assign n972 = ( n486 & n539 ) | ( n486 & n971 ) | ( n539 & n971 ) ;
  assign n973 = ( ~n491 & n542 ) | ( ~n491 & n543 ) | ( n542 & n543 ) ;
  assign n974 = n491 & n973 ;
  assign n975 = n501 & n974 ;
  assign n976 = ~n532 & n975 ;
  assign n977 = ~n536 & n976 ;
  assign n978 = n539 & ~n977 ;
  assign n979 = ( ~n971 & n972 ) | ( ~n971 & n978 ) | ( n972 & n978 ) ;
  assign n980 = ( n962 & ~n970 ) | ( n962 & n979 ) | ( ~n970 & n979 ) ;
  assign n981 = ~n977 & n979 ;
  assign n982 = ( ~n962 & n980 ) | ( ~n962 & n981 ) | ( n980 & n981 ) ;
  assign n983 = ~n302 & n311 ;
  assign n984 = x205 & ~n308 ;
  assign n985 = ( n230 & ~n302 ) | ( n230 & n984 ) | ( ~n302 & n984 ) ;
  assign n986 = ~n230 & n985 ;
  assign n987 = n299 & ~n314 ;
  assign n988 = n307 | n987 ;
  assign n989 = ( ~x189 & n319 ) | ( ~x189 & n988 ) | ( n319 & n988 ) ;
  assign n990 = ( ~n983 & n986 ) | ( ~n983 & n989 ) | ( n986 & n989 ) ;
  assign n991 = n323 & ~n989 ;
  assign n992 = ( n983 & n990 ) | ( n983 & ~n991 ) | ( n990 & ~n991 ) ;
  assign n993 = n296 | n992 ;
  assign n994 = ~n296 & n992 ;
  assign n995 = ( ~n992 & n993 ) | ( ~n992 & n994 ) | ( n993 & n994 ) ;
  assign n996 = n983 | n986 ;
  assign n997 = n988 | n996 ;
  assign n998 = n323 & n997 ;
  assign n999 = n323 | n997 ;
  assign n1000 = ~n998 & n999 ;
  assign n1001 = ( ~x187 & n299 ) | ( ~x187 & n310 ) | ( n299 & n310 ) ;
  assign n1002 = ( n230 & n302 ) | ( n230 & ~n1001 ) | ( n302 & ~n1001 ) ;
  assign n1003 = x205 & n1002 ;
  assign n1004 = ( x205 & n1001 ) | ( x205 & ~n1003 ) | ( n1001 & ~n1003 ) ;
  assign n1005 = n308 | n1004 ;
  assign n1006 = ~n308 & n1004 ;
  assign n1007 = ( ~n1004 & n1005 ) | ( ~n1004 & n1006 ) | ( n1005 & n1006 ) ;
  assign n1008 = n230 & ~n310 ;
  assign n1009 = ( x205 & n310 ) | ( x205 & ~n1008 ) | ( n310 & ~n1008 ) ;
  assign n1010 = ~n302 & n1009 ;
  assign n1011 = n302 | n1009 ;
  assign n1012 = ( ~n1009 & n1010 ) | ( ~n1009 & n1011 ) | ( n1010 & n1011 ) ;
  assign n1013 = ~n341 & n352 ;
  assign n1014 = ( ~n340 & n346 ) | ( ~n340 & n1013 ) | ( n346 & n1013 ) ;
  assign n1015 = ~n346 & n347 ;
  assign n1016 = ( n340 & n1014 ) | ( n340 & ~n1015 ) | ( n1014 & ~n1015 ) ;
  assign n1017 = x205 | n329 ;
  assign n1018 = ( n329 & ~n432 ) | ( n329 & n1017 ) | ( ~n432 & n1017 ) ;
  assign n1019 = n1016 & ~n1018 ;
  assign n1020 = n341 | n347 ;
  assign n1021 = ( ~n350 & n351 ) | ( ~n350 & n1020 ) | ( n351 & n1020 ) ;
  assign n1022 = ( ~x193 & n340 ) | ( ~x193 & n344 ) | ( n340 & n344 ) ;
  assign n1023 = n1021 & ~n1022 ;
  assign n1024 = n1018 & ~n1023 ;
  assign n1025 = ( n335 & n1019 ) | ( n335 & n1024 ) | ( n1019 & n1024 ) ;
  assign n1026 = ( n335 & n1024 ) | ( n335 & ~n1025 ) | ( n1024 & ~n1025 ) ;
  assign n1027 = ( n1019 & ~n1025 ) | ( n1019 & n1026 ) | ( ~n1025 & n1026 ) ;
  assign n1028 = n340 | n1013 ;
  assign n1029 = ~n1018 & n1028 ;
  assign n1030 = n353 & ~n1028 ;
  assign n1031 = ( n341 & ~n1028 ) | ( n341 & n1030 ) | ( ~n1028 & n1030 ) ;
  assign n1032 = n1018 & ~n1031 ;
  assign n1033 = ( n347 & n1029 ) | ( n347 & n1032 ) | ( n1029 & n1032 ) ;
  assign n1034 = ( n347 & n1032 ) | ( n347 & ~n1033 ) | ( n1032 & ~n1033 ) ;
  assign n1035 = ( n1029 & ~n1033 ) | ( n1029 & n1034 ) | ( ~n1033 & n1034 ) ;
  assign n1036 = ( ~x191 & n350 ) | ( ~x191 & n1018 ) | ( n350 & n1018 ) ;
  assign n1037 = n341 & n1036 ;
  assign n1038 = n341 | n1036 ;
  assign n1039 = ~n1037 & n1038 ;
  assign n1040 = n353 | n1018 ;
  assign n1041 = ~n353 & n1018 ;
  assign n1042 = ( ~n1018 & n1040 ) | ( ~n1018 & n1041 ) | ( n1040 & n1041 ) ;
  assign n1043 = x5 & ~x150 ;
  assign n1044 = x5 | x60 ;
  assign n1045 = ( n371 & ~n1043 ) | ( n371 & n1044 ) | ( ~n1043 & n1044 ) ;
  assign n1046 = ( n371 & n1044 ) | ( n371 & ~n1045 ) | ( n1044 & ~n1045 ) ;
  assign n1047 = ( n1043 & n1045 ) | ( n1043 & ~n1046 ) | ( n1045 & ~n1046 ) ;
  assign n1048 = ( n359 & ~n381 ) | ( n359 & n382 ) | ( ~n381 & n382 ) ;
  assign n1049 = ( n359 & n382 ) | ( n359 & ~n1048 ) | ( n382 & ~n1048 ) ;
  assign n1050 = ( n381 & n1048 ) | ( n381 & ~n1049 ) | ( n1048 & ~n1049 ) ;
  assign n1051 = ( n365 & n1047 ) | ( n365 & n1050 ) | ( n1047 & n1050 ) ;
  assign n1052 = ( n1047 & n1050 ) | ( n1047 & ~n1051 ) | ( n1050 & ~n1051 ) ;
  assign n1053 = ( n365 & ~n1051 ) | ( n365 & n1052 ) | ( ~n1051 & n1052 ) ;
  assign n1054 = n377 & ~n1053 ;
  assign n1055 = ~n377 & n1053 ;
  assign n1056 = n1054 | n1055 ;
  assign n1057 = ( n392 & n398 ) | ( n392 & n404 ) | ( n398 & n404 ) ;
  assign n1058 = ( n392 & n404 ) | ( n392 & ~n1057 ) | ( n404 & ~n1057 ) ;
  assign n1059 = ( n398 & ~n1057 ) | ( n398 & n1058 ) | ( ~n1057 & n1058 ) ;
  assign n1060 = n410 & ~n1059 ;
  assign n1061 = ~n410 & n1059 ;
  assign n1062 = n1060 | n1061 ;
  assign n1063 = ~n1056 & n1062 ;
  assign n1064 = n1056 & n1062 ;
  assign n1065 = ( n1056 & n1063 ) | ( n1056 & ~n1064 ) | ( n1063 & ~n1064 ) ;
  assign n1066 = ( n236 & ~n258 ) | ( n236 & n259 ) | ( ~n258 & n259 ) ;
  assign n1067 = ( n236 & n259 ) | ( n236 & ~n1066 ) | ( n259 & ~n1066 ) ;
  assign n1068 = ( n258 & n1066 ) | ( n258 & ~n1067 ) | ( n1066 & ~n1067 ) ;
  assign n1069 = x5 & ~x84 ;
  assign n1070 = x5 | x70 ;
  assign n1071 = ( n248 & ~n1069 ) | ( n248 & n1070 ) | ( ~n1069 & n1070 ) ;
  assign n1072 = ( n248 & n1070 ) | ( n248 & ~n1071 ) | ( n1070 & ~n1071 ) ;
  assign n1073 = ( n1069 & n1071 ) | ( n1069 & ~n1072 ) | ( n1071 & ~n1072 ) ;
  assign n1074 = ( n268 & n273 ) | ( n268 & n278 ) | ( n273 & n278 ) ;
  assign n1075 = ( n268 & n278 ) | ( n268 & ~n1074 ) | ( n278 & ~n1074 ) ;
  assign n1076 = ( n273 & ~n1074 ) | ( n273 & n1075 ) | ( ~n1074 & n1075 ) ;
  assign n1077 = n283 & ~n1076 ;
  assign n1078 = ~n283 & n1076 ;
  assign n1079 = n1077 | n1078 ;
  assign n1080 = ~n242 & n254 ;
  assign n1081 = n242 & n254 ;
  assign n1082 = ( n242 & n1080 ) | ( n242 & ~n1081 ) | ( n1080 & ~n1081 ) ;
  assign n1083 = ( n1073 & n1079 ) | ( n1073 & ~n1082 ) | ( n1079 & ~n1082 ) ;
  assign n1084 = ( ~n1079 & n1082 ) | ( ~n1079 & n1083 ) | ( n1082 & n1083 ) ;
  assign n1085 = ( ~n1073 & n1083 ) | ( ~n1073 & n1084 ) | ( n1083 & n1084 ) ;
  assign n1086 = n1068 & n1085 ;
  assign n1087 = n1068 | n1085 ;
  assign n1088 = ~n1086 & n1087 ;
  assign n1089 = ( ~x5 & x138 ) | ( ~x5 & x139 ) | ( x138 & x139 ) ;
  assign n1090 = ( x138 & x139 ) | ( x138 & ~n240 ) | ( x139 & ~n240 ) ;
  assign n1091 = ~n1089 & n1090 ;
  assign n1092 = ( ~x5 & x134 ) | ( ~x5 & x135 ) | ( x134 & x135 ) ;
  assign n1093 = ( x134 & x135 ) | ( x134 & ~n240 ) | ( x135 & ~n240 ) ;
  assign n1094 = ~n1092 & n1093 ;
  assign n1095 = ~n498 & n515 ;
  assign n1096 = n498 & n515 ;
  assign n1097 = ( n498 & n1095 ) | ( n498 & ~n1096 ) | ( n1095 & ~n1096 ) ;
  assign n1098 = n240 | n503 ;
  assign n1099 = ~n240 & n503 ;
  assign n1100 = ( ~n503 & n1098 ) | ( ~n503 & n1099 ) | ( n1098 & n1099 ) ;
  assign n1101 = ( n1094 & n1097 ) | ( n1094 & ~n1100 ) | ( n1097 & ~n1100 ) ;
  assign n1102 = ( ~n1097 & n1100 ) | ( ~n1097 & n1101 ) | ( n1100 & n1101 ) ;
  assign n1103 = ( ~n1094 & n1101 ) | ( ~n1094 & n1102 ) | ( n1101 & n1102 ) ;
  assign n1104 = n1091 & n1103 ;
  assign n1105 = n1091 | n1103 ;
  assign n1106 = ~n1104 & n1105 ;
  assign n1107 = ~n299 & n305 ;
  assign n1108 = n299 & n305 ;
  assign n1109 = ( n299 & n1107 ) | ( n299 & ~n1108 ) | ( n1107 & ~n1108 ) ;
  assign n1110 = x5 & ~x162 ;
  assign n1111 = x5 | x13 ;
  assign n1112 = ( n227 & ~n1110 ) | ( n227 & n1111 ) | ( ~n1110 & n1111 ) ;
  assign n1113 = ( n227 & n1111 ) | ( n227 & ~n1112 ) | ( n1111 & ~n1112 ) ;
  assign n1114 = ( n1110 & n1112 ) | ( n1110 & ~n1113 ) | ( n1112 & ~n1113 ) ;
  assign n1115 = ( n332 & n338 ) | ( n332 & n344 ) | ( n338 & n344 ) ;
  assign n1116 = ( n332 & n344 ) | ( n332 & ~n1115 ) | ( n344 & ~n1115 ) ;
  assign n1117 = ( n338 & ~n1115 ) | ( n338 & n1116 ) | ( ~n1115 & n1116 ) ;
  assign n1118 = n350 & ~n1117 ;
  assign n1119 = ~n350 & n1117 ;
  assign n1120 = n1118 | n1119 ;
  assign n1121 = n293 & ~n319 ;
  assign n1122 = n293 & n319 ;
  assign n1123 = ( n319 & n1121 ) | ( n319 & ~n1122 ) | ( n1121 & ~n1122 ) ;
  assign n1124 = ( n1114 & n1120 ) | ( n1114 & n1123 ) | ( n1120 & n1123 ) ;
  assign n1125 = ( n1120 & n1123 ) | ( n1120 & ~n1124 ) | ( n1123 & ~n1124 ) ;
  assign n1126 = ( n1114 & ~n1124 ) | ( n1114 & n1125 ) | ( ~n1124 & n1125 ) ;
  assign n1127 = n1109 & ~n1126 ;
  assign n1128 = ~n1109 & n1126 ;
  assign n1129 = n1127 | n1128 ;
  assign n1130 = ~n1106 & n1129 ;
  assign n1131 = ( n1065 & n1088 ) | ( n1065 & ~n1130 ) | ( n1088 & ~n1130 ) ;
  assign n1132 = n1065 & ~n1131 ;
  assign n1133 = ( ~n756 & n760 ) | ( ~n756 & n773 ) | ( n760 & n773 ) ;
  assign n1134 = ( n760 & n773 ) | ( n760 & ~n1133 ) | ( n773 & ~n1133 ) ;
  assign n1135 = ( n756 & n1133 ) | ( n756 & ~n1134 ) | ( n1133 & ~n1134 ) ;
  assign n1136 = ( n750 & ~n764 ) | ( n750 & n767 ) | ( ~n764 & n767 ) ;
  assign n1137 = ( n750 & n767 ) | ( n750 & ~n1136 ) | ( n767 & ~n1136 ) ;
  assign n1138 = ( n764 & n1136 ) | ( n764 & ~n1137 ) | ( n1136 & ~n1137 ) ;
  assign n1139 = x5 & x195 ;
  assign n1140 = x5 | x21 ;
  assign n1141 = ( n778 & ~n1139 ) | ( n778 & n1140 ) | ( ~n1139 & n1140 ) ;
  assign n1142 = ( n778 & n1140 ) | ( n778 & ~n1141 ) | ( n1140 & ~n1141 ) ;
  assign n1143 = ( n1139 & n1141 ) | ( n1139 & ~n1142 ) | ( n1141 & ~n1142 ) ;
  assign n1144 = ( n1135 & n1138 ) | ( n1135 & ~n1143 ) | ( n1138 & ~n1143 ) ;
  assign n1145 = ( ~n1138 & n1143 ) | ( ~n1138 & n1144 ) | ( n1143 & n1144 ) ;
  assign n1146 = ( ~n1135 & n1144 ) | ( ~n1135 & n1145 ) | ( n1144 & n1145 ) ;
  assign n1147 = ( n716 & n724 ) | ( n716 & n734 ) | ( n724 & n734 ) ;
  assign n1148 = ( n716 & n724 ) | ( n716 & ~n1147 ) | ( n724 & ~n1147 ) ;
  assign n1149 = ( n734 & ~n1147 ) | ( n734 & n1148 ) | ( ~n1147 & n1148 ) ;
  assign n1150 = n742 & ~n1149 ;
  assign n1151 = ~n742 & n1149 ;
  assign n1152 = n1150 | n1151 ;
  assign n1153 = ( n891 & ~n892 ) | ( n891 & n895 ) | ( ~n892 & n895 ) ;
  assign n1154 = ( n891 & n895 ) | ( n891 & ~n1153 ) | ( n895 & ~n1153 ) ;
  assign n1155 = ( n892 & n1153 ) | ( n892 & ~n1154 ) | ( n1153 & ~n1154 ) ;
  assign n1156 = x5 & x167 ;
  assign n1157 = x5 | x59 ;
  assign n1158 = ( n906 & ~n1156 ) | ( n906 & n1157 ) | ( ~n1156 & n1157 ) ;
  assign n1159 = ( n906 & n1157 ) | ( n906 & ~n1158 ) | ( n1157 & ~n1158 ) ;
  assign n1160 = ( n1156 & n1158 ) | ( n1156 & ~n1159 ) | ( n1158 & ~n1159 ) ;
  assign n1161 = x5 & x172 ;
  assign n1162 = x5 & ~x173 ;
  assign n1163 = x5 | x174 ;
  assign n1164 = ( ~x5 & n1162 ) | ( ~x5 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1165 = x5 | x166 ;
  assign n1166 = ( ~n1161 & n1164 ) | ( ~n1161 & n1165 ) | ( n1164 & n1165 ) ;
  assign n1167 = ( n1164 & n1165 ) | ( n1164 & ~n1166 ) | ( n1165 & ~n1166 ) ;
  assign n1168 = ( n1161 & n1166 ) | ( n1161 & ~n1167 ) | ( n1166 & ~n1167 ) ;
  assign n1169 = ~n885 & n919 ;
  assign n1170 = n885 & n919 ;
  assign n1171 = ( n885 & n1169 ) | ( n885 & ~n1170 ) | ( n1169 & ~n1170 ) ;
  assign n1172 = ( n1160 & n1168 ) | ( n1160 & n1171 ) | ( n1168 & n1171 ) ;
  assign n1173 = ( n1168 & n1171 ) | ( n1168 & ~n1172 ) | ( n1171 & ~n1172 ) ;
  assign n1174 = ( n1160 & ~n1172 ) | ( n1160 & n1173 ) | ( ~n1172 & n1173 ) ;
  assign n1175 = n1155 & ~n1174 ;
  assign n1176 = ~n1155 & n1174 ;
  assign n1177 = n1175 | n1176 ;
  assign n1178 = ( ~n562 & n566 ) | ( ~n562 & n572 ) | ( n566 & n572 ) ;
  assign n1179 = ( n566 & n572 ) | ( n566 & ~n1178 ) | ( n572 & ~n1178 ) ;
  assign n1180 = ( n562 & n1178 ) | ( n562 & ~n1179 ) | ( n1178 & ~n1179 ) ;
  assign n1181 = x5 & x175 ;
  assign n1182 = x5 | x41 ;
  assign n1183 = ( n578 & ~n1181 ) | ( n578 & n1182 ) | ( ~n1181 & n1182 ) ;
  assign n1184 = ( n578 & n1182 ) | ( n578 & ~n1183 ) | ( n1182 & ~n1183 ) ;
  assign n1185 = ( n1181 & n1183 ) | ( n1181 & ~n1184 ) | ( n1183 & ~n1184 ) ;
  assign n1186 = ( n597 & n605 ) | ( n597 & n616 ) | ( n605 & n616 ) ;
  assign n1187 = ( n597 & n605 ) | ( n597 & ~n1186 ) | ( n605 & ~n1186 ) ;
  assign n1188 = ( n616 & ~n1186 ) | ( n616 & n1187 ) | ( ~n1186 & n1187 ) ;
  assign n1189 = n611 & ~n1188 ;
  assign n1190 = ~n611 & n1188 ;
  assign n1191 = n1189 | n1190 ;
  assign n1192 = ( n558 & ~n586 ) | ( n558 & n589 ) | ( ~n586 & n589 ) ;
  assign n1193 = ( n558 & n589 ) | ( n558 & ~n1192 ) | ( n589 & ~n1192 ) ;
  assign n1194 = ( n586 & n1192 ) | ( n586 & ~n1193 ) | ( n1192 & ~n1193 ) ;
  assign n1195 = ( n1185 & n1191 ) | ( n1185 & n1194 ) | ( n1191 & n1194 ) ;
  assign n1196 = ( n1191 & n1194 ) | ( n1191 & ~n1195 ) | ( n1194 & ~n1195 ) ;
  assign n1197 = ( n1185 & ~n1195 ) | ( n1185 & n1196 ) | ( ~n1195 & n1196 ) ;
  assign n1198 = n1180 & ~n1197 ;
  assign n1199 = ~n1180 & n1197 ;
  assign n1200 = n1198 | n1199 ;
  assign n1201 = n1177 & n1200 ;
  assign n1202 = ( n1146 & n1152 ) | ( n1146 & n1201 ) | ( n1152 & n1201 ) ;
  assign n1203 = ~n640 & n643 ;
  assign n1204 = n640 & n643 ;
  assign n1205 = ( n640 & n1203 ) | ( n640 & ~n1204 ) | ( n1203 & ~n1204 ) ;
  assign n1206 = x5 & x185 ;
  assign n1207 = x5 & ~x186 ;
  assign n1208 = x5 | x31 ;
  assign n1209 = ( ~x5 & n1207 ) | ( ~x5 & n1208 ) | ( n1207 & n1208 ) ;
  assign n1210 = x5 | x30 ;
  assign n1211 = ( ~n1206 & n1209 ) | ( ~n1206 & n1210 ) | ( n1209 & n1210 ) ;
  assign n1212 = ( n1209 & n1210 ) | ( n1209 & ~n1211 ) | ( n1210 & ~n1211 ) ;
  assign n1213 = ( n1206 & n1211 ) | ( n1206 & ~n1212 ) | ( n1211 & ~n1212 ) ;
  assign n1214 = ( n682 & n690 ) | ( n682 & n700 ) | ( n690 & n700 ) ;
  assign n1215 = ( n682 & n690 ) | ( n682 & ~n1214 ) | ( n690 & ~n1214 ) ;
  assign n1216 = ( n700 & ~n1214 ) | ( n700 & n1215 ) | ( ~n1214 & n1215 ) ;
  assign n1217 = n708 & ~n1216 ;
  assign n1218 = ~n708 & n1216 ;
  assign n1219 = n1217 | n1218 ;
  assign n1220 = n632 & ~n666 ;
  assign n1221 = n632 & n666 ;
  assign n1222 = ( n666 & n1220 ) | ( n666 & ~n1221 ) | ( n1220 & ~n1221 ) ;
  assign n1223 = ( n1213 & n1219 ) | ( n1213 & n1222 ) | ( n1219 & n1222 ) ;
  assign n1224 = ( n1219 & n1222 ) | ( n1219 & ~n1223 ) | ( n1222 & ~n1223 ) ;
  assign n1225 = ( n1213 & ~n1223 ) | ( n1213 & n1224 ) | ( ~n1223 & n1224 ) ;
  assign n1226 = n1205 & ~n1225 ;
  assign n1227 = ~n1205 & n1225 ;
  assign n1228 = n1226 | n1227 ;
  assign n1229 = ( n1146 & n1152 ) | ( n1146 & ~n1228 ) | ( n1152 & ~n1228 ) ;
  assign n1230 = n1202 & ~n1229 ;
  assign n1231 = x5 & ~x120 ;
  assign n1232 = ( n780 & n1044 ) | ( n780 & ~n1231 ) | ( n1044 & ~n1231 ) ;
  assign n1233 = ( n780 & n1044 ) | ( n780 & ~n1232 ) | ( n1044 & ~n1232 ) ;
  assign n1234 = ( n1231 & n1232 ) | ( n1231 & ~n1233 ) | ( n1232 & ~n1233 ) ;
  assign n1235 = ~n759 & n775 ;
  assign n1236 = n759 & n775 ;
  assign n1237 = ( n759 & n1235 ) | ( n759 & ~n1236 ) | ( n1235 & ~n1236 ) ;
  assign n1238 = ( n752 & n1234 ) | ( n752 & n1237 ) | ( n1234 & n1237 ) ;
  assign n1239 = ( n1234 & n1237 ) | ( n1234 & ~n1238 ) | ( n1237 & ~n1238 ) ;
  assign n1240 = ( n752 & ~n1238 ) | ( n752 & n1239 ) | ( ~n1238 & n1239 ) ;
  assign n1241 = n766 & ~n1240 ;
  assign n1242 = ~n766 & n1240 ;
  assign n1243 = n1241 | n1242 ;
  assign n1244 = ( n718 & n726 ) | ( n718 & n736 ) | ( n726 & n736 ) ;
  assign n1245 = ( n718 & n726 ) | ( n718 & ~n1244 ) | ( n726 & ~n1244 ) ;
  assign n1246 = ( n736 & ~n1244 ) | ( n736 & n1245 ) | ( ~n1244 & n1245 ) ;
  assign n1247 = n731 & ~n1246 ;
  assign n1248 = ~n731 & n1246 ;
  assign n1249 = n1247 | n1248 ;
  assign n1250 = ~n1243 & n1249 ;
  assign n1251 = n1243 & n1249 ;
  assign n1252 = ( n1243 & n1250 ) | ( n1243 & ~n1251 ) | ( n1250 & ~n1251 ) ;
  assign n1253 = ~n565 & n574 ;
  assign n1254 = n565 & n574 ;
  assign n1255 = ( n565 & n1253 ) | ( n565 & ~n1254 ) | ( n1253 & ~n1254 ) ;
  assign n1256 = x5 & ~x104 ;
  assign n1257 = ( n580 & n1070 ) | ( n580 & ~n1256 ) | ( n1070 & ~n1256 ) ;
  assign n1258 = ( n580 & n1070 ) | ( n580 & ~n1257 ) | ( n1070 & ~n1257 ) ;
  assign n1259 = ( n1256 & n1257 ) | ( n1256 & ~n1258 ) | ( n1257 & ~n1258 ) ;
  assign n1260 = ( n594 & n602 ) | ( n594 & n613 ) | ( n602 & n613 ) ;
  assign n1261 = ( n594 & n602 ) | ( n594 & ~n1260 ) | ( n602 & ~n1260 ) ;
  assign n1262 = ( n613 & ~n1260 ) | ( n613 & n1261 ) | ( ~n1260 & n1261 ) ;
  assign n1263 = n621 & ~n1262 ;
  assign n1264 = ~n621 & n1262 ;
  assign n1265 = n1263 | n1264 ;
  assign n1266 = ~n555 & n588 ;
  assign n1267 = n555 & n588 ;
  assign n1268 = ( n555 & n1266 ) | ( n555 & ~n1267 ) | ( n1266 & ~n1267 ) ;
  assign n1269 = ( n1259 & n1265 ) | ( n1259 & ~n1268 ) | ( n1265 & ~n1268 ) ;
  assign n1270 = ( ~n1265 & n1268 ) | ( ~n1265 & n1269 ) | ( n1268 & n1269 ) ;
  assign n1271 = ( ~n1259 & n1269 ) | ( ~n1259 & n1270 ) | ( n1269 & n1270 ) ;
  assign n1272 = n1255 & n1271 ;
  assign n1273 = n1255 | n1271 ;
  assign n1274 = ~n1272 & n1273 ;
  assign n1275 = x5 & ~n240 ;
  assign n1276 = ~x93 & n1275 ;
  assign n1277 = ( ~x5 & x87 ) | ( ~x5 & x88 ) | ( x87 & x88 ) ;
  assign n1278 = ( x87 & x88 ) | ( x87 & ~n240 ) | ( x88 & ~n240 ) ;
  assign n1279 = ~n1277 & n1278 ;
  assign n1280 = ~n882 & n916 ;
  assign n1281 = n882 & n916 ;
  assign n1282 = ( n882 & n1280 ) | ( n882 & ~n1281 ) | ( n1280 & ~n1281 ) ;
  assign n1283 = ~n894 & n900 ;
  assign n1284 = n894 & n900 ;
  assign n1285 = ( n894 & n1283 ) | ( n894 & ~n1284 ) | ( n1283 & ~n1284 ) ;
  assign n1286 = ( n1279 & n1282 ) | ( n1279 & n1285 ) | ( n1282 & n1285 ) ;
  assign n1287 = ( n1282 & n1285 ) | ( n1282 & ~n1286 ) | ( n1285 & ~n1286 ) ;
  assign n1288 = ( n1279 & ~n1286 ) | ( n1279 & n1287 ) | ( ~n1286 & n1287 ) ;
  assign n1289 = n1276 | n1288 ;
  assign n1290 = n1276 & n1288 ;
  assign n1291 = n1289 & ~n1290 ;
  assign n1292 = n645 & ~n650 ;
  assign n1293 = n645 & n650 ;
  assign n1294 = ( n650 & n1292 ) | ( n650 & ~n1293 ) | ( n1292 & ~n1293 ) ;
  assign n1295 = x5 & ~x131 ;
  assign n1296 = ( n658 & n1111 ) | ( n658 & ~n1295 ) | ( n1111 & ~n1295 ) ;
  assign n1297 = ( n658 & n1111 ) | ( n658 & ~n1296 ) | ( n1111 & ~n1296 ) ;
  assign n1298 = ( n1295 & n1296 ) | ( n1295 & ~n1297 ) | ( n1296 & ~n1297 ) ;
  assign n1299 = ( n684 & n692 ) | ( n684 & n702 ) | ( n692 & n702 ) ;
  assign n1300 = ( n684 & n692 ) | ( n684 & ~n1299 ) | ( n692 & ~n1299 ) ;
  assign n1301 = ( n702 & ~n1299 ) | ( n702 & n1300 ) | ( ~n1299 & n1300 ) ;
  assign n1302 = n697 & ~n1301 ;
  assign n1303 = ~n697 & n1301 ;
  assign n1304 = n1302 | n1303 ;
  assign n1305 = n634 & ~n668 ;
  assign n1306 = n634 & n668 ;
  assign n1307 = ( n668 & n1305 ) | ( n668 & ~n1306 ) | ( n1305 & ~n1306 ) ;
  assign n1308 = ( n1298 & n1304 ) | ( n1298 & n1307 ) | ( n1304 & n1307 ) ;
  assign n1309 = ( n1304 & n1307 ) | ( n1304 & ~n1308 ) | ( n1307 & ~n1308 ) ;
  assign n1310 = ( n1298 & ~n1308 ) | ( n1298 & n1309 ) | ( ~n1308 & n1309 ) ;
  assign n1311 = n1294 & ~n1310 ;
  assign n1312 = ~n1294 & n1310 ;
  assign n1313 = n1311 | n1312 ;
  assign n1314 = ~n1291 & n1313 ;
  assign n1315 = ( n1252 & n1274 ) | ( n1252 & ~n1314 ) | ( n1274 & ~n1314 ) ;
  assign n1316 = n1252 & ~n1315 ;
  assign n1317 = n813 | n878 ;
  assign n1318 = ( ~n803 & n847 ) | ( ~n803 & n1317 ) | ( n847 & n1317 ) ;
  assign n1319 = n803 | n1318 ;
  assign n1320 = ~n929 & n941 ;
  assign n1321 = ( n929 & n1319 ) | ( n929 & ~n1320 ) | ( n1319 & ~n1320 ) ;
  assign n1322 = ( n879 & n880 ) | ( n879 & ~n1321 ) | ( n880 & ~n1321 ) ;
  assign n1323 = ( ~n880 & n1321 ) | ( ~n880 & n1322 ) | ( n1321 & n1322 ) ;
  assign n1324 = ( x11 & ~n879 ) | ( x11 & n1323 ) | ( ~n879 & n1323 ) ;
  assign n1325 = n427 | n460 ;
  assign n1326 = n435 | n1325 ;
  assign n1327 = n251 | n1326 ;
  assign n1328 = ~n251 & n1326 ;
  assign n1329 = ( ~n1326 & n1327 ) | ( ~n1326 & n1328 ) | ( n1327 & n1328 ) ;
  assign n1330 = ~n436 & n486 ;
  assign n1331 = ( n428 & ~n461 ) | ( n428 & n1330 ) | ( ~n461 & n1330 ) ;
  assign n1332 = ~n428 & n1331 ;
  assign n1333 = n542 & n1332 ;
  assign n1334 = n542 & ~n1332 ;
  assign n1335 = ( n1332 & ~n1333 ) | ( n1332 & n1334 ) | ( ~n1333 & n1334 ) ;
  assign n1336 = x48 | n679 ;
  assign n1337 = ( n679 & n809 ) | ( n679 & n1336 ) | ( n809 & n1336 ) ;
  assign n1338 = n713 | n800 ;
  assign n1339 = ( n800 & n1337 ) | ( n800 & n1338 ) | ( n1337 & n1338 ) ;
  assign n1340 = n788 | n834 ;
  assign n1341 = ( n834 & n1339 ) | ( n834 & n1340 ) | ( n1339 & n1340 ) ;
  assign n1342 = n845 | n1341 ;
  assign n1343 = ( n747 & n845 ) | ( n747 & n1342 ) | ( n845 & n1342 ) ;
  assign n1344 = n486 & ~n970 ;
  assign n1345 = ( n962 & ~n971 ) | ( n962 & n1344 ) | ( ~n971 & n1344 ) ;
  assign n1346 = ~n962 & n1345 ;
  assign n1347 = n525 & ~n975 ;
  assign n1348 = ( n525 & n1346 ) | ( n525 & n1347 ) | ( n1346 & n1347 ) ;
  assign n1349 = n528 & n1348 ;
  assign n1350 = ~n528 & n536 ;
  assign n1351 = ( ~n528 & n532 ) | ( ~n528 & n1350 ) | ( n532 & n1350 ) ;
  assign n1352 = ~n1348 & n1351 ;
  assign n1353 = ( n1348 & ~n1349 ) | ( n1348 & n1352 ) | ( ~n1349 & n1352 ) ;
  assign n1354 = ~n262 & n462 ;
  assign n1355 = ~n239 & n1328 ;
  assign n1356 = ~n262 & n1355 ;
  assign n1357 = n238 & ~n262 ;
  assign n1358 = n469 | n1357 ;
  assign n1359 = ( ~x179 & n254 ) | ( ~x179 & n1358 ) | ( n254 & n1358 ) ;
  assign n1360 = ( ~n1354 & n1356 ) | ( ~n1354 & n1359 ) | ( n1356 & n1359 ) ;
  assign n1361 = n257 & ~n1359 ;
  assign n1362 = ( n1354 & n1360 ) | ( n1354 & ~n1361 ) | ( n1360 & ~n1361 ) ;
  assign n1363 = n245 & ~n1362 ;
  assign n1364 = n245 & n1362 ;
  assign n1365 = ( n1362 & n1363 ) | ( n1362 & ~n1364 ) | ( n1363 & ~n1364 ) ;
  assign n1366 = n1354 | n1356 ;
  assign n1367 = n1358 | n1366 ;
  assign n1368 = n257 & n1367 ;
  assign n1369 = n257 | n1367 ;
  assign n1370 = ~n1368 & n1369 ;
  assign n1371 = ( ~x177 & n236 ) | ( ~x177 & n250 ) | ( n236 & n250 ) ;
  assign n1372 = n1328 | n1371 ;
  assign n1373 = ( ~n239 & n1371 ) | ( ~n239 & n1372 ) | ( n1371 & n1372 ) ;
  assign n1374 = ~n262 & n1373 ;
  assign n1375 = n262 | n1373 ;
  assign n1376 = ( ~n1373 & n1374 ) | ( ~n1373 & n1375 ) | ( n1374 & n1375 ) ;
  assign n1377 = n250 & ~n1328 ;
  assign n1378 = ( n239 & ~n1328 ) | ( n239 & n1377 ) | ( ~n1328 & n1377 ) ;
  assign n1379 = ( n239 & n1328 ) | ( n239 & n1377 ) | ( n1328 & n1377 ) ;
  assign n1380 = ( n1328 & n1378 ) | ( n1328 & ~n1379 ) | ( n1378 & ~n1379 ) ;
  assign n1381 = n491 & ~n504 ;
  assign n1382 = n496 & n1381 ;
  assign n1383 = n491 & n1334 ;
  assign n1384 = n496 & n1383 ;
  assign n1385 = ~x169 & n508 ;
  assign n1386 = n513 & ~n1385 ;
  assign n1387 = ( x170 & n515 ) | ( x170 & n1386 ) | ( n515 & n1386 ) ;
  assign n1388 = ( n1382 & ~n1384 ) | ( n1382 & n1387 ) | ( ~n1384 & n1387 ) ;
  assign n1389 = ~n519 & n1387 ;
  assign n1390 = ( ~n1382 & n1388 ) | ( ~n1382 & n1389 ) | ( n1388 & n1389 ) ;
  assign n1391 = n501 & n1390 ;
  assign n1392 = n501 & ~n1390 ;
  assign n1393 = ( n1390 & ~n1391 ) | ( n1390 & n1392 ) | ( ~n1391 & n1392 ) ;
  assign n1394 = n1382 | n1384 ;
  assign n1395 = n1386 & ~n1394 ;
  assign n1396 = n519 | n1395 ;
  assign n1397 = n519 & n1395 ;
  assign n1398 = n1396 & ~n1397 ;
  assign n1399 = ( x169 & n488 ) | ( x169 & n504 ) | ( n488 & n504 ) ;
  assign n1400 = ~n1334 & n1399 ;
  assign n1401 = ( ~n491 & n1399 ) | ( ~n491 & n1400 ) | ( n1399 & n1400 ) ;
  assign n1402 = n496 & ~n1401 ;
  assign n1403 = n496 & n1401 ;
  assign n1404 = ( n1401 & n1402 ) | ( n1401 & ~n1403 ) | ( n1402 & ~n1403 ) ;
  assign n1405 = n504 | n1334 ;
  assign n1406 = ( n491 & n1334 ) | ( n491 & n1405 ) | ( n1334 & n1405 ) ;
  assign n1407 = ( n491 & ~n1334 ) | ( n491 & n1405 ) | ( ~n1334 & n1405 ) ;
  assign n1408 = ( n1334 & ~n1406 ) | ( n1334 & n1407 ) | ( ~n1406 & n1407 ) ;
  assign n1409 = n214 & n220 ;
  assign n1410 = ( ~n211 & n217 ) | ( ~n211 & n1409 ) | ( n217 & n1409 ) ;
  assign n1411 = n211 & n1410 ;
  assign n1412 = n1230 & n1411 ;
  assign n1413 = ( ~n1132 & n1316 ) | ( ~n1132 & n1412 ) | ( n1316 & n1412 ) ;
  assign n1414 = n1132 & n1413 ;
  assign n1415 = n525 & ~n546 ;
  assign n1416 = ( n525 & n1332 ) | ( n525 & n1415 ) | ( n1332 & n1415 ) ;
  assign n1417 = n528 & n1416 ;
  assign n1418 = n1351 & ~n1416 ;
  assign n1419 = ( n1416 & ~n1417 ) | ( n1416 & n1418 ) | ( ~n1417 & n1418 ) ;
  assign n1420 = ~x181 & n478 ;
  assign n1421 = n279 & ~n1420 ;
  assign n1422 = ( x183 & n273 ) | ( x183 & n1421 ) | ( n273 & n1421 ) ;
  assign n1423 = ~n266 & n476 ;
  assign n1424 = ( n476 & ~n1326 ) | ( n476 & n1423 ) | ( ~n1326 & n1423 ) ;
  assign n1425 = ~n1422 & n1424 ;
  assign n1426 = n276 & n281 ;
  assign n1427 = ( ~n283 & n285 ) | ( ~n283 & n1426 ) | ( n285 & n1426 ) ;
  assign n1428 = ( x183 & n273 ) | ( x183 & n279 ) | ( n273 & n279 ) ;
  assign n1429 = ~n1427 & n1428 ;
  assign n1430 = n1424 | n1429 ;
  assign n1431 = ( n271 & ~n1425 ) | ( n271 & n1430 ) | ( ~n1425 & n1430 ) ;
  assign n1432 = ( n271 & n1430 ) | ( n271 & ~n1431 ) | ( n1430 & ~n1431 ) ;
  assign n1433 = ( n1425 & n1431 ) | ( n1425 & ~n1432 ) | ( n1431 & ~n1432 ) ;
  assign n1434 = ~n1421 & n1424 ;
  assign n1435 = ~n286 & n1421 ;
  assign n1436 = ( ~n281 & n1421 ) | ( ~n281 & n1435 ) | ( n1421 & n1435 ) ;
  assign n1437 = n1424 | n1436 ;
  assign n1438 = ( n276 & ~n1434 ) | ( n276 & n1437 ) | ( ~n1434 & n1437 ) ;
  assign n1439 = ( n276 & n1437 ) | ( n276 & ~n1438 ) | ( n1437 & ~n1438 ) ;
  assign n1440 = ( n1434 & n1438 ) | ( n1434 & ~n1439 ) | ( n1438 & ~n1439 ) ;
  assign n1441 = ( x181 & n283 ) | ( x181 & n1424 ) | ( n283 & n1424 ) ;
  assign n1442 = n281 | n1441 ;
  assign n1443 = n281 & n1441 ;
  assign n1444 = n1442 & ~n1443 ;
  assign n1445 = n286 & n1424 ;
  assign n1446 = n286 & ~n1424 ;
  assign n1447 = ( n1424 & ~n1445 ) | ( n1424 & n1446 ) | ( ~n1445 & n1446 ) ;
  assign n1448 = n356 & ~n425 ;
  assign n1449 = ( n425 & n1018 ) | ( n425 & ~n1448 ) | ( n1018 & ~n1448 ) ;
  assign n1450 = n374 | n1449 ;
  assign n1451 = ~n374 & n1449 ;
  assign n1452 = ( ~n1449 & n1450 ) | ( ~n1449 & n1451 ) | ( n1450 & n1451 ) ;
  assign n1453 = ( ~x11 & n529 ) | ( ~x11 & n1416 ) | ( n529 & n1416 ) ;
  assign n1454 = n536 & ~n1453 ;
  assign n1455 = ~n536 & n1453 ;
  assign n1456 = n1454 | n1455 ;
  assign n1457 = ~n532 & n1416 ;
  assign n1458 = n532 | n1416 ;
  assign n1459 = ( ~n1416 & n1457 ) | ( ~n1416 & n1458 ) | ( n1457 & n1458 ) ;
  assign n1460 = ~n362 & n373 ;
  assign n1461 = ~n385 & n1460 ;
  assign n1462 = ~n362 & n1451 ;
  assign n1463 = ~n385 & n1462 ;
  assign n1464 = n361 & ~n385 ;
  assign n1465 = n444 | n1464 ;
  assign n1466 = ( ~x199 & n377 ) | ( ~x199 & n1465 ) | ( n377 & n1465 ) ;
  assign n1467 = ( ~n1461 & n1463 ) | ( ~n1461 & n1466 ) | ( n1463 & n1466 ) ;
  assign n1468 = n380 & ~n1466 ;
  assign n1469 = ( n1461 & n1467 ) | ( n1461 & ~n1468 ) | ( n1467 & ~n1468 ) ;
  assign n1470 = n368 | n1469 ;
  assign n1471 = ~n368 & n1469 ;
  assign n1472 = ( ~n1469 & n1470 ) | ( ~n1469 & n1471 ) | ( n1470 & n1471 ) ;
  assign n1473 = n1461 | n1463 ;
  assign n1474 = n1465 | n1473 ;
  assign n1475 = n380 & n1474 ;
  assign n1476 = n380 | n1474 ;
  assign n1477 = ~n1475 & n1476 ;
  assign n1478 = ( ~x197 & n359 ) | ( ~x197 & n373 ) | ( n359 & n373 ) ;
  assign n1479 = n1451 | n1478 ;
  assign n1480 = ( ~n362 & n1478 ) | ( ~n362 & n1479 ) | ( n1478 & n1479 ) ;
  assign n1481 = ~n385 & n1480 ;
  assign n1482 = n385 | n1480 ;
  assign n1483 = ( ~n1480 & n1481 ) | ( ~n1480 & n1482 ) | ( n1481 & n1482 ) ;
  assign n1484 = n373 & ~n1451 ;
  assign n1485 = ( n362 & ~n1451 ) | ( n362 & n1484 ) | ( ~n1451 & n1484 ) ;
  assign n1486 = ( n362 & n1451 ) | ( n362 & n1484 ) | ( n1451 & n1484 ) ;
  assign n1487 = ( n1451 & n1485 ) | ( n1451 & ~n1486 ) | ( n1485 & ~n1486 ) ;
  assign n1488 = ~n407 & n412 ;
  assign n1489 = ( n400 & n406 ) | ( n400 & ~n1488 ) | ( n406 & ~n1488 ) ;
  assign n1490 = ~n400 & n401 ;
  assign n1491 = ( n1488 & n1489 ) | ( n1488 & ~n1490 ) | ( n1489 & ~n1490 ) ;
  assign n1492 = n389 & ~n451 ;
  assign n1493 = ( n451 & n1449 ) | ( n451 & ~n1492 ) | ( n1449 & ~n1492 ) ;
  assign n1494 = n1491 & ~n1493 ;
  assign n1495 = n401 | n407 ;
  assign n1496 = ( ~n410 & n411 ) | ( ~n410 & n1495 ) | ( n411 & n1495 ) ;
  assign n1497 = ( ~x203 & n398 ) | ( ~x203 & n406 ) | ( n398 & n406 ) ;
  assign n1498 = n1496 & ~n1497 ;
  assign n1499 = n1493 & ~n1498 ;
  assign n1500 = ( n395 & n1494 ) | ( n395 & n1499 ) | ( n1494 & n1499 ) ;
  assign n1501 = ( n395 & n1499 ) | ( n395 & ~n1500 ) | ( n1499 & ~n1500 ) ;
  assign n1502 = ( n1494 & ~n1500 ) | ( n1494 & n1501 ) | ( ~n1500 & n1501 ) ;
  assign n1503 = n406 | n1488 ;
  assign n1504 = ~n1493 & n1503 ;
  assign n1505 = n413 & ~n1503 ;
  assign n1506 = ( n407 & ~n1503 ) | ( n407 & n1505 ) | ( ~n1503 & n1505 ) ;
  assign n1507 = n1493 & ~n1506 ;
  assign n1508 = ( n401 & n1504 ) | ( n401 & n1507 ) | ( n1504 & n1507 ) ;
  assign n1509 = ( n401 & n1507 ) | ( n401 & ~n1508 ) | ( n1507 & ~n1508 ) ;
  assign n1510 = ( n1504 & ~n1508 ) | ( n1504 & n1509 ) | ( ~n1508 & n1509 ) ;
  assign n1511 = ( ~x201 & n410 ) | ( ~x201 & n1493 ) | ( n410 & n1493 ) ;
  assign n1512 = n407 & n1511 ;
  assign n1513 = n407 | n1511 ;
  assign n1514 = ~n1512 & n1513 ;
  assign n1515 = n413 | n1493 ;
  assign n1516 = ~n413 & n1493 ;
  assign n1517 = ( ~n1493 & n1515 ) | ( ~n1493 & n1516 ) | ( n1515 & n1516 ) ;
  assign n1518 = x181 & n283 ;
  assign n1519 = ( n1421 & n1422 ) | ( n1421 & ~n1518 ) | ( n1422 & ~n1518 ) ;
  assign n1520 = ( ~n1422 & n1518 ) | ( ~n1422 & n1519 ) | ( n1518 & n1519 ) ;
  assign n1521 = ( ~n1421 & n1519 ) | ( ~n1421 & n1520 ) | ( n1519 & n1520 ) ;
  assign n1522 = ( n271 & n281 ) | ( n271 & ~n1521 ) | ( n281 & ~n1521 ) ;
  assign n1523 = ( ~n271 & n1521 ) | ( ~n271 & n1522 ) | ( n1521 & n1522 ) ;
  assign n1524 = ( ~n281 & n1522 ) | ( ~n281 & n1523 ) | ( n1522 & n1523 ) ;
  assign n1525 = n276 & n1524 ;
  assign n1526 = n276 | n1524 ;
  assign n1527 = ~n1525 & n1526 ;
  assign n1528 = n460 | n957 ;
  assign n1529 = n969 | n1528 ;
  assign n1530 = ( n476 & n1527 ) | ( n476 & n1529 ) | ( n1527 & n1529 ) ;
  assign n1531 = ( n284 & n1429 ) | ( n284 & n1436 ) | ( n1429 & n1436 ) ;
  assign n1532 = ( n284 & n1436 ) | ( n284 & ~n1531 ) | ( n1436 & ~n1531 ) ;
  assign n1533 = ( n1429 & ~n1531 ) | ( n1429 & n1532 ) | ( ~n1531 & n1532 ) ;
  assign n1534 = ( n271 & n281 ) | ( n271 & n1533 ) | ( n281 & n1533 ) ;
  assign n1535 = ( n271 & n1533 ) | ( n271 & ~n1534 ) | ( n1533 & ~n1534 ) ;
  assign n1536 = ( n281 & ~n1534 ) | ( n281 & n1535 ) | ( ~n1534 & n1535 ) ;
  assign n1537 = n276 & ~n1536 ;
  assign n1538 = ~n276 & n1536 ;
  assign n1539 = n1537 | n1538 ;
  assign n1540 = ( n476 & ~n1529 ) | ( n476 & n1539 ) | ( ~n1529 & n1539 ) ;
  assign n1541 = ~n1530 & n1540 ;
  assign n1542 = ( n1354 & n1359 ) | ( n1354 & ~n1361 ) | ( n1359 & ~n1361 ) ;
  assign n1543 = ~n1354 & n1358 ;
  assign n1544 = ( n250 & ~n1354 ) | ( n250 & n1543 ) | ( ~n1354 & n1543 ) ;
  assign n1545 = ( n250 & n1354 ) | ( n250 & n1543 ) | ( n1354 & n1543 ) ;
  assign n1546 = ( n1354 & n1544 ) | ( n1354 & ~n1545 ) | ( n1544 & ~n1545 ) ;
  assign n1547 = ( n1371 & n1542 ) | ( n1371 & ~n1546 ) | ( n1542 & ~n1546 ) ;
  assign n1548 = ( ~n1542 & n1546 ) | ( ~n1542 & n1547 ) | ( n1546 & n1547 ) ;
  assign n1549 = ( ~n1371 & n1547 ) | ( ~n1371 & n1548 ) | ( n1547 & n1548 ) ;
  assign n1550 = ~n251 & n1549 ;
  assign n1551 = n251 & ~n1549 ;
  assign n1552 = n1550 | n1551 ;
  assign n1553 = ( ~n239 & n245 ) | ( ~n239 & n1552 ) | ( n245 & n1552 ) ;
  assign n1554 = ( n245 & n1552 ) | ( n245 & ~n1553 ) | ( n1552 & ~n1553 ) ;
  assign n1555 = ( n239 & n1553 ) | ( n239 & ~n1554 ) | ( n1553 & ~n1554 ) ;
  assign n1556 = ~n262 & n1555 ;
  assign n1557 = n262 & ~n1555 ;
  assign n1558 = n1556 | n1557 ;
  assign n1559 = ~n1529 & n1558 ;
  assign n1560 = n239 & ~n1371 ;
  assign n1561 = ( n251 & ~n1371 ) | ( n251 & n1560 ) | ( ~n1371 & n1560 ) ;
  assign n1562 = x176 & ~n248 ;
  assign n1563 = n1358 & ~n1562 ;
  assign n1564 = n251 | n262 ;
  assign n1565 = n239 & ~n1354 ;
  assign n1566 = ( ~n1354 & n1564 ) | ( ~n1354 & n1565 ) | ( n1564 & n1565 ) ;
  assign n1567 = ~n1562 & n1566 ;
  assign n1568 = ( n1358 & n1562 ) | ( n1358 & ~n1566 ) | ( n1562 & ~n1566 ) ;
  assign n1569 = ( ~n1563 & n1567 ) | ( ~n1563 & n1568 ) | ( n1567 & n1568 ) ;
  assign n1570 = n1561 | n1569 ;
  assign n1571 = n1561 & ~n1569 ;
  assign n1572 = ( ~n1561 & n1570 ) | ( ~n1561 & n1571 ) | ( n1570 & n1571 ) ;
  assign n1573 = ( ~n239 & n257 ) | ( ~n239 & n1564 ) | ( n257 & n1564 ) ;
  assign n1574 = ~n257 & n1354 ;
  assign n1575 = ( n239 & n1573 ) | ( n239 & ~n1574 ) | ( n1573 & ~n1574 ) ;
  assign n1576 = ~n1359 & n1575 ;
  assign n1577 = ( ~n251 & n1572 ) | ( ~n251 & n1576 ) | ( n1572 & n1576 ) ;
  assign n1578 = ( n1572 & n1576 ) | ( n1572 & ~n1577 ) | ( n1576 & ~n1577 ) ;
  assign n1579 = ( n251 & n1577 ) | ( n251 & ~n1578 ) | ( n1577 & ~n1578 ) ;
  assign n1580 = ( ~n239 & n245 ) | ( ~n239 & n1579 ) | ( n245 & n1579 ) ;
  assign n1581 = ( n245 & n1579 ) | ( n245 & ~n1580 ) | ( n1579 & ~n1580 ) ;
  assign n1582 = ( n239 & n1580 ) | ( n239 & ~n1581 ) | ( n1580 & ~n1581 ) ;
  assign n1583 = ~n262 & n1582 ;
  assign n1584 = n262 & ~n1582 ;
  assign n1585 = n1583 | n1584 ;
  assign n1586 = n1529 & ~n1585 ;
  assign n1587 = ( n257 & n1559 ) | ( n257 & n1586 ) | ( n1559 & n1586 ) ;
  assign n1588 = ( n257 & n1586 ) | ( n257 & ~n1587 ) | ( n1586 & ~n1587 ) ;
  assign n1589 = ( n1559 & ~n1587 ) | ( n1559 & n1588 ) | ( ~n1587 & n1588 ) ;
  assign n1590 = n476 & ~n960 ;
  assign n1591 = ( n1529 & n1539 ) | ( n1529 & n1590 ) | ( n1539 & n1590 ) ;
  assign n1592 = ( n1527 & ~n1529 ) | ( n1527 & n1590 ) | ( ~n1529 & n1590 ) ;
  assign n1593 = n1591 & ~n1592 ;
  assign n1594 = ~n1541 & n1593 ;
  assign n1595 = ( n1541 & n1589 ) | ( n1541 & ~n1594 ) | ( n1589 & ~n1594 ) ;
  assign n1596 = ( n1541 & ~n1589 ) | ( n1541 & n1594 ) | ( ~n1589 & n1594 ) ;
  assign n1597 = ( ~n1541 & n1595 ) | ( ~n1541 & n1596 ) | ( n1595 & n1596 ) ;
  assign n1598 = x11 | x206 ;
  assign n1599 = ( x11 & x172 ) | ( x11 & x206 ) | ( x172 & x206 ) ;
  assign n1600 = x173 & ~n1599 ;
  assign n1601 = ( x173 & x206 ) | ( x173 & ~n1599 ) | ( x206 & ~n1599 ) ;
  assign n1602 = ( n1598 & n1600 ) | ( n1598 & ~n1601 ) | ( n1600 & ~n1601 ) ;
  assign n1603 = ( ~n525 & n1346 ) | ( ~n525 & n1602 ) | ( n1346 & n1602 ) ;
  assign n1604 = ( x11 & x172 ) | ( x11 & ~x206 ) | ( x172 & ~x206 ) ;
  assign n1605 = ~x173 & n1604 ;
  assign n1606 = ( ~x173 & x206 ) | ( ~x173 & n1604 ) | ( x206 & n1604 ) ;
  assign n1607 = ( x206 & n1605 ) | ( x206 & ~n1606 ) | ( n1605 & ~n1606 ) ;
  assign n1608 = ( n525 & n1346 ) | ( n525 & n1607 ) | ( n1346 & n1607 ) ;
  assign n1609 = n1603 & n1608 ;
  assign n1610 = ( ~n1382 & n1387 ) | ( ~n1382 & n1389 ) | ( n1387 & n1389 ) ;
  assign n1611 = n1382 | n1386 ;
  assign n1612 = ( n504 & n1382 ) | ( n504 & n1611 ) | ( n1382 & n1611 ) ;
  assign n1613 = ( n504 & ~n1382 ) | ( n504 & n1611 ) | ( ~n1382 & n1611 ) ;
  assign n1614 = ( n1382 & ~n1612 ) | ( n1382 & n1613 ) | ( ~n1612 & n1613 ) ;
  assign n1615 = ( n1399 & n1610 ) | ( n1399 & n1614 ) | ( n1610 & n1614 ) ;
  assign n1616 = ( n1610 & n1614 ) | ( n1610 & ~n1615 ) | ( n1614 & ~n1615 ) ;
  assign n1617 = ( n1399 & ~n1615 ) | ( n1399 & n1616 ) | ( ~n1615 & n1616 ) ;
  assign n1618 = n542 & n1617 ;
  assign n1619 = n542 | n1617 ;
  assign n1620 = ~n1618 & n1619 ;
  assign n1621 = ( n491 & n501 ) | ( n491 & ~n1620 ) | ( n501 & ~n1620 ) ;
  assign n1622 = ( ~n491 & n1620 ) | ( ~n491 & n1621 ) | ( n1620 & n1621 ) ;
  assign n1623 = ( ~n501 & n1621 ) | ( ~n501 & n1622 ) | ( n1621 & n1622 ) ;
  assign n1624 = n496 & n1623 ;
  assign n1625 = n496 | n1623 ;
  assign n1626 = ~n1624 & n1625 ;
  assign n1627 = n1346 & ~n1626 ;
  assign n1628 = ~n491 & n1399 ;
  assign n1629 = ( ~n542 & n1399 ) | ( ~n542 & n1628 ) | ( n1399 & n1628 ) ;
  assign n1630 = x168 & n503 ;
  assign n1631 = n1386 | n1630 ;
  assign n1632 = n496 & n542 ;
  assign n1633 = n491 | n1382 ;
  assign n1634 = ( n1382 & n1632 ) | ( n1382 & n1633 ) | ( n1632 & n1633 ) ;
  assign n1635 = n1630 | n1634 ;
  assign n1636 = ( ~n1386 & n1630 ) | ( ~n1386 & n1634 ) | ( n1630 & n1634 ) ;
  assign n1637 = ( n1631 & ~n1635 ) | ( n1631 & n1636 ) | ( ~n1635 & n1636 ) ;
  assign n1638 = n1629 | n1637 ;
  assign n1639 = n1629 & ~n1637 ;
  assign n1640 = ( ~n1629 & n1638 ) | ( ~n1629 & n1639 ) | ( n1638 & n1639 ) ;
  assign n1641 = ( ~n491 & n519 ) | ( ~n491 & n1632 ) | ( n519 & n1632 ) ;
  assign n1642 = n519 & n1382 ;
  assign n1643 = ( n491 & n1641 ) | ( n491 & n1642 ) | ( n1641 & n1642 ) ;
  assign n1644 = n1387 & ~n1643 ;
  assign n1645 = ( n542 & n1640 ) | ( n542 & n1644 ) | ( n1640 & n1644 ) ;
  assign n1646 = ( n1640 & n1644 ) | ( n1640 & ~n1645 ) | ( n1644 & ~n1645 ) ;
  assign n1647 = ( n542 & ~n1645 ) | ( n542 & n1646 ) | ( ~n1645 & n1646 ) ;
  assign n1648 = ( n491 & n501 ) | ( n491 & ~n1647 ) | ( n501 & ~n1647 ) ;
  assign n1649 = ( ~n491 & n1647 ) | ( ~n491 & n1648 ) | ( n1647 & n1648 ) ;
  assign n1650 = ( ~n501 & n1648 ) | ( ~n501 & n1649 ) | ( n1648 & n1649 ) ;
  assign n1651 = n496 & n1650 ;
  assign n1652 = n496 | n1650 ;
  assign n1653 = ~n1651 & n1652 ;
  assign n1654 = ~n1346 & n1653 ;
  assign n1655 = ( ~n519 & n1627 ) | ( ~n519 & n1654 ) | ( n1627 & n1654 ) ;
  assign n1656 = ( n519 & ~n1654 ) | ( n519 & n1655 ) | ( ~n1654 & n1655 ) ;
  assign n1657 = ( ~n1627 & n1655 ) | ( ~n1627 & n1656 ) | ( n1655 & n1656 ) ;
  assign n1658 = ( ~n1346 & n1347 ) | ( ~n1346 & n1607 ) | ( n1347 & n1607 ) ;
  assign n1659 = ( n1346 & n1347 ) | ( n1346 & ~n1602 ) | ( n1347 & ~n1602 ) ;
  assign n1660 = n1658 & ~n1659 ;
  assign n1661 = ~n1609 & n1660 ;
  assign n1662 = ( ~n1609 & n1657 ) | ( ~n1609 & n1661 ) | ( n1657 & n1661 ) ;
  assign n1663 = ( n1609 & n1657 ) | ( n1609 & n1661 ) | ( n1657 & n1661 ) ;
  assign n1664 = ( n1609 & n1662 ) | ( n1609 & ~n1663 ) | ( n1662 & ~n1663 ) ;
  assign n1665 = x201 & ~n410 ;
  assign n1666 = ( n1491 & n1503 ) | ( n1491 & n1665 ) | ( n1503 & n1665 ) ;
  assign n1667 = ( n1491 & n1665 ) | ( n1491 & ~n1666 ) | ( n1665 & ~n1666 ) ;
  assign n1668 = ( n1503 & ~n1666 ) | ( n1503 & n1667 ) | ( ~n1666 & n1667 ) ;
  assign n1669 = ( n395 & n407 ) | ( n395 & n1668 ) | ( n407 & n1668 ) ;
  assign n1670 = ( n395 & n1668 ) | ( n395 & ~n1669 ) | ( n1668 & ~n1669 ) ;
  assign n1671 = ( n407 & ~n1669 ) | ( n407 & n1670 ) | ( ~n1669 & n1670 ) ;
  assign n1672 = ~n401 & n1671 ;
  assign n1673 = n401 & ~n1671 ;
  assign n1674 = n1672 | n1673 ;
  assign n1675 = ( n329 & ~n966 ) | ( n329 & n1017 ) | ( ~n966 & n1017 ) ;
  assign n1676 = ( n425 & ~n1448 ) | ( n425 & n1675 ) | ( ~n1448 & n1675 ) ;
  assign n1677 = ( n451 & n1674 ) | ( n451 & ~n1676 ) | ( n1674 & ~n1676 ) ;
  assign n1678 = ( ~n412 & n1498 ) | ( ~n412 & n1506 ) | ( n1498 & n1506 ) ;
  assign n1679 = ( n412 & ~n1506 ) | ( n412 & n1678 ) | ( ~n1506 & n1678 ) ;
  assign n1680 = ( ~n1498 & n1678 ) | ( ~n1498 & n1679 ) | ( n1678 & n1679 ) ;
  assign n1681 = ( n395 & n407 ) | ( n395 & n1680 ) | ( n407 & n1680 ) ;
  assign n1682 = ( n395 & n1680 ) | ( n395 & ~n1681 ) | ( n1680 & ~n1681 ) ;
  assign n1683 = ( n407 & ~n1681 ) | ( n407 & n1682 ) | ( ~n1681 & n1682 ) ;
  assign n1684 = ~n401 & n1683 ;
  assign n1685 = n401 & ~n1683 ;
  assign n1686 = n1684 | n1685 ;
  assign n1687 = ( n451 & n1676 ) | ( n451 & ~n1686 ) | ( n1676 & ~n1686 ) ;
  assign n1688 = n1677 & ~n1687 ;
  assign n1689 = ( n1461 & n1466 ) | ( n1461 & ~n1468 ) | ( n1466 & ~n1468 ) ;
  assign n1690 = ~n1461 & n1465 ;
  assign n1691 = ( n373 & ~n1461 ) | ( n373 & n1690 ) | ( ~n1461 & n1690 ) ;
  assign n1692 = ( n373 & n1461 ) | ( n373 & n1690 ) | ( n1461 & n1690 ) ;
  assign n1693 = ( n1461 & n1691 ) | ( n1461 & ~n1692 ) | ( n1691 & ~n1692 ) ;
  assign n1694 = ( n1478 & n1689 ) | ( n1478 & ~n1693 ) | ( n1689 & ~n1693 ) ;
  assign n1695 = ( ~n1689 & n1693 ) | ( ~n1689 & n1694 ) | ( n1693 & n1694 ) ;
  assign n1696 = ( ~n1478 & n1694 ) | ( ~n1478 & n1695 ) | ( n1694 & n1695 ) ;
  assign n1697 = ~n374 & n1696 ;
  assign n1698 = n374 & ~n1696 ;
  assign n1699 = n1697 | n1698 ;
  assign n1700 = ( n362 & n368 ) | ( n362 & ~n1699 ) | ( n368 & ~n1699 ) ;
  assign n1701 = ( ~n362 & n1699 ) | ( ~n362 & n1700 ) | ( n1699 & n1700 ) ;
  assign n1702 = ( ~n368 & n1700 ) | ( ~n368 & n1701 ) | ( n1700 & n1701 ) ;
  assign n1703 = n385 | n1702 ;
  assign n1704 = n385 & n1702 ;
  assign n1705 = n1703 & ~n1704 ;
  assign n1706 = n1676 | n1705 ;
  assign n1707 = n362 & ~n1478 ;
  assign n1708 = ( n374 & ~n1478 ) | ( n374 & n1707 ) | ( ~n1478 & n1707 ) ;
  assign n1709 = x196 & ~n371 ;
  assign n1710 = n1465 & ~n1709 ;
  assign n1711 = n374 | n385 ;
  assign n1712 = n362 & ~n1461 ;
  assign n1713 = ( ~n1461 & n1711 ) | ( ~n1461 & n1712 ) | ( n1711 & n1712 ) ;
  assign n1714 = ~n1709 & n1713 ;
  assign n1715 = ( n1465 & n1709 ) | ( n1465 & ~n1713 ) | ( n1709 & ~n1713 ) ;
  assign n1716 = ( ~n1710 & n1714 ) | ( ~n1710 & n1715 ) | ( n1714 & n1715 ) ;
  assign n1717 = n1708 | n1716 ;
  assign n1718 = n1708 & ~n1716 ;
  assign n1719 = ( ~n1708 & n1717 ) | ( ~n1708 & n1718 ) | ( n1717 & n1718 ) ;
  assign n1720 = ( ~n362 & n380 ) | ( ~n362 & n1711 ) | ( n380 & n1711 ) ;
  assign n1721 = ~n380 & n1461 ;
  assign n1722 = ( n362 & n1720 ) | ( n362 & ~n1721 ) | ( n1720 & ~n1721 ) ;
  assign n1723 = ~n1466 & n1722 ;
  assign n1724 = ( ~n374 & n1719 ) | ( ~n374 & n1723 ) | ( n1719 & n1723 ) ;
  assign n1725 = ( n1719 & n1723 ) | ( n1719 & ~n1724 ) | ( n1723 & ~n1724 ) ;
  assign n1726 = ( n374 & n1724 ) | ( n374 & ~n1725 ) | ( n1724 & ~n1725 ) ;
  assign n1727 = ( n362 & n368 ) | ( n362 & ~n1726 ) | ( n368 & ~n1726 ) ;
  assign n1728 = ( ~n362 & n1726 ) | ( ~n362 & n1727 ) | ( n1726 & n1727 ) ;
  assign n1729 = ( ~n368 & n1727 ) | ( ~n368 & n1728 ) | ( n1727 & n1728 ) ;
  assign n1730 = n385 | n1729 ;
  assign n1731 = n385 & n1729 ;
  assign n1732 = n1730 & ~n1731 ;
  assign n1733 = n1676 & n1732 ;
  assign n1734 = ( n380 & ~n1706 ) | ( n380 & n1733 ) | ( ~n1706 & n1733 ) ;
  assign n1735 = ( n380 & n1733 ) | ( n380 & ~n1734 ) | ( n1733 & ~n1734 ) ;
  assign n1736 = ( n1706 & n1734 ) | ( n1706 & ~n1735 ) | ( n1734 & ~n1735 ) ;
  assign n1737 = ~n451 & n953 ;
  assign n1738 = ( n1676 & n1686 ) | ( n1676 & n1737 ) | ( n1686 & n1737 ) ;
  assign n1739 = ( n1674 & n1676 ) | ( n1674 & ~n1737 ) | ( n1676 & ~n1737 ) ;
  assign n1740 = n1738 & n1739 ;
  assign n1741 = ~n1688 & n1740 ;
  assign n1742 = ( ~n1688 & n1736 ) | ( ~n1688 & n1741 ) | ( n1736 & n1741 ) ;
  assign n1743 = ( n1688 & n1736 ) | ( n1688 & n1741 ) | ( n1736 & n1741 ) ;
  assign n1744 = ( n1688 & n1742 ) | ( n1688 & ~n1743 ) | ( n1742 & ~n1743 ) ;
  assign n1745 = x191 & ~n350 ;
  assign n1746 = ( n1016 & n1028 ) | ( n1016 & n1745 ) | ( n1028 & n1745 ) ;
  assign n1747 = ( n1016 & n1745 ) | ( n1016 & ~n1746 ) | ( n1745 & ~n1746 ) ;
  assign n1748 = ( n1028 & ~n1746 ) | ( n1028 & n1747 ) | ( ~n1746 & n1747 ) ;
  assign n1749 = ( n335 & n347 ) | ( n335 & n1748 ) | ( n347 & n1748 ) ;
  assign n1750 = ( n335 & n1748 ) | ( n335 & ~n1749 ) | ( n1748 & ~n1749 ) ;
  assign n1751 = ( n347 & ~n1749 ) | ( n347 & n1750 ) | ( ~n1749 & n1750 ) ;
  assign n1752 = ~n341 & n1751 ;
  assign n1753 = n341 & ~n1751 ;
  assign n1754 = n1752 | n1753 ;
  assign n1755 = ~n329 & n966 ;
  assign n1756 = ( x205 & n1754 ) | ( x205 & ~n1755 ) | ( n1754 & ~n1755 ) ;
  assign n1757 = ( ~n352 & n1023 ) | ( ~n352 & n1031 ) | ( n1023 & n1031 ) ;
  assign n1758 = ( n352 & ~n1031 ) | ( n352 & n1757 ) | ( ~n1031 & n1757 ) ;
  assign n1759 = ( ~n1023 & n1757 ) | ( ~n1023 & n1758 ) | ( n1757 & n1758 ) ;
  assign n1760 = ( n335 & n347 ) | ( n335 & n1759 ) | ( n347 & n1759 ) ;
  assign n1761 = ( n335 & n1759 ) | ( n335 & ~n1760 ) | ( n1759 & ~n1760 ) ;
  assign n1762 = ( n347 & ~n1760 ) | ( n347 & n1761 ) | ( ~n1760 & n1761 ) ;
  assign n1763 = ~n341 & n1762 ;
  assign n1764 = n341 & ~n1762 ;
  assign n1765 = n1763 | n1764 ;
  assign n1766 = ( x205 & n1755 ) | ( x205 & n1765 ) | ( n1755 & n1765 ) ;
  assign n1767 = n1756 & n1766 ;
  assign n1768 = ( n983 & n989 ) | ( n983 & ~n991 ) | ( n989 & ~n991 ) ;
  assign n1769 = ~n983 & n988 ;
  assign n1770 = ( n310 & ~n983 ) | ( n310 & n1769 ) | ( ~n983 & n1769 ) ;
  assign n1771 = ( n310 & n983 ) | ( n310 & n1769 ) | ( n983 & n1769 ) ;
  assign n1772 = ( n983 & n1770 ) | ( n983 & ~n1771 ) | ( n1770 & ~n1771 ) ;
  assign n1773 = ( n1001 & n1768 ) | ( n1001 & ~n1772 ) | ( n1768 & ~n1772 ) ;
  assign n1774 = ( ~n1768 & n1772 ) | ( ~n1768 & n1773 ) | ( n1772 & n1773 ) ;
  assign n1775 = ( ~n1001 & n1773 ) | ( ~n1001 & n1774 ) | ( n1773 & n1774 ) ;
  assign n1776 = ~n230 & n1775 ;
  assign n1777 = n230 & ~n1775 ;
  assign n1778 = n1776 | n1777 ;
  assign n1779 = ( n296 & n308 ) | ( n296 & ~n1778 ) | ( n308 & ~n1778 ) ;
  assign n1780 = ( ~n296 & n1778 ) | ( ~n296 & n1779 ) | ( n1778 & n1779 ) ;
  assign n1781 = ( ~n308 & n1779 ) | ( ~n308 & n1780 ) | ( n1779 & n1780 ) ;
  assign n1782 = n302 | n1781 ;
  assign n1783 = n302 & n1781 ;
  assign n1784 = n1782 & ~n1783 ;
  assign n1785 = ( x205 & ~n323 ) | ( x205 & n1784 ) | ( ~n323 & n1784 ) ;
  assign n1786 = n323 | n1785 ;
  assign n1787 = ( ~n1784 & n1785 ) | ( ~n1784 & n1786 ) | ( n1785 & n1786 ) ;
  assign n1788 = ~x5 & x186 ;
  assign n1789 = ~n227 & n1788 ;
  assign n1790 = n302 & ~n1001 ;
  assign n1791 = ( n230 & ~n1001 ) | ( n230 & n1790 ) | ( ~n1001 & n1790 ) ;
  assign n1792 = n230 | n308 ;
  assign n1793 = n302 & ~n983 ;
  assign n1794 = ( ~n983 & n1792 ) | ( ~n983 & n1793 ) | ( n1792 & n1793 ) ;
  assign n1795 = ~n988 & n1794 ;
  assign n1796 = ( n1789 & n1791 ) | ( n1789 & ~n1795 ) | ( n1791 & ~n1795 ) ;
  assign n1797 = ( ~n1791 & n1795 ) | ( ~n1791 & n1796 ) | ( n1795 & n1796 ) ;
  assign n1798 = ( ~n1789 & n1796 ) | ( ~n1789 & n1797 ) | ( n1796 & n1797 ) ;
  assign n1799 = ( ~n302 & n323 ) | ( ~n302 & n1792 ) | ( n323 & n1792 ) ;
  assign n1800 = ~n323 & n983 ;
  assign n1801 = ( n302 & n1799 ) | ( n302 & ~n1800 ) | ( n1799 & ~n1800 ) ;
  assign n1802 = ~n989 & n1801 ;
  assign n1803 = ( ~n230 & n1798 ) | ( ~n230 & n1802 ) | ( n1798 & n1802 ) ;
  assign n1804 = ( n1798 & n1802 ) | ( n1798 & ~n1803 ) | ( n1802 & ~n1803 ) ;
  assign n1805 = ( n230 & n1803 ) | ( n230 & ~n1804 ) | ( n1803 & ~n1804 ) ;
  assign n1806 = ( n296 & n308 ) | ( n296 & ~n1805 ) | ( n308 & ~n1805 ) ;
  assign n1807 = ( ~n296 & n1805 ) | ( ~n296 & n1806 ) | ( n1805 & n1806 ) ;
  assign n1808 = ( ~n308 & n1806 ) | ( ~n308 & n1807 ) | ( n1806 & n1807 ) ;
  assign n1809 = n302 | n1808 ;
  assign n1810 = n302 & n1808 ;
  assign n1811 = n1809 & ~n1810 ;
  assign n1812 = ( x205 & n323 ) | ( x205 & n1811 ) | ( n323 & n1811 ) ;
  assign n1813 = ~n323 & n1812 ;
  assign n1814 = ( ~n1811 & n1812 ) | ( ~n1811 & n1813 ) | ( n1812 & n1813 ) ;
  assign n1815 = n1787 & ~n1814 ;
  assign n1816 = n1767 & ~n1815 ;
  assign n1817 = ( x205 & n329 ) | ( x205 & ~n1765 ) | ( n329 & ~n1765 ) ;
  assign n1818 = ( ~x205 & n329 ) | ( ~x205 & n1754 ) | ( n329 & n1754 ) ;
  assign n1819 = ~n1817 & n1818 ;
  assign n1820 = n1815 | n1819 ;
  assign n1821 = ( n1767 & n1815 ) | ( n1767 & n1819 ) | ( n1815 & n1819 ) ;
  assign n1822 = ( n1816 & n1820 ) | ( n1816 & ~n1821 ) | ( n1820 & ~n1821 ) ;
  assign y0 = x164 ;
  assign y1 = x0 ;
  assign y2 = x0 ;
  assign y3 = x167 ;
  assign y4 = x169 ;
  assign y5 = x170 ;
  assign y6 = x171 ;
  assign y7 = x172 ;
  assign y8 = x173 ;
  assign y9 = x175 ;
  assign y10 = x177 ;
  assign y11 = x178 ;
  assign y12 = x179 ;
  assign y13 = x180 ;
  assign y14 = x181 ;
  assign y15 = x182 ;
  assign y16 = x183 ;
  assign y17 = x184 ;
  assign y18 = x185 ;
  assign y19 = x186 ;
  assign y20 = x187 ;
  assign y21 = x188 ;
  assign y22 = x189 ;
  assign y23 = x190 ;
  assign y24 = x191 ;
  assign y25 = x192 ;
  assign y26 = x193 ;
  assign y27 = x194 ;
  assign y28 = x195 ;
  assign y29 = x197 ;
  assign y30 = x198 ;
  assign y31 = x199 ;
  assign y32 = x200 ;
  assign y33 = x201 ;
  assign y34 = x202 ;
  assign y35 = x203 ;
  assign y36 = x204 ;
  assign y37 = ~x4 ;
  assign y38 = x168 ;
  assign y39 = x176 ;
  assign y40 = x196 ;
  assign y41 = n208 ;
  assign y42 = ~n211 ;
  assign y43 = ~n214 ;
  assign y44 = ~n217 ;
  assign y45 = ~n220 ;
  assign y46 = x0 ;
  assign y47 = x53 ;
  assign y48 = ~n221 ;
  assign y49 = ~x4 ;
  assign y50 = ~n221 ;
  assign y51 = ~n223 ;
  assign y52 = ~x4 ;
  assign y53 = ~n223 ;
  assign y54 = x0 ;
  assign y55 = n224 ;
  assign y56 = ~n233 ;
  assign y57 = ~n553 ;
  assign y58 = n950 ;
  assign y59 = n950 ;
  assign y60 = ~n982 ;
  assign y61 = ~n995 ;
  assign y62 = ~n1000 ;
  assign y63 = ~n1007 ;
  assign y64 = ~n1012 ;
  assign y65 = ~n1027 ;
  assign y66 = ~n1035 ;
  assign y67 = ~n1039 ;
  assign y68 = ~n1042 ;
  assign y69 = ~n1132 ;
  assign y70 = ~n1230 ;
  assign y71 = ~n1316 ;
  assign y72 = n1324 ;
  assign y73 = ~n1329 ;
  assign y74 = ~n1335 ;
  assign y75 = n1343 ;
  assign y76 = ~n1353 ;
  assign y77 = n1365 ;
  assign y78 = ~n1370 ;
  assign y79 = ~n1376 ;
  assign y80 = ~n1380 ;
  assign y81 = ~n1393 ;
  assign y82 = ~n1398 ;
  assign y83 = ~n1404 ;
  assign y84 = ~n1408 ;
  assign y85 = ~n1414 ;
  assign y86 = ~n1419 ;
  assign y87 = ~n1433 ;
  assign y88 = ~n1440 ;
  assign y89 = ~n1444 ;
  assign y90 = ~n1447 ;
  assign y91 = ~n1452 ;
  assign y92 = n1456 ;
  assign y93 = n1456 ;
  assign y94 = n1459 ;
  assign y95 = n1459 ;
  assign y96 = ~n1472 ;
  assign y97 = ~n1477 ;
  assign y98 = ~n1483 ;
  assign y99 = ~n1487 ;
  assign y100 = ~n1502 ;
  assign y101 = ~n1510 ;
  assign y102 = ~n1514 ;
  assign y103 = ~n1517 ;
  assign y104 = ~n1597 ;
  assign y105 = n1664 ;
  assign y106 = n1744 ;
  assign y107 = n1822 ;
endmodule
