module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, y0, y1, y2, y3, y4, y5, y6);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10;
  output y0, y1, y2, y3, y4, y5, y6;
  wire n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212;
  assign n40 = x7 ^ x6;
  assign n41 = x8 & x9;
  assign n42 = x7 & n41;
  assign n43 = ~n40 & n42;
  assign n44 = n43 ^ n40;
  assign n30 = x5 ^ x4;
  assign n13 = x3 ^ x2;
  assign n14 = n13 ^ x6;
  assign n15 = n14 ^ n13;
  assign n16 = x1 & x4;
  assign n17 = n16 ^ x0;
  assign n18 = n17 ^ x5;
  assign n19 = n18 ^ n17;
  assign n20 = x2 ^ x1;
  assign n21 = n20 ^ n17;
  assign n22 = n19 & n21;
  assign n23 = n22 ^ n17;
  assign n24 = n23 ^ n13;
  assign n25 = ~n15 & n24;
  assign n26 = n25 ^ n13;
  assign n12 = x4 ^ x3;
  assign n27 = n26 ^ n12;
  assign n28 = x7 & n27;
  assign n29 = n28 ^ n26;
  assign n31 = n30 ^ n29;
  assign n32 = ~x8 & n31;
  assign n33 = n32 ^ n30;
  assign n34 = n33 ^ x9;
  assign n35 = n34 ^ n33;
  assign n36 = x6 ^ x5;
  assign n37 = n36 ^ n33;
  assign n38 = n35 & n37;
  assign n39 = n38 ^ n33;
  assign n45 = n44 ^ n39;
  assign n46 = x10 & n45;
  assign n47 = n46 ^ n39;
  assign n48 = ~x7 & ~x8;
  assign n55 = x1 & x2;
  assign n56 = n55 ^ x3;
  assign n52 = ~x0 & n16;
  assign n53 = n52 ^ x1;
  assign n51 = x2 & x4;
  assign n54 = n53 ^ n51;
  assign n57 = n56 ^ n54;
  assign n58 = x5 & n57;
  assign n59 = n58 ^ n54;
  assign n49 = x2 & x3;
  assign n50 = n49 ^ x4;
  assign n60 = n59 ^ n50;
  assign n61 = n60 ^ n59;
  assign n62 = n59 ^ x9;
  assign n63 = n62 ^ n59;
  assign n64 = ~n61 & ~n63;
  assign n65 = n64 ^ n59;
  assign n66 = x6 & ~n65;
  assign n67 = n66 ^ n59;
  assign n68 = n48 & ~n67;
  assign n71 = x4 & x5;
  assign n72 = n71 ^ x6;
  assign n73 = n72 ^ x8;
  assign n74 = n73 ^ n72;
  assign n75 = n74 ^ x9;
  assign n76 = x3 & x4;
  assign n77 = n76 ^ x5;
  assign n78 = n77 ^ x7;
  assign n79 = x7 & ~n78;
  assign n80 = n79 ^ n72;
  assign n81 = n80 ^ x7;
  assign n82 = n75 & ~n81;
  assign n83 = n82 ^ n79;
  assign n84 = n83 ^ x7;
  assign n69 = x5 & x6;
  assign n70 = n69 ^ x7;
  assign n85 = n84 ^ n70;
  assign n86 = ~x9 & ~n85;
  assign n87 = n86 ^ n70;
  assign n88 = ~x10 & n87;
  assign n89 = ~n68 & n88;
  assign n90 = x6 & x7;
  assign n91 = x8 & n90;
  assign n92 = ~x9 & n91;
  assign n93 = ~x8 & ~n90;
  assign n94 = x10 & ~n93;
  assign n95 = ~n92 & n94;
  assign n96 = ~n89 & ~n95;
  assign n97 = n91 ^ x10;
  assign n98 = n97 ^ n91;
  assign n99 = x5 & n90;
  assign n100 = n99 ^ x8;
  assign n101 = n100 ^ n91;
  assign n102 = ~n98 & ~n101;
  assign n103 = n102 ^ n91;
  assign n104 = n103 ^ x9;
  assign n105 = n104 ^ x10;
  assign n106 = n105 ^ n103;
  assign n107 = n103 ^ x10;
  assign n108 = n107 ^ n103;
  assign n109 = x6 & n71;
  assign n110 = n49 & n109;
  assign n111 = ~x7 & ~n110;
  assign n112 = x5 ^ x2;
  assign n114 = n112 ^ x2;
  assign n115 = n114 ^ n112;
  assign n116 = n115 ^ x6;
  assign n117 = n114 ^ x4;
  assign n118 = n117 ^ n114;
  assign n119 = n118 ^ n116;
  assign n120 = ~n116 & ~n119;
  assign n113 = n112 ^ x6;
  assign n121 = n120 ^ n113;
  assign n122 = n121 ^ n116;
  assign n123 = x6 ^ x3;
  assign n124 = n120 ^ n116;
  assign n125 = ~n123 & ~n124;
  assign n126 = n125 ^ x6;
  assign n127 = ~n122 & ~n126;
  assign n128 = n127 ^ x6;
  assign n129 = n128 ^ x5;
  assign n130 = n129 ^ x6;
  assign n131 = n111 & n130;
  assign n132 = ~x0 & ~x5;
  assign n133 = x1 & ~n132;
  assign n134 = ~x3 & x5;
  assign n135 = n133 & ~n134;
  assign n138 = n36 ^ x6;
  assign n139 = n36 ^ x3;
  assign n140 = n139 ^ n36;
  assign n141 = ~n138 & ~n140;
  assign n142 = n141 ^ n36;
  assign n143 = x4 & n142;
  assign n144 = n143 ^ n36;
  assign n136 = x3 & ~x6;
  assign n137 = n51 & n136;
  assign n145 = n144 ^ n137;
  assign n146 = n135 & n145;
  assign n147 = n146 ^ n144;
  assign n148 = n131 & ~n147;
  assign n149 = ~x3 & n90;
  assign n150 = ~n148 & ~n149;
  assign n151 = ~x8 & ~n150;
  assign n152 = x7 & ~n109;
  assign n153 = ~n93 & n152;
  assign n154 = n71 ^ n40;
  assign n155 = x8 ^ x7;
  assign n156 = n155 ^ x8;
  assign n157 = x8 ^ x3;
  assign n158 = n156 & n157;
  assign n159 = n158 ^ x8;
  assign n160 = n159 ^ n40;
  assign n161 = n154 & n160;
  assign n162 = n161 ^ n158;
  assign n163 = n162 ^ x8;
  assign n164 = n163 ^ n71;
  assign n165 = n40 & n164;
  assign n166 = n165 ^ n40;
  assign n167 = ~n153 & ~n166;
  assign n168 = ~n151 & n167;
  assign n169 = n168 ^ n103;
  assign n170 = n169 ^ n103;
  assign n171 = ~n108 & ~n170;
  assign n172 = n171 ^ n103;
  assign n173 = ~n106 & n172;
  assign n174 = n173 ^ n104;
  assign n175 = ~x5 & ~x6;
  assign n176 = n48 & n175;
  assign n177 = ~x4 & n176;
  assign n178 = ~x2 & n71;
  assign n179 = n91 & n178;
  assign n180 = ~n177 & ~n179;
  assign n181 = ~x9 & ~x10;
  assign n182 = ~x3 & n181;
  assign n183 = ~n180 & n182;
  assign n184 = n133 & n175;
  assign n185 = n49 & n184;
  assign n186 = n55 & n76;
  assign n187 = x4 & n175;
  assign n188 = n187 ^ x6;
  assign n189 = ~n186 & ~n188;
  assign n190 = ~n185 & ~n189;
  assign n191 = n111 & n190;
  assign n192 = ~x8 & ~n191;
  assign n193 = ~x2 & ~x3;
  assign n194 = n71 & ~n193;
  assign n195 = n90 & n194;
  assign n196 = ~x9 & ~n195;
  assign n197 = ~n192 & n196;
  assign n198 = x9 ^ x8;
  assign n199 = ~x9 & ~n76;
  assign n200 = ~n198 & n199;
  assign n201 = n200 ^ n198;
  assign n202 = n99 & ~n201;
  assign n203 = ~x10 & ~n202;
  assign n204 = ~n197 & n203;
  assign n205 = n135 & n137;
  assign n206 = n175 & ~n205;
  assign n207 = n48 & ~n110;
  assign n208 = ~n206 & n207;
  assign n209 = x8 & n195;
  assign n210 = n181 & ~n209;
  assign n211 = ~n208 & n210;
  assign n212 = n181 & n207;
  assign y0 = n47;
  assign y1 = ~n96;
  assign y2 = n174;
  assign y3 = ~n183;
  assign y4 = ~n204;
  assign y5 = ~n211;
  assign y6 = ~n212;
endmodule
