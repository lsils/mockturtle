module top( in_0_ , in_1_ , in_2_ , in_3_ , in_4_ , in_5_ , in_6_ , in_7_ , in_8_ , in_9_ , in_10_ , in_11_ , in_12_ , in_13_ , in_14_ , in_15_ , out_0_ , out_1_ , out_2_ , out_3_ , out_4_ );
  input in_0_ , in_1_ , in_2_ , in_3_ , in_4_ , in_5_ , in_6_ , in_7_ , in_8_ , in_9_ , in_10_ , in_11_ , in_12_ , in_13_ , in_14_ , in_15_ ;
  output out_0_ , out_1_ , out_2_ , out_3_ , out_4_ ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 ;
  assign n17 = in_14_ & in_15_ ;
  assign n18 = in_12_ | in_13_ ;
  assign n19 = in_4_ | in_5_ ;
  assign n20 = in_0_ | in_1_ ;
  assign n21 = in_2_ & in_3_ ;
  assign n22 = ( n19 & n20 ) | ( n19 & n21 ) | ( n20 & n21 ) ;
  assign n23 = ( ~n19 & n20 ) | ( ~n19 & n21 ) | ( n20 & n21 ) ;
  assign n24 = ( n19 & ~n22 ) | ( n19 & n23 ) | ( ~n22 & n23 ) ;
  assign n25 = in_10_ & in_11_ ;
  assign n26 = in_6_ & in_7_ ;
  assign n27 = in_8_ | in_9_ ;
  assign n28 = ( n25 & n26 ) | ( n25 & n27 ) | ( n26 & n27 ) ;
  assign n29 = ( ~n25 & n26 ) | ( ~n25 & n27 ) | ( n26 & n27 ) ;
  assign n30 = ( n25 & ~n28 ) | ( n25 & n29 ) | ( ~n28 & n29 ) ;
  assign n31 = ( n18 & n24 ) | ( n18 & n30 ) | ( n24 & n30 ) ;
  assign n32 = ( ~n18 & n24 ) | ( ~n18 & n30 ) | ( n24 & n30 ) ;
  assign n33 = ( n18 & ~n31 ) | ( n18 & n32 ) | ( ~n31 & n32 ) ;
  assign n34 = n17 & n33 ;
  assign n35 = n17 | n33 ;
  assign n36 = ~n34 & n35 ;
  assign n37 = ( n22 & n28 ) | ( n22 & n31 ) | ( n28 & n31 ) ;
  assign n38 = ( n22 & n28 ) | ( n22 & ~n31 ) | ( n28 & ~n31 ) ;
  assign n39 = ( n31 & ~n37 ) | ( n31 & n38 ) | ( ~n37 & n38 ) ;
  assign n40 = n34 & n39 ;
  assign n41 = n34 | n39 ;
  assign n42 = ~n40 & n41 ;
  assign n43 = n37 & n40 ;
  assign n44 = n37 | n40 ;
  assign n45 = ~n43 & n44 ;
  assign out_0_ = 1'b0 ;
  assign out_1_ = n36 ;
  assign out_2_ = n42 ;
  assign out_3_ = n45 ;
  assign out_4_ = n43 ;
endmodule
