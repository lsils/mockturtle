module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 ;
  wire n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 ;
  assign n13 = x2 | x3 ;
  assign n14 = x6 & x7 ;
  assign n15 = ~x5 & n14 ;
  assign n16 = x4 & n15 ;
  assign n17 = ~x1 & n16 ;
  assign n18 = ~n13 & n17 ;
  assign n9 = x4 & x5 ;
  assign n10 = x1 | x3 ;
  assign n11 = ( x2 & ~n9 ) | ( x2 & n10 ) | ( ~n9 & n10 ) ;
  assign n12 = n9 | n11 ;
  assign n19 = ~x0 & n12 ;
  assign n20 = ( ~x0 & n18 ) | ( ~x0 & n19 ) | ( n18 & n19 ) ;
  assign n25 = ~x6 & x7 ;
  assign n26 = x2 & x5 ;
  assign n27 = ( x4 & n25 ) | ( x4 & n26 ) | ( n25 & n26 ) ;
  assign n28 = ~x4 & n27 ;
  assign n21 = x6 & ~x7 ;
  assign n22 = ~x5 & n21 ;
  assign n23 = ( x2 & x4 ) | ( x2 & n22 ) | ( x4 & n22 ) ;
  assign n24 = ~x2 & n23 ;
  assign n29 = ~x3 & n24 ;
  assign n30 = ( ~x3 & n28 ) | ( ~x3 & n29 ) | ( n28 & n29 ) ;
  assign n43 = ( ~x0 & x1 ) | ( ~x0 & n30 ) | ( x1 & n30 ) ;
  assign n36 = ( ~x1 & x3 ) | ( ~x1 & x4 ) | ( x3 & x4 ) ;
  assign n37 = x2 & ~n36 ;
  assign n38 = ( x1 & ~x2 ) | ( x1 & n36 ) | ( ~x2 & n36 ) ;
  assign n39 = ( ~x1 & n37 ) | ( ~x1 & n38 ) | ( n37 & n38 ) ;
  assign n31 = ( x2 & x4 ) | ( x2 & ~x5 ) | ( x4 & ~x5 ) ;
  assign n32 = ( x2 & ~x6 ) | ( x2 & n31 ) | ( ~x6 & n31 ) ;
  assign n33 = x2 & ~n32 ;
  assign n34 = n32 | n33 ;
  assign n35 = ( ~x2 & n33 ) | ( ~x2 & n34 ) | ( n33 & n34 ) ;
  assign n40 = ( x1 & ~n35 ) | ( x1 & n39 ) | ( ~n35 & n39 ) ;
  assign n41 = ~x3 & n40 ;
  assign n42 = ( x3 & n39 ) | ( x3 & n41 ) | ( n39 & n41 ) ;
  assign n44 = x0 | n42 ;
  assign n45 = ( x1 & ~n43 ) | ( x1 & n44 ) | ( ~n43 & n44 ) ;
  assign n65 = x3 | x5 ;
  assign n66 = x3 & x4 ;
  assign n67 = x4 & ~x5 ;
  assign n68 = ( n65 & ~n66 ) | ( n65 & n67 ) | ( ~n66 & n67 ) ;
  assign n69 = x2 & ~n68 ;
  assign n70 = ( x1 & ~n68 ) | ( x1 & n69 ) | ( ~n68 & n69 ) ;
  assign n75 = ( ~x1 & x3 ) | ( ~x1 & x5 ) | ( x3 & x5 ) ;
  assign n76 = ( x4 & x5 ) | ( x4 & ~n75 ) | ( x5 & ~n75 ) ;
  assign n77 = ( ~x3 & x4 ) | ( ~x3 & n75 ) | ( x4 & n75 ) ;
  assign n78 = n76 & ~n77 ;
  assign n71 = ~x3 & x5 ;
  assign n72 = ~x4 & n71 ;
  assign n73 = ~x1 & n72 ;
  assign n74 = ~x2 & n73 ;
  assign n79 = ( x3 & x4 ) | ( x3 & ~n36 ) | ( x4 & ~n36 ) ;
  assign n80 = x2 & n36 ;
  assign n81 = ( x1 & n36 ) | ( x1 & n80 ) | ( n36 & n80 ) ;
  assign n82 = n79 & ~n81 ;
  assign n83 = n74 | n82 ;
  assign n84 = ( ~n70 & n78 ) | ( ~n70 & n83 ) | ( n78 & n83 ) ;
  assign n85 = n70 | n84 ;
  assign n46 = ( x2 & x3 ) | ( x2 & ~x5 ) | ( x3 & ~x5 ) ;
  assign n47 = ( x2 & x4 ) | ( x2 & ~n46 ) | ( x4 & ~n46 ) ;
  assign n48 = ( ~x3 & x5 ) | ( ~x3 & n47 ) | ( x5 & n47 ) ;
  assign n49 = n46 | n48 ;
  assign n50 = ( ~n47 & n48 ) | ( ~n47 & n49 ) | ( n48 & n49 ) ;
  assign n54 = ( ~x1 & x6 ) | ( ~x1 & n50 ) | ( x6 & n50 ) ;
  assign n51 = x5 | x6 ;
  assign n52 = x4 & ~n13 ;
  assign n53 = ~n51 & n52 ;
  assign n55 = ~x1 & n53 ;
  assign n56 = ( ~n50 & n54 ) | ( ~n50 & n55 ) | ( n54 & n55 ) ;
  assign n57 = ( x2 & x5 ) | ( x2 & x6 ) | ( x5 & x6 ) ;
  assign n58 = ( ~x4 & x6 ) | ( ~x4 & n57 ) | ( x6 & n57 ) ;
  assign n59 = x6 & ~n58 ;
  assign n60 = n58 | n59 ;
  assign n61 = ( ~x6 & n59 ) | ( ~x6 & n60 ) | ( n59 & n60 ) ;
  assign n62 = x1 | x7 ;
  assign n63 = ( x3 & n61 ) | ( x3 & n62 ) | ( n61 & n62 ) ;
  assign n64 = n61 & ~n63 ;
  assign n86 = ( ~x0 & n56 ) | ( ~x0 & n64 ) | ( n56 & n64 ) ;
  assign n87 = ~n85 & n86 ;
  assign n88 = ( ~x0 & n85 ) | ( ~x0 & n87 ) | ( n85 & n87 ) ;
  assign n111 = ( x3 & x5 ) | ( x3 & x6 ) | ( x5 & x6 ) ;
  assign n112 = x3 & n111 ;
  assign n113 = ( x2 & ~x3 ) | ( x2 & n111 ) | ( ~x3 & n111 ) ;
  assign n114 = ~n111 & n113 ;
  assign n115 = n112 | n114 ;
  assign n134 = ~x1 & n115 ;
  assign n116 = x2 | n51 ;
  assign n117 = ( ~x1 & x3 ) | ( ~x1 & n116 ) | ( x3 & n116 ) ;
  assign n118 = x1 | n117 ;
  assign n122 = ( x2 & ~x3 ) | ( x2 & x5 ) | ( ~x3 & x5 ) ;
  assign n123 = ( x2 & x3 ) | ( x2 & ~x6 ) | ( x3 & ~x6 ) ;
  assign n124 = n122 | n123 ;
  assign n125 = ( x3 & ~x5 ) | ( x3 & n124 ) | ( ~x5 & n124 ) ;
  assign n126 = x4 | n125 ;
  assign n120 = ~x2 & x3 ;
  assign n121 = x5 & x6 ;
  assign n127 = n120 & n121 ;
  assign n128 = x4 & ~n127 ;
  assign n129 = n126 & ~n128 ;
  assign n130 = x1 | n129 ;
  assign n119 = x4 | n51 ;
  assign n131 = ~n119 & n120 ;
  assign n132 = x1 & ~n131 ;
  assign n133 = n130 & ~n132 ;
  assign n135 = n118 & ~n133 ;
  assign n136 = ( ~n115 & n134 ) | ( ~n115 & n135 ) | ( n134 & n135 ) ;
  assign n89 = ( x1 & x2 ) | ( x1 & x4 ) | ( x2 & x4 ) ;
  assign n90 = ( x3 & x6 ) | ( x3 & n89 ) | ( x6 & n89 ) ;
  assign n91 = ( x5 & ~x6 ) | ( x5 & n90 ) | ( ~x6 & n90 ) ;
  assign n92 = ( x3 & x5 ) | ( x3 & ~n90 ) | ( x5 & ~n90 ) ;
  assign n93 = n91 & ~n92 ;
  assign n94 = ~x2 & x4 ;
  assign n95 = x3 & n94 ;
  assign n96 = x5 & n25 ;
  assign n97 = n95 & n96 ;
  assign n98 = ( ~x4 & x6 ) | ( ~x4 & x7 ) | ( x6 & x7 ) ;
  assign n99 = ( x2 & ~x6 ) | ( x2 & n98 ) | ( ~x6 & n98 ) ;
  assign n100 = ( ~x4 & x7 ) | ( ~x4 & n99 ) | ( x7 & n99 ) ;
  assign n101 = ~n98 & n100 ;
  assign n102 = ( ~n99 & n100 ) | ( ~n99 & n101 ) | ( n100 & n101 ) ;
  assign n103 = ( x3 & ~x5 ) | ( x3 & n102 ) | ( ~x5 & n102 ) ;
  assign n104 = ( n29 & n102 ) | ( n29 & ~n103 ) | ( n102 & ~n103 ) ;
  assign n105 = x1 & ~n13 ;
  assign n106 = ( ~n9 & n25 ) | ( ~n9 & n105 ) | ( n25 & n105 ) ;
  assign n107 = n9 & n106 ;
  assign n108 = ( ~n97 & n104 ) | ( ~n97 & n107 ) | ( n104 & n107 ) ;
  assign n109 = x1 & ~n107 ;
  assign n110 = ( n97 & n108 ) | ( n97 & ~n109 ) | ( n108 & ~n109 ) ;
  assign n137 = ( ~x0 & n93 ) | ( ~x0 & n110 ) | ( n93 & n110 ) ;
  assign n138 = n136 & n137 ;
  assign n139 = ( x0 & n136 ) | ( x0 & ~n138 ) | ( n136 & ~n138 ) ;
  assign n191 = x3 & x5 ;
  assign n192 = x5 & ~x7 ;
  assign n193 = ( x1 & n191 ) | ( x1 & n192 ) | ( n191 & n192 ) ;
  assign n194 = ( ~x1 & x7 ) | ( ~x1 & n193 ) | ( x7 & n193 ) ;
  assign n195 = ( ~x5 & n191 ) | ( ~x5 & n194 ) | ( n191 & n194 ) ;
  assign n196 = ( ~n191 & n193 ) | ( ~n191 & n195 ) | ( n193 & n195 ) ;
  assign n197 = ~x3 & n21 ;
  assign n198 = ( x1 & ~x5 ) | ( x1 & n197 ) | ( ~x5 & n197 ) ;
  assign n199 = ~x1 & n198 ;
  assign n200 = x6 & ~n199 ;
  assign n201 = ( n196 & n199 ) | ( n196 & ~n200 ) | ( n199 & ~n200 ) ;
  assign n202 = x4 & ~n201 ;
  assign n186 = ( x3 & x6 ) | ( x3 & x7 ) | ( x6 & x7 ) ;
  assign n187 = ( ~x3 & x5 ) | ( ~x3 & n186 ) | ( x5 & n186 ) ;
  assign n188 = ( x6 & x7 ) | ( x6 & n187 ) | ( x7 & n187 ) ;
  assign n189 = ~n186 & n188 ;
  assign n190 = ( ~n187 & n188 ) | ( ~n187 & n189 ) | ( n188 & n189 ) ;
  assign n203 = ~x1 & n190 ;
  assign n204 = x4 | n203 ;
  assign n205 = ~n202 & n204 ;
  assign n206 = x2 | n205 ;
  assign n178 = ( x5 & ~x6 ) | ( x5 & x7 ) | ( ~x6 & x7 ) ;
  assign n179 = ~x7 & n178 ;
  assign n180 = ( x4 & ~x5 ) | ( x4 & n179 ) | ( ~x5 & n179 ) ;
  assign n181 = ( n178 & n179 ) | ( n178 & n180 ) | ( n179 & n180 ) ;
  assign n182 = x3 | n181 ;
  assign n183 = ~x4 & n15 ;
  assign n184 = x3 & ~n183 ;
  assign n185 = n182 & ~n184 ;
  assign n207 = ~x1 & n185 ;
  assign n208 = x2 & ~n207 ;
  assign n209 = n206 & ~n208 ;
  assign n140 = ( ~x1 & x2 ) | ( ~x1 & n13 ) | ( x2 & n13 ) ;
  assign n141 = ( x1 & x2 ) | ( x1 & ~n13 ) | ( x2 & ~n13 ) ;
  assign n142 = ( ~x2 & n140 ) | ( ~x2 & n141 ) | ( n140 & n141 ) ;
  assign n143 = ( x5 & x6 ) | ( x5 & n142 ) | ( x6 & n142 ) ;
  assign n144 = ( x4 & ~x6 ) | ( x4 & n143 ) | ( ~x6 & n143 ) ;
  assign n145 = ( x4 & x5 ) | ( x4 & ~n143 ) | ( x5 & ~n143 ) ;
  assign n146 = n144 & ~n145 ;
  assign n154 = ~x1 & x2 ;
  assign n155 = ~x1 & x4 ;
  assign n156 = ( n94 & n154 ) | ( n94 & ~n155 ) | ( n154 & ~n155 ) ;
  assign n157 = ( ~x3 & x6 ) | ( ~x3 & n156 ) | ( x6 & n156 ) ;
  assign n158 = ( x5 & ~x6 ) | ( x5 & n157 ) | ( ~x6 & n157 ) ;
  assign n159 = ( x3 & ~x5 ) | ( x3 & n157 ) | ( ~x5 & n157 ) ;
  assign n160 = n158 & n159 ;
  assign n147 = x1 & ~x2 ;
  assign n148 = x1 | n13 ;
  assign n149 = ( ~x1 & n147 ) | ( ~x1 & n148 ) | ( n147 & n148 ) ;
  assign n150 = ( x4 & ~x6 ) | ( x4 & n149 ) | ( ~x6 & n149 ) ;
  assign n151 = ( ~x5 & x6 ) | ( ~x5 & n150 ) | ( x6 & n150 ) ;
  assign n152 = ( ~x4 & x5 ) | ( ~x4 & n150 ) | ( x5 & n150 ) ;
  assign n153 = n151 | n152 ;
  assign n166 = x4 | x6 ;
  assign n167 = ( ~x2 & x4 ) | ( ~x2 & x6 ) | ( x4 & x6 ) ;
  assign n168 = ( x3 & x4 ) | ( x3 & n167 ) | ( x4 & n167 ) ;
  assign n169 = n167 & n168 ;
  assign n170 = n166 & ~n169 ;
  assign n171 = x1 & ~n170 ;
  assign n161 = x3 & ~x6 ;
  assign n162 = x4 & ~x6 ;
  assign n163 = ( ~x5 & x6 ) | ( ~x5 & n162 ) | ( x6 & n162 ) ;
  assign n164 = ( x3 & ~x5 ) | ( x3 & n162 ) | ( ~x5 & n162 ) ;
  assign n165 = ( n161 & n163 ) | ( n161 & ~n164 ) | ( n163 & ~n164 ) ;
  assign n172 = x2 & n165 ;
  assign n173 = x1 | n172 ;
  assign n174 = ~n171 & n173 ;
  assign n175 = n153 & ~n174 ;
  assign n176 = ( n146 & ~n160 ) | ( n146 & n175 ) | ( ~n160 & n175 ) ;
  assign n177 = ~n146 & n176 ;
  assign n210 = x0 | n177 ;
  assign n211 = ( x0 & ~n209 ) | ( x0 & n210 ) | ( ~n209 & n210 ) ;
  assign n212 = ( ~x0 & x2 ) | ( ~x0 & n10 ) | ( x2 & n10 ) ;
  assign n213 = x0 | n212 ;
  assign n214 = x5 | n213 ;
  assign n215 = ( ~x4 & x6 ) | ( ~x4 & n214 ) | ( x6 & n214 ) ;
  assign n216 = x4 | n215 ;
  assign n217 = x7 | n216 ;
  assign n218 = x5 & ~x6 ;
  assign n219 = ~x7 & n218 ;
  assign n220 = x5 | n219 ;
  assign n221 = x3 | x4 ;
  assign n222 = ( ~n219 & n220 ) | ( ~n219 & n221 ) | ( n220 & n221 ) ;
  assign n223 = x1 | n222 ;
  assign n224 = ( ~x0 & x2 ) | ( ~x0 & n223 ) | ( x2 & n223 ) ;
  assign n225 = x0 | n224 ;
  assign n226 = ( x4 & ~x5 ) | ( x4 & x6 ) | ( ~x5 & x6 ) ;
  assign n227 = ( ~x4 & x5 ) | ( ~x4 & n226 ) | ( x5 & n226 ) ;
  assign n228 = x7 & ~n226 ;
  assign n229 = ( x6 & ~n226 ) | ( x6 & n228 ) | ( ~n226 & n228 ) ;
  assign n230 = n227 & ~n229 ;
  assign n231 = ( x2 & n10 ) | ( x2 & ~n230 ) | ( n10 & ~n230 ) ;
  assign n232 = n230 | n231 ;
  assign n233 = x0 | n232 ;
  assign n234 = ( x3 & x5 ) | ( x3 & ~x7 ) | ( x5 & ~x7 ) ;
  assign n235 = ( x3 & x4 ) | ( x3 & ~n234 ) | ( x4 & ~n234 ) ;
  assign n236 = ( ~x5 & x7 ) | ( ~x5 & n235 ) | ( x7 & n235 ) ;
  assign n237 = n234 | n236 ;
  assign n238 = ( ~n235 & n236 ) | ( ~n235 & n237 ) | ( n236 & n237 ) ;
  assign n244 = x6 & ~n238 ;
  assign n239 = n22 & ~n221 ;
  assign n240 = ( ~x3 & x4 ) | ( ~x3 & x5 ) | ( x4 & x5 ) ;
  assign n241 = x3 & ~n240 ;
  assign n242 = ( x6 & n71 ) | ( x6 & n241 ) | ( n71 & n241 ) ;
  assign n243 = n241 | n242 ;
  assign n245 = n239 | n243 ;
  assign n246 = ( n238 & n244 ) | ( n238 & ~n245 ) | ( n244 & ~n245 ) ;
  assign n247 = x0 | x2 ;
  assign n248 = ( x1 & ~n246 ) | ( x1 & n247 ) | ( ~n246 & n247 ) ;
  assign n249 = n246 | n248 ;
  assign n250 = ~x5 & x6 ;
  assign n251 = x6 & ~n250 ;
  assign n252 = x4 & n251 ;
  assign n253 = ( x3 & n250 ) | ( x3 & ~n251 ) | ( n250 & ~n251 ) ;
  assign n254 = ( x5 & ~n252 ) | ( x5 & n253 ) | ( ~n252 & n253 ) ;
  assign n258 = ( x3 & ~x5 ) | ( x3 & x6 ) | ( ~x5 & x6 ) ;
  assign n259 = ( x3 & ~x7 ) | ( x3 & n258 ) | ( ~x7 & n258 ) ;
  assign n260 = x3 & ~n259 ;
  assign n261 = n259 | n260 ;
  assign n262 = ( ~x3 & n260 ) | ( ~x3 & n261 ) | ( n260 & n261 ) ;
  assign n263 = x4 & ~n262 ;
  assign n255 = ( x5 & x6 ) | ( x5 & x7 ) | ( x6 & x7 ) ;
  assign n256 = ~x6 & n255 ;
  assign n257 = ( ~x5 & n255 ) | ( ~x5 & n256 ) | ( n255 & n256 ) ;
  assign n264 = ~x3 & n257 ;
  assign n265 = x4 | n264 ;
  assign n266 = ~n263 & n265 ;
  assign n267 = x2 & ~x3 ;
  assign n268 = ~x4 & x5 ;
  assign n269 = ( x3 & x4 ) | ( x3 & n268 ) | ( x4 & n268 ) ;
  assign n270 = ( ~x2 & x3 ) | ( ~x2 & n269 ) | ( x3 & n269 ) ;
  assign n271 = ( n267 & ~n269 ) | ( n267 & n270 ) | ( ~n269 & n270 ) ;
  assign n272 = ( n254 & n266 ) | ( n254 & n271 ) | ( n266 & n271 ) ;
  assign n273 = x2 & ~n271 ;
  assign n274 = ( n254 & ~n272 ) | ( n254 & n273 ) | ( ~n272 & n273 ) ;
  assign n275 = x1 | n274 ;
  assign n276 = x0 | n275 ;
  assign n280 = ( x3 & ~x4 ) | ( x3 & x6 ) | ( ~x4 & x6 ) ;
  assign n281 = ( x3 & ~x7 ) | ( x3 & n280 ) | ( ~x7 & n280 ) ;
  assign n282 = x3 & ~n281 ;
  assign n283 = n281 | n282 ;
  assign n284 = ( ~x3 & n282 ) | ( ~x3 & n283 ) | ( n282 & n283 ) ;
  assign n285 = x5 & ~n284 ;
  assign n277 = ( x4 & x7 ) | ( x4 & n162 ) | ( x7 & n162 ) ;
  assign n278 = ( ~x4 & x7 ) | ( ~x4 & n162 ) | ( x7 & n162 ) ;
  assign n279 = ( x4 & ~n277 ) | ( x4 & n278 ) | ( ~n277 & n278 ) ;
  assign n286 = x3 | n279 ;
  assign n287 = ~x5 & n286 ;
  assign n288 = n285 | n287 ;
  assign n289 = ~x2 & n288 ;
  assign n290 = n219 & ~n221 ;
  assign n291 = x2 & ~n290 ;
  assign n292 = n289 | n291 ;
  assign n311 = ( x0 & x1 ) | ( x0 & ~n292 ) | ( x1 & ~n292 ) ;
  assign n293 = ( x1 & ~x3 ) | ( x1 & x5 ) | ( ~x3 & x5 ) ;
  assign n294 = ( x2 & ~x5 ) | ( x2 & n293 ) | ( ~x5 & n293 ) ;
  assign n295 = ( ~x1 & x5 ) | ( ~x1 & n294 ) | ( x5 & n294 ) ;
  assign n296 = ~n293 & n295 ;
  assign n297 = x2 & ~n296 ;
  assign n298 = ( n294 & n296 ) | ( n294 & ~n297 ) | ( n296 & ~n297 ) ;
  assign n308 = x4 & n298 ;
  assign n299 = x2 & x4 ;
  assign n300 = ( x1 & x3 ) | ( x1 & n299 ) | ( x3 & n299 ) ;
  assign n301 = ~x1 & n300 ;
  assign n302 = x4 & x6 ;
  assign n303 = x1 & ~x6 ;
  assign n304 = x1 & n221 ;
  assign n305 = ( n302 & n303 ) | ( n302 & ~n304 ) | ( n303 & ~n304 ) ;
  assign n306 = x5 & n305 ;
  assign n307 = ~x2 & n306 ;
  assign n309 = n301 | n307 ;
  assign n310 = ( n298 & ~n308 ) | ( n298 & n309 ) | ( ~n308 & n309 ) ;
  assign n312 = ~x0 & n310 ;
  assign n313 = ( n292 & n311 ) | ( n292 & ~n312 ) | ( n311 & ~n312 ) ;
  assign n346 = ( x1 & x5 ) | ( x1 & ~x6 ) | ( x5 & ~x6 ) ;
  assign n347 = ( x1 & x4 ) | ( x1 & ~n250 ) | ( x4 & ~n250 ) ;
  assign n348 = ~n346 & n347 ;
  assign n352 = ( ~x2 & x3 ) | ( ~x2 & n348 ) | ( x3 & n348 ) ;
  assign n349 = ( ~x5 & n155 ) | ( ~x5 & n302 ) | ( n155 & n302 ) ;
  assign n350 = ( x5 & x6 ) | ( x5 & ~n155 ) | ( x6 & ~n155 ) ;
  assign n351 = ( ~x6 & n349 ) | ( ~x6 & n350 ) | ( n349 & n350 ) ;
  assign n353 = ( x2 & x3 ) | ( x2 & ~n351 ) | ( x3 & ~n351 ) ;
  assign n354 = n352 & ~n353 ;
  assign n339 = x1 | x2 ;
  assign n340 = x2 & ~n10 ;
  assign n341 = ( ~x2 & n339 ) | ( ~x2 & n340 ) | ( n339 & n340 ) ;
  assign n342 = ( x4 & x6 ) | ( x4 & n341 ) | ( x6 & n341 ) ;
  assign n343 = ( x5 & ~x6 ) | ( x5 & n342 ) | ( ~x6 & n342 ) ;
  assign n344 = ( x4 & x5 ) | ( x4 & ~n342 ) | ( x5 & ~n342 ) ;
  assign n345 = n343 & ~n344 ;
  assign n355 = ( x4 & x5 ) | ( x4 & ~n293 ) | ( x5 & ~n293 ) ;
  assign n356 = ( ~x1 & x3 ) | ( ~x1 & n355 ) | ( x3 & n355 ) ;
  assign n357 = n293 | n356 ;
  assign n358 = ( ~n355 & n356 ) | ( ~n355 & n357 ) | ( n356 & n357 ) ;
  assign n359 = ~x2 & n358 ;
  assign n325 = x3 & ~x4 ;
  assign n360 = ~x1 & n325 ;
  assign n361 = x2 & ~n360 ;
  assign n362 = n359 | n361 ;
  assign n363 = ~n345 & n362 ;
  assign n364 = ~n354 & n363 ;
  assign n317 = ( x1 & x3 ) | ( x1 & ~x7 ) | ( x3 & ~x7 ) ;
  assign n318 = ( x1 & x6 ) | ( x1 & ~n317 ) | ( x6 & ~n317 ) ;
  assign n319 = ( ~x3 & x7 ) | ( ~x3 & n318 ) | ( x7 & n318 ) ;
  assign n320 = n317 | n319 ;
  assign n321 = ( ~n318 & n319 ) | ( ~n318 & n320 ) | ( n319 & n320 ) ;
  assign n322 = x4 & ~n321 ;
  assign n314 = ( ~x3 & x6 ) | ( ~x3 & x7 ) | ( x6 & x7 ) ;
  assign n315 = ( x4 & x6 ) | ( x4 & x7 ) | ( x6 & x7 ) ;
  assign n316 = n314 & ~n315 ;
  assign n323 = n316 | n322 ;
  assign n324 = ( ~x1 & n322 ) | ( ~x1 & n323 ) | ( n322 & n323 ) ;
  assign n329 = ( x2 & ~x5 ) | ( x2 & n324 ) | ( ~x5 & n324 ) ;
  assign n326 = ~x5 & n325 ;
  assign n327 = ( x1 & n25 ) | ( x1 & n326 ) | ( n25 & n326 ) ;
  assign n328 = ~x1 & n327 ;
  assign n330 = ~x2 & n328 ;
  assign n331 = ( n324 & ~n329 ) | ( n324 & n330 ) | ( ~n329 & n330 ) ;
  assign n332 = ~x3 & x4 ;
  assign n333 = ( x5 & ~x7 ) | ( x5 & n332 ) | ( ~x7 & n332 ) ;
  assign n334 = ( x4 & x5 ) | ( x4 & ~n332 ) | ( x5 & ~n332 ) ;
  assign n335 = ( x3 & x7 ) | ( x3 & ~n334 ) | ( x7 & ~n334 ) ;
  assign n336 = n333 | n335 ;
  assign n337 = ( ~x6 & n154 ) | ( ~x6 & n336 ) | ( n154 & n336 ) ;
  assign n338 = ~n336 & n337 ;
  assign n365 = ( ~x0 & n331 ) | ( ~x0 & n338 ) | ( n331 & n338 ) ;
  assign n366 = n364 & n365 ;
  assign n367 = ( x0 & n364 ) | ( x0 & ~n366 ) | ( n364 & ~n366 ) ;
  assign n399 = ( x2 & ~x4 ) | ( x2 & x7 ) | ( ~x4 & x7 ) ;
  assign n397 = ~x3 & x6 ;
  assign n398 = ( n71 & n250 ) | ( n71 & ~n397 ) | ( n250 & ~n397 ) ;
  assign n400 = x2 | x7 ;
  assign n401 = ( ~x4 & n398 ) | ( ~x4 & n400 ) | ( n398 & n400 ) ;
  assign n402 = ~n399 & n401 ;
  assign n407 = ( x2 & n25 ) | ( x2 & n326 ) | ( n25 & n326 ) ;
  assign n408 = ~x2 & n407 ;
  assign n409 = x6 | x7 ;
  assign n403 = x2 & ~x4 ;
  assign n404 = ~x2 & x5 ;
  assign n405 = x3 & ~n404 ;
  assign n406 = ( n66 & n403 ) | ( n66 & ~n405 ) | ( n403 & ~n405 ) ;
  assign n410 = ( x6 & x7 ) | ( x6 & ~n406 ) | ( x7 & ~n406 ) ;
  assign n411 = ( n408 & n409 ) | ( n408 & ~n410 ) | ( n409 & ~n410 ) ;
  assign n412 = n402 | n411 ;
  assign n413 = x1 | n412 ;
  assign n396 = n9 & n14 ;
  assign n414 = n120 & n396 ;
  assign n415 = x1 & ~n414 ;
  assign n416 = n413 & ~n415 ;
  assign n369 = ( x5 & x6 ) | ( x5 & ~n280 ) | ( x6 & ~n280 ) ;
  assign n370 = ( ~x3 & x5 ) | ( ~x3 & n280 ) | ( x5 & n280 ) ;
  assign n371 = n369 & ~n370 ;
  assign n372 = x2 & ~n371 ;
  assign n373 = x3 | n119 ;
  assign n374 = ~x2 & n373 ;
  assign n375 = n372 | n374 ;
  assign n376 = ~x1 & n375 ;
  assign n368 = ~x4 & n121 ;
  assign n377 = ~n13 & n368 ;
  assign n378 = x1 & ~n377 ;
  assign n379 = n376 | n378 ;
  assign n384 = ( x3 & x7 ) | ( x3 & n9 ) | ( x7 & n9 ) ;
  assign n385 = ( x3 & x7 ) | ( x3 & ~n9 ) | ( x7 & ~n9 ) ;
  assign n386 = ( x4 & x5 ) | ( x4 & n385 ) | ( x5 & n385 ) ;
  assign n387 = ~n384 & n386 ;
  assign n388 = x2 | n387 ;
  assign n382 = ~x5 & x7 ;
  assign n383 = x4 & n382 ;
  assign n389 = x3 & n383 ;
  assign n390 = x2 & ~n389 ;
  assign n391 = n388 & ~n390 ;
  assign n392 = n154 & n326 ;
  assign n393 = ( ~x1 & n391 ) | ( ~x1 & n392 ) | ( n391 & n392 ) ;
  assign n380 = x2 | x4 ;
  assign n381 = ( x2 & ~x3 ) | ( x2 & n380 ) | ( ~x3 & n380 ) ;
  assign n394 = ( x1 & n381 ) | ( x1 & n392 ) | ( n381 & n392 ) ;
  assign n395 = n393 | n394 ;
  assign n417 = ( x0 & n379 ) | ( x0 & ~n395 ) | ( n379 & ~n395 ) ;
  assign n418 = n416 | n417 ;
  assign n419 = ( x0 & ~n416 ) | ( x0 & n418 ) | ( ~n416 & n418 ) ;
  assign y0 = ~x0 ;
  assign y1 = ~x0 ;
  assign y2 = ~x0 ;
  assign y3 = n20 ;
  assign y4 = ~n45 ;
  assign y5 = n88 ;
  assign y6 = ~n139 ;
  assign y7 = ~n211 ;
  assign y8 = ~n217 ;
  assign y9 = ~n225 ;
  assign y10 = ~n233 ;
  assign y11 = ~n249 ;
  assign y12 = ~n276 ;
  assign y13 = ~n313 ;
  assign y14 = ~n367 ;
  assign y15 = ~n419 ;
endmodule
