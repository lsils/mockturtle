module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159;
  wire n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770, n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778, n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794, n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802, n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842, n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866, n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874, n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914, n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922, n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930, n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938, n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946, n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986, n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994, n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010, n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018, n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058, n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066, n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074, n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082, n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090, n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130, n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138, n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146, n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154, n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162, n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202, n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218, n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226, n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234, n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274, n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282, n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306, n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346, n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362, n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370, n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378, n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418, n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426, n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442, n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450, n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490, n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514, n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522, n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562, n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722, n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730, n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738, n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746, n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754, n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762, n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770, n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778, n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786, n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794, n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802, n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810, n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818, n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826, n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834, n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842, n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850, n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858, n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866, n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874, n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882, n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890, n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898, n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906, n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914, n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922, n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930, n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938, n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946, n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954, n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962, n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970, n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978, n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986, n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994, n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002, n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010, n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018, n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026, n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034, n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042, n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050, n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058, n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066, n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074, n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082, n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090, n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098, n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106, n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114, n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122, n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130, n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138, n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146, n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154, n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162, n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170, n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178, n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186, n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194, n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202, n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210, n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218, n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226, n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234, n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242, n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250, n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258, n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266, n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274, n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282, n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290, n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298, n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306, n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314, n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322, n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330, n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338, n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346, n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354, n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362, n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370, n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378, n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386, n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394, n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402, n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410, n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418, n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426, n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434, n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442, n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450, n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458, n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466, n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474, n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482, n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490, n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498, n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506, n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514, n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522, n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530, n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538, n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546, n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554, n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562, n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570, n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578, n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586, n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594, n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602, n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610, n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618, n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626, n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634, n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642, n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650, n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658, n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666, n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674, n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682, n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690, n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698, n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706, n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714, n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722, n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730, n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738, n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746, n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754, n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762, n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770, n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778, n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786, n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794, n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802, n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810, n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818, n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826, n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834, n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842, n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850, n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858, n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866, n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874, n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882, n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890, n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898, n54899, n54900, n54901, n54902, n54903, n54904, n54905, n54906, n54907, n54908, n54909, n54910, n54911, n54912, n54913, n54914, n54915, n54916, n54917, n54918, n54919, n54920, n54921, n54922, n54923, n54924, n54925, n54926, n54927, n54928, n54929, n54930, n54931, n54932, n54933, n54934, n54935, n54936, n54937, n54938, n54939, n54940, n54941, n54942, n54943, n54944, n54945, n54946, n54947, n54948, n54949, n54950, n54951, n54952, n54953, n54954, n54955, n54956, n54957, n54958, n54959, n54960, n54961, n54962, n54963, n54964, n54965, n54966, n54967, n54968, n54969, n54970, n54971, n54972, n54973, n54974, n54975, n54976, n54977, n54978, n54979, n54980, n54981, n54982, n54983, n54984, n54985, n54986, n54987, n54988, n54989, n54990, n54991, n54992, n54993, n54994, n54995, n54996, n54997, n54998, n54999, n55000, n55001, n55002, n55003, n55004, n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012, n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020, n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028, n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036, n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044, n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052, n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060, n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068, n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076, n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084, n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092, n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100, n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108, n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116, n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124, n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132, n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140, n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148, n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156, n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164, n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172, n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180, n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188, n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196, n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204, n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212, n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220, n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228, n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236, n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244, n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252, n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260, n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268, n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276, n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284, n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292, n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300, n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308, n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316, n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324, n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332, n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340, n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348, n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356, n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364, n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372, n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380, n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388, n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396, n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404, n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412, n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420, n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428, n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436, n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444, n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452, n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460, n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468, n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476, n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484, n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492, n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500, n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508, n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516, n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524, n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532, n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540, n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548, n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556, n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564, n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572, n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580, n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588, n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596, n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604, n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612, n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620, n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628, n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636, n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644, n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652, n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660, n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668, n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676, n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684, n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692, n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700, n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708, n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716, n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724, n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732, n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740, n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748, n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756, n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764, n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772, n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780, n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788, n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796, n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804, n55805, n55806, n55807, n55808, n55809, n55810, n55811, n55812, n55813, n55814, n55815, n55816, n55817, n55818, n55819, n55820, n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828, n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836, n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844, n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852, n55853, n55854, n55855, n55856, n55857, n55858, n55859, n55860, n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868, n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876, n55877, n55878, n55879, n55880, n55881, n55882, n55883, n55884, n55885, n55886, n55887, n55888, n55889, n55890, n55891, n55892, n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900, n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908, n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916, n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924, n55925, n55926, n55927, n55928, n55929, n55930, n55931, n55932, n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940, n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948, n55949, n55950, n55951, n55952, n55953, n55954, n55955, n55956, n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964, n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972, n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980, n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988, n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996, n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004, n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012, n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020, n56021, n56022, n56023, n56024, n56025, n56026, n56027, n56028, n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036, n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044, n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052, n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060, n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068, n56069, n56070, n56071, n56072, n56073, n56074, n56075, n56076, n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084, n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092, n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100, n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108, n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116, n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124, n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132, n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140, n56141, n56142, n56143, n56144, n56145, n56146, n56147, n56148, n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156, n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164, n56165, n56166, n56167, n56168, n56169, n56170, n56171, n56172, n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180, n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188, n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196, n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204, n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212, n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220, n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228, n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236, n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244, n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252, n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260, n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268, n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276, n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284, n56285, n56286, n56287, n56288, n56289, n56290, n56291, n56292, n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300, n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308, n56309, n56310, n56311, n56312, n56313, n56314, n56315, n56316, n56317, n56318, n56319, n56320, n56321, n56322, n56323, n56324, n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332, n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340, n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348, n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356, n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364, n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372, n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380, n56381, n56382, n56383, n56384, n56385, n56386, n56387, n56388, n56389, n56390, n56391, n56392, n56393, n56394, n56395, n56396, n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404, n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412, n56413, n56414, n56415, n56416, n56417, n56418, n56419, n56420, n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428, n56429, n56430, n56431, n56432, n56433, n56434, n56435, n56436, n56437, n56438, n56439, n56440, n56441, n56442, n56443, n56444, n56445, n56446, n56447, n56448, n56449, n56450, n56451, n56452, n56453, n56454, n56455, n56456, n56457, n56458, n56459, n56460, n56461, n56462, n56463, n56464, n56465, n56466, n56467, n56468, n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476, n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484, n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492, n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500, n56501, n56502, n56503, n56504, n56505, n56506, n56507, n56508, n56509, n56510, n56511, n56512, n56513, n56514, n56515, n56516, n56517, n56518, n56519, n56520, n56521, n56522, n56523, n56524, n56525, n56526, n56527, n56528, n56529, n56530, n56531, n56532, n56533, n56534, n56535, n56536, n56537, n56538, n56539, n56540, n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548, n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556, n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564, n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572, n56573, n56574, n56575, n56576, n56577, n56578, n56579, n56580, n56581, n56582, n56583, n56584, n56585, n56586, n56587, n56588, n56589, n56590, n56591, n56592, n56593, n56594, n56595, n56596, n56597, n56598, n56599, n56600, n56601, n56602, n56603, n56604, n56605, n56606, n56607, n56608, n56609, n56610, n56611, n56612, n56613, n56614, n56615, n56616, n56617, n56618, n56619, n56620, n56621, n56622, n56623, n56624, n56625, n56626, n56627, n56628, n56629, n56630, n56631, n56632, n56633, n56634, n56635, n56636, n56637, n56638, n56639, n56640, n56641, n56642, n56643;
  assign n13252 = x449 ^ x97;
  assign n13253 = n13252 ^ x289;
  assign n13254 = n13253 ^ x33;
  assign n14745 = n13254 ^ x192;
  assign n14746 = n14745 ^ x384;
  assign n14747 = n14746 ^ x128;
  assign n16787 = n14747 ^ x319;
  assign n16788 = n16787 ^ x511;
  assign n16789 = n16788 ^ x255;
  assign n18368 = n16789 ^ x414;
  assign n13341 = x511 ^ x159;
  assign n13342 = n13341 ^ x351;
  assign n13343 = n13342 ^ x95;
  assign n18369 = n18368 ^ n13343;
  assign n18370 = n18369 ^ x350;
  assign n20264 = n18370 ^ x509;
  assign n15253 = n13343 ^ x254;
  assign n15254 = n15253 ^ x446;
  assign n15255 = n15254 ^ x190;
  assign n20265 = n20264 ^ n15255;
  assign n20266 = n20265 ^ x445;
  assign n1715 = x509 ^ x157;
  assign n1716 = n1715 ^ x349;
  assign n1717 = n1716 ^ x93;
  assign n22379 = n20266 ^ n1717;
  assign n17476 = n15255 ^ x349;
  assign n1442 = x446 ^ x94;
  assign n1443 = n1442 ^ x286;
  assign n1444 = n1443 ^ x30;
  assign n17477 = n17476 ^ n1444;
  assign n17478 = n17477 ^ x285;
  assign n22380 = n22379 ^ n17478;
  assign n1593 = x445 ^ x93;
  assign n1594 = n1593 ^ x285;
  assign n1595 = n1594 ^ x29;
  assign n22381 = n22380 ^ n1595;
  assign n1781 = n1717 ^ x252;
  assign n1782 = n1781 ^ x444;
  assign n1783 = n1782 ^ x188;
  assign n24186 = n22381 ^ n1783;
  assign n19349 = n17478 ^ x444;
  assign n1457 = n1444 ^ x189;
  assign n1458 = n1457 ^ x381;
  assign n1459 = n1458 ^ x125;
  assign n19350 = n19349 ^ n1459;
  assign n19351 = n19350 ^ x380;
  assign n24187 = n24186 ^ n19351;
  assign n1638 = n1595 ^ x188;
  assign n1639 = n1638 ^ x380;
  assign n1640 = n1639 ^ x124;
  assign n24188 = n24187 ^ n1640;
  assign n1856 = n1783 ^ x347;
  assign n1853 = x444 ^ x92;
  assign n1854 = n1853 ^ x284;
  assign n1855 = n1854 ^ x28;
  assign n1857 = n1856 ^ n1855;
  assign n1858 = n1857 ^ x283;
  assign n26140 = n24188 ^ n1858;
  assign n20827 = n19351 ^ n1855;
  assign n1626 = n1459 ^ x284;
  assign n1627 = n1626 ^ x476;
  assign n1628 = n1627 ^ x220;
  assign n20828 = n20827 ^ n1628;
  assign n20829 = n20828 ^ x475;
  assign n26141 = n26140 ^ n20829;
  assign n1686 = n1640 ^ x283;
  assign n1687 = n1686 ^ x475;
  assign n1688 = n1687 ^ x219;
  assign n26142 = n26141 ^ n1688;
  assign n1940 = n1858 ^ x442;
  assign n1937 = n1855 ^ x187;
  assign n1938 = n1937 ^ x379;
  assign n1939 = n1938 ^ x123;
  assign n1941 = n1940 ^ n1939;
  assign n1942 = n1941 ^ x378;
  assign n28554 = n26142 ^ n1942;
  assign n23098 = n20829 ^ n1939;
  assign n1655 = n1628 ^ x379;
  assign n1650 = x476 ^ x124;
  assign n1651 = n1650 ^ x316;
  assign n1652 = n1651 ^ x60;
  assign n1656 = n1655 ^ n1652;
  assign n1657 = n1656 ^ x315;
  assign n23099 = n23098 ^ n1657;
  assign n1749 = x475 ^ x123;
  assign n1750 = n1749 ^ x315;
  assign n1751 = n1750 ^ x59;
  assign n23100 = n23099 ^ n1751;
  assign n28555 = n28554 ^ n23100;
  assign n1752 = n1688 ^ x378;
  assign n1753 = n1752 ^ n1751;
  assign n1754 = n1753 ^ x314;
  assign n28556 = n28555 ^ n1754;
  assign n1869 = x442 ^ x90;
  assign n1870 = n1869 ^ x282;
  assign n1871 = n1870 ^ x26;
  assign n2030 = n1942 ^ n1871;
  assign n2027 = n1939 ^ x282;
  assign n2028 = n2027 ^ x474;
  assign n2029 = n2028 ^ x218;
  assign n2031 = n2030 ^ n2029;
  assign n2032 = n2031 ^ x473;
  assign n30587 = n28556 ^ n2032;
  assign n24992 = n23100 ^ n2029;
  assign n1706 = n1657 ^ x474;
  assign n1701 = n1652 ^ x155;
  assign n1702 = n1701 ^ x411;
  assign n1703 = n1702 ^ x219;
  assign n1707 = n1706 ^ n1703;
  assign n1708 = n1707 ^ x410;
  assign n24993 = n24992 ^ n1708;
  assign n1815 = n1751 ^ x218;
  assign n1816 = n1815 ^ x410;
  assign n1817 = n1816 ^ x154;
  assign n24994 = n24993 ^ n1817;
  assign n30588 = n30587 ^ n24994;
  assign n1818 = n1754 ^ x473;
  assign n1819 = n1818 ^ n1817;
  assign n1820 = n1819 ^ x409;
  assign n30589 = n30588 ^ n1820;
  assign n1689 = x443 ^ x91;
  assign n1690 = n1689 ^ x283;
  assign n1691 = n1690 ^ x27;
  assign n1755 = n1691 ^ x186;
  assign n1756 = n1755 ^ x378;
  assign n1757 = n1756 ^ x122;
  assign n1821 = n1757 ^ x281;
  assign n1822 = n1821 ^ x473;
  assign n1823 = n1822 ^ x217;
  assign n1437 = x510 ^ x158;
  assign n1438 = n1437 ^ x350;
  assign n1439 = n1438 ^ x94;
  assign n1446 = n1439 ^ x253;
  assign n1447 = n1446 ^ x445;
  assign n1448 = n1447 ^ x189;
  assign n1621 = n1448 ^ x348;
  assign n1622 = n1621 ^ n1595;
  assign n1623 = n1622 ^ x284;
  assign n1641 = n1623 ^ x443;
  assign n1642 = n1641 ^ n1640;
  assign n1643 = n1642 ^ x379;
  assign n1692 = n1691 ^ n1643;
  assign n1693 = n1692 ^ n1688;
  assign n1694 = n1693 ^ x474;
  assign n1758 = n1757 ^ n1694;
  assign n1759 = n1758 ^ n1754;
  assign n1746 = x474 ^ x122;
  assign n1747 = n1746 ^ x314;
  assign n1748 = n1747 ^ x58;
  assign n1760 = n1759 ^ n1748;
  assign n1824 = n1823 ^ n1760;
  assign n1825 = n1824 ^ n1820;
  assign n1812 = n1748 ^ x217;
  assign n1813 = n1812 ^ x409;
  assign n1814 = n1813 ^ x153;
  assign n1826 = n1825 ^ n1814;
  assign n36689 = n30589 ^ n1826;
  assign n2536 = x419 ^ x67;
  assign n2537 = n2536 ^ x259;
  assign n2538 = n2537 ^ x3;
  assign n2614 = n2538 ^ x162;
  assign n2615 = n2614 ^ x354;
  assign n2616 = n2615 ^ x98;
  assign n16399 = n2616 ^ x257;
  assign n16400 = n16399 ^ x449;
  assign n16401 = n16400 ^ x193;
  assign n17762 = n16401 ^ x352;
  assign n17763 = n17762 ^ n13254;
  assign n17764 = n17763 ^ x288;
  assign n19682 = n17764 ^ x479;
  assign n19683 = n19682 ^ n14747;
  assign n19684 = n19683 ^ x415;
  assign n1570 = x479 ^ x127;
  assign n1571 = n1570 ^ x319;
  assign n1572 = n1571 ^ x63;
  assign n21562 = n19684 ^ n1572;
  assign n21563 = n21562 ^ n16789;
  assign n21564 = n21563 ^ x510;
  assign n1605 = n1572 ^ x222;
  assign n1606 = n1605 ^ x414;
  assign n1607 = n1606 ^ x158;
  assign n23390 = n21564 ^ n1607;
  assign n23391 = n23390 ^ n18370;
  assign n23392 = n23391 ^ n1439;
  assign n1663 = n1607 ^ x317;
  assign n1664 = n1663 ^ x509;
  assign n1665 = n1664 ^ x253;
  assign n25644 = n23392 ^ n1665;
  assign n25645 = n25644 ^ n20266;
  assign n25646 = n25645 ^ n1448;
  assign n1714 = n1665 ^ x412;
  assign n1718 = n1717 ^ n1714;
  assign n1719 = n1718 ^ x348;
  assign n27623 = n25646 ^ n1719;
  assign n27624 = n27623 ^ n22381;
  assign n27625 = n27624 ^ n1623;
  assign n1780 = n1719 ^ x507;
  assign n1784 = n1783 ^ n1780;
  assign n1785 = n1784 ^ x443;
  assign n29702 = n27625 ^ n1785;
  assign n29703 = n29702 ^ n24188;
  assign n29704 = n29703 ^ n1643;
  assign n1733 = x507 ^ x155;
  assign n1734 = n1733 ^ x347;
  assign n1735 = n1734 ^ x91;
  assign n1852 = n1785 ^ n1735;
  assign n1859 = n1858 ^ n1852;
  assign n1860 = n1859 ^ n1691;
  assign n31887 = n29704 ^ n1860;
  assign n31888 = n31887 ^ n26142;
  assign n31889 = n31888 ^ n1694;
  assign n1799 = n1735 ^ x250;
  assign n1800 = n1799 ^ x442;
  assign n1801 = n1800 ^ x186;
  assign n1936 = n1860 ^ n1801;
  assign n1943 = n1942 ^ n1936;
  assign n1944 = n1943 ^ n1757;
  assign n34735 = n31889 ^ n1944;
  assign n34736 = n34735 ^ n28556;
  assign n34737 = n34736 ^ n1760;
  assign n1877 = n1801 ^ x345;
  assign n1878 = n1877 ^ n1871;
  assign n1879 = n1878 ^ x281;
  assign n2026 = n1944 ^ n1879;
  assign n2033 = n2032 ^ n2026;
  assign n2034 = n2033 ^ n1823;
  assign n36688 = n34737 ^ n2034;
  assign n36690 = n36689 ^ n36688;
  assign n1961 = n1879 ^ x440;
  assign n1953 = n1871 ^ x185;
  assign n1954 = n1953 ^ x377;
  assign n1955 = n1954 ^ x121;
  assign n1962 = n1961 ^ n1955;
  assign n1963 = n1962 ^ x376;
  assign n2122 = n2034 ^ n1963;
  assign n2119 = n2032 ^ n1955;
  assign n2116 = n2029 ^ x377;
  assign n2117 = n2116 ^ n1748;
  assign n2118 = n2117 ^ x313;
  assign n2120 = n2119 ^ n2118;
  assign n1897 = x473 ^ x121;
  assign n1898 = n1897 ^ x313;
  assign n1899 = n1898 ^ x57;
  assign n2121 = n2120 ^ n1899;
  assign n2123 = n2122 ^ n2121;
  assign n1896 = n1823 ^ x376;
  assign n1900 = n1899 ^ n1896;
  assign n1901 = n1900 ^ x312;
  assign n2124 = n2123 ^ n1901;
  assign n39186 = n36690 ^ n2124;
  assign n27010 = n24994 ^ n2118;
  assign n1772 = n1748 ^ n1708;
  assign n1767 = n1703 ^ x314;
  assign n1768 = n1767 ^ x506;
  assign n1769 = n1768 ^ x250;
  assign n1773 = n1772 ^ n1769;
  assign n1774 = n1773 ^ x505;
  assign n27011 = n27010 ^ n1774;
  assign n1904 = n1817 ^ x313;
  assign n1905 = n1904 ^ x505;
  assign n1906 = n1905 ^ x249;
  assign n27012 = n27011 ^ n1906;
  assign n32745 = n27012 ^ n2121;
  assign n32746 = n32745 ^ n30589;
  assign n1903 = n1899 ^ n1820;
  assign n1907 = n1906 ^ n1903;
  assign n1908 = n1907 ^ x504;
  assign n32747 = n32746 ^ n1908;
  assign n39187 = n39186 ^ n32747;
  assign n1902 = n1901 ^ n1826;
  assign n1909 = n1908 ^ n1902;
  assign n1893 = n1814 ^ x312;
  assign n1894 = n1893 ^ x504;
  assign n1895 = n1894 ^ x248;
  assign n1910 = n1909 ^ n1895;
  assign n39188 = n39187 ^ n1910;
  assign n2009 = x440 ^ x88;
  assign n2010 = n2009 ^ x280;
  assign n2011 = n2010 ^ x24;
  assign n2051 = n2011 ^ n1963;
  assign n2043 = n1955 ^ x280;
  assign n2044 = n2043 ^ x472;
  assign n2045 = n2044 ^ x216;
  assign n2052 = n2051 ^ n2045;
  assign n2053 = n2052 ^ x471;
  assign n2227 = n2124 ^ n2053;
  assign n2224 = n2121 ^ n2045;
  assign n2221 = n2118 ^ x472;
  assign n2222 = n2221 ^ n1814;
  assign n2223 = n2222 ^ x408;
  assign n2225 = n2224 ^ n2223;
  assign n1984 = n1899 ^ x216;
  assign n1985 = n1984 ^ x408;
  assign n1986 = n1985 ^ x152;
  assign n2226 = n2225 ^ n1986;
  assign n2228 = n2227 ^ n2226;
  assign n1983 = n1901 ^ x471;
  assign n1987 = n1986 ^ n1983;
  assign n1988 = n1987 ^ x407;
  assign n2229 = n2228 ^ n1988;
  assign n41509 = n39188 ^ n2229;
  assign n35669 = n32747 ^ n2226;
  assign n28864 = n27012 ^ n2223;
  assign n1844 = n1814 ^ n1774;
  assign n1836 = n1769 ^ x409;
  assign n1831 = x506 ^ x154;
  assign n1832 = n1831 ^ x346;
  assign n1833 = n1832 ^ x90;
  assign n1837 = n1836 ^ n1833;
  assign n1838 = n1837 ^ x345;
  assign n1845 = n1844 ^ n1838;
  assign n1841 = x505 ^ x153;
  assign n1842 = n1841 ^ x345;
  assign n1843 = n1842 ^ x89;
  assign n1846 = n1845 ^ n1843;
  assign n28865 = n28864 ^ n1846;
  assign n1991 = n1906 ^ x408;
  assign n1992 = n1991 ^ n1843;
  assign n1993 = n1992 ^ x344;
  assign n28866 = n28865 ^ n1993;
  assign n35670 = n35669 ^ n28866;
  assign n1990 = n1986 ^ n1908;
  assign n1994 = n1993 ^ n1990;
  assign n1978 = x504 ^ x152;
  assign n1979 = n1978 ^ x344;
  assign n1980 = n1979 ^ x88;
  assign n1995 = n1994 ^ n1980;
  assign n35671 = n35670 ^ n1995;
  assign n41510 = n41509 ^ n35671;
  assign n1989 = n1988 ^ n1910;
  assign n1996 = n1995 ^ n1989;
  assign n1977 = n1895 ^ x407;
  assign n1981 = n1980 ^ n1977;
  assign n1982 = n1981 ^ x343;
  assign n1997 = n1996 ^ n1982;
  assign n41511 = n41510 ^ n1997;
  assign n2099 = n2011 ^ x183;
  assign n2100 = n2099 ^ x375;
  assign n2101 = n2100 ^ x119;
  assign n2144 = n2101 ^ n2053;
  assign n2136 = n2045 ^ x375;
  assign n2128 = x472 ^ x120;
  assign n2129 = n2128 ^ x312;
  assign n2130 = n2129 ^ x56;
  assign n2137 = n2136 ^ n2130;
  assign n2138 = n2137 ^ x311;
  assign n2145 = n2144 ^ n2138;
  assign n576 = x471 ^ x119;
  assign n577 = n576 ^ x311;
  assign n578 = n577 ^ x55;
  assign n2146 = n2145 ^ n578;
  assign n33218 = n2229 ^ n2146;
  assign n26953 = n2226 ^ n2138;
  assign n21605 = n2223 ^ n2130;
  assign n21606 = n21605 ^ n1895;
  assign n21607 = n21606 ^ x503;
  assign n26954 = n26953 ^ n21607;
  assign n2074 = n1986 ^ x311;
  assign n2075 = n2074 ^ x503;
  assign n2076 = n2075 ^ x247;
  assign n26955 = n26954 ^ n2076;
  assign n33219 = n33218 ^ n26955;
  assign n2073 = n1988 ^ n578;
  assign n2077 = n2076 ^ n2073;
  assign n2078 = n2077 ^ x502;
  assign n33220 = n33219 ^ n2078;
  assign n43557 = n41511 ^ n33220;
  assign n37938 = n35671 ^ n26955;
  assign n31217 = n28866 ^ n21607;
  assign n1928 = n1895 ^ n1846;
  assign n1920 = n1838 ^ x504;
  assign n1915 = n1833 ^ x249;
  assign n1916 = n1915 ^ x441;
  assign n1917 = n1916 ^ x185;
  assign n1921 = n1920 ^ n1917;
  assign n1922 = n1921 ^ x440;
  assign n1929 = n1928 ^ n1922;
  assign n1925 = n1843 ^ x248;
  assign n1926 = n1925 ^ x440;
  assign n1927 = n1926 ^ x184;
  assign n1930 = n1929 ^ n1927;
  assign n31218 = n31217 ^ n1930;
  assign n2081 = n1993 ^ x503;
  assign n2082 = n2081 ^ n1927;
  assign n2083 = n2082 ^ x439;
  assign n31219 = n31218 ^ n2083;
  assign n37939 = n37938 ^ n31219;
  assign n2080 = n2076 ^ n1995;
  assign n2084 = n2083 ^ n2080;
  assign n2068 = n1980 ^ x247;
  assign n2069 = n2068 ^ x439;
  assign n2070 = n2069 ^ x183;
  assign n2085 = n2084 ^ n2070;
  assign n37940 = n37939 ^ n2085;
  assign n43558 = n43557 ^ n37940;
  assign n2079 = n2078 ^ n1997;
  assign n2086 = n2085 ^ n2079;
  assign n2067 = n1982 ^ x502;
  assign n2071 = n2070 ^ n2067;
  assign n2072 = n2071 ^ x438;
  assign n2087 = n2086 ^ n2072;
  assign n43559 = n43558 ^ n2087;
  assign n2204 = n2101 ^ x278;
  assign n2205 = n2204 ^ x470;
  assign n2206 = n2205 ^ x214;
  assign n2248 = n2206 ^ n2146;
  assign n2241 = n2138 ^ x470;
  assign n2233 = n2130 ^ x215;
  assign n2234 = n2233 ^ x407;
  assign n2235 = n2234 ^ x151;
  assign n2242 = n2241 ^ n2235;
  assign n2243 = n2242 ^ x406;
  assign n2249 = n2248 ^ n2243;
  assign n579 = n578 ^ x214;
  assign n580 = n579 ^ x406;
  assign n581 = n580 ^ x150;
  assign n2250 = n2249 ^ n581;
  assign n35659 = n33220 ^ n2250;
  assign n2179 = n2076 ^ x406;
  assign n2176 = x503 ^ x151;
  assign n2177 = n2176 ^ x343;
  assign n2178 = n2177 ^ x87;
  assign n2180 = n2179 ^ n2178;
  assign n2181 = n2180 ^ x342;
  assign n29322 = n26955 ^ n2181;
  assign n23450 = n21607 ^ n2235;
  assign n23451 = n23450 ^ n1982;
  assign n23452 = n23451 ^ n2178;
  assign n29323 = n29322 ^ n23452;
  assign n29324 = n29323 ^ n2243;
  assign n35660 = n35659 ^ n29324;
  assign n2175 = n2078 ^ n581;
  assign n2182 = n2181 ^ n2175;
  assign n2163 = x502 ^ x150;
  assign n2164 = n2163 ^ x342;
  assign n2165 = n2164 ^ x86;
  assign n2183 = n2182 ^ n2165;
  assign n35661 = n35660 ^ n2183;
  assign n45602 = n43559 ^ n35661;
  assign n39963 = n37940 ^ n29324;
  assign n2018 = n1982 ^ n1930;
  assign n2007 = n1980 ^ n1922;
  assign n2002 = n1917 ^ x344;
  assign n1887 = x441 ^ x89;
  assign n1888 = n1887 ^ x281;
  assign n1889 = n1888 ^ x25;
  assign n2003 = n2002 ^ n1889;
  assign n2004 = n2003 ^ x280;
  assign n2008 = n2007 ^ n2004;
  assign n2012 = n2011 ^ n2008;
  assign n2019 = n2018 ^ n2012;
  assign n2015 = n1927 ^ x343;
  assign n2016 = n2015 ^ n2011;
  assign n2017 = n2016 ^ x279;
  assign n2020 = n2019 ^ n2017;
  assign n33654 = n31219 ^ n2020;
  assign n2186 = n2178 ^ n2083;
  assign n2187 = n2186 ^ n2017;
  assign n2168 = x439 ^ x87;
  assign n2169 = n2168 ^ x279;
  assign n2170 = n2169 ^ x23;
  assign n2188 = n2187 ^ n2170;
  assign n33655 = n33654 ^ n2188;
  assign n33656 = n33655 ^ n23452;
  assign n39964 = n39963 ^ n33656;
  assign n2185 = n2181 ^ n2085;
  assign n2189 = n2188 ^ n2185;
  assign n2167 = n2070 ^ x342;
  assign n2171 = n2170 ^ n2167;
  assign n2172 = n2171 ^ x278;
  assign n2190 = n2189 ^ n2172;
  assign n39965 = n39964 ^ n2190;
  assign n45603 = n45602 ^ n39965;
  assign n2184 = n2183 ^ n2087;
  assign n2191 = n2190 ^ n2184;
  assign n2166 = n2165 ^ n2072;
  assign n2173 = n2172 ^ n2166;
  assign n2160 = x438 ^ x86;
  assign n2161 = n2160 ^ x278;
  assign n2162 = n2161 ^ x22;
  assign n2174 = n2173 ^ n2162;
  assign n2192 = n2191 ^ n2174;
  assign n45604 = n45603 ^ n2192;
  assign n17816 = n2206 ^ x373;
  assign n12790 = x470 ^ x118;
  assign n12791 = n12790 ^ x310;
  assign n12792 = n12791 ^ x54;
  assign n17817 = n17816 ^ n12792;
  assign n17818 = n17817 ^ x309;
  assign n26943 = n17818 ^ n2250;
  assign n21546 = n12792 ^ n2243;
  assign n16828 = n2235 ^ x310;
  assign n16829 = n16828 ^ x502;
  assign n16830 = n16829 ^ x246;
  assign n21547 = n21546 ^ n16830;
  assign n21548 = n21547 ^ x501;
  assign n26944 = n26943 ^ n21548;
  assign n582 = n581 ^ x309;
  assign n583 = n582 ^ x501;
  assign n584 = n583 ^ x245;
  assign n26945 = n26944 ^ n584;
  assign n37933 = n35661 ^ n26945;
  assign n31210 = n29324 ^ n21548;
  assign n25693 = n23452 ^ n16830;
  assign n25694 = n25693 ^ n2072;
  assign n15307 = n2178 ^ x246;
  assign n15308 = n15307 ^ x438;
  assign n15309 = n15308 ^ x182;
  assign n25695 = n25694 ^ n15309;
  assign n31211 = n31210 ^ n25695;
  assign n20326 = n2181 ^ x501;
  assign n20327 = n20326 ^ n15309;
  assign n20328 = n20327 ^ x437;
  assign n31212 = n31211 ^ n20328;
  assign n37934 = n37933 ^ n31212;
  assign n25699 = n2183 ^ n584;
  assign n25700 = n25699 ^ n20328;
  assign n15597 = n2165 ^ x245;
  assign n15598 = n15597 ^ x437;
  assign n15599 = n15598 ^ x181;
  assign n25701 = n25700 ^ n15599;
  assign n37935 = n37934 ^ n25701;
  assign n47748 = n45604 ^ n37935;
  assign n42127 = n39965 ^ n31212;
  assign n35951 = n33656 ^ n25695;
  assign n2108 = n2072 ^ n2020;
  assign n2097 = n2070 ^ n2012;
  assign n2092 = n2004 ^ x439;
  assign n1971 = n1889 ^ x184;
  assign n1972 = n1971 ^ x376;
  assign n1973 = n1972 ^ x120;
  assign n2093 = n2092 ^ n1973;
  assign n2094 = n2093 ^ x375;
  assign n2098 = n2097 ^ n2094;
  assign n2102 = n2101 ^ n2098;
  assign n2109 = n2108 ^ n2102;
  assign n2105 = n2017 ^ x438;
  assign n2106 = n2105 ^ n2101;
  assign n2107 = n2106 ^ x374;
  assign n2110 = n2109 ^ n2107;
  assign n35952 = n35951 ^ n2110;
  assign n24172 = n15309 ^ n2188;
  assign n24173 = n24172 ^ n2107;
  assign n14145 = n2170 ^ x182;
  assign n14146 = n14145 ^ x374;
  assign n14147 = n14146 ^ x118;
  assign n24174 = n24173 ^ n14147;
  assign n35953 = n35952 ^ n24174;
  assign n42128 = n42127 ^ n35953;
  assign n29644 = n20328 ^ n2190;
  assign n29645 = n29644 ^ n24174;
  assign n19336 = n2172 ^ x437;
  assign n19337 = n19336 ^ n14147;
  assign n19338 = n19337 ^ x373;
  assign n29646 = n29645 ^ n19338;
  assign n42129 = n42128 ^ n29646;
  assign n47749 = n47748 ^ n42129;
  assign n36038 = n25701 ^ n2192;
  assign n36039 = n36038 ^ n29646;
  assign n24247 = n15599 ^ n2174;
  assign n24248 = n24247 ^ n19338;
  assign n14093 = n2162 ^ x181;
  assign n14094 = n14093 ^ x373;
  assign n14095 = n14094 ^ x117;
  assign n24249 = n24248 ^ n14095;
  assign n36040 = n36039 ^ n24249;
  assign n47750 = n47749 ^ n36040;
  assign n19657 = n17818 ^ x468;
  assign n14729 = n12792 ^ x213;
  assign n14730 = n14729 ^ x405;
  assign n14731 = n14730 ^ x149;
  assign n19658 = n19657 ^ n14731;
  assign n19659 = n19658 ^ x404;
  assign n29312 = n26945 ^ n19659;
  assign n23845 = n21548 ^ n14731;
  assign n18704 = n16830 ^ x405;
  assign n18705 = n18704 ^ n2165;
  assign n18706 = n18705 ^ x341;
  assign n23846 = n23845 ^ n18706;
  assign n586 = x501 ^ x149;
  assign n587 = n586 ^ x341;
  assign n588 = n587 ^ x85;
  assign n23847 = n23846 ^ n588;
  assign n29313 = n29312 ^ n23847;
  assign n585 = n584 ^ x404;
  assign n589 = n588 ^ n585;
  assign n590 = n589 ^ x340;
  assign n29314 = n29313 ^ n590;
  assign n39866 = n37935 ^ n29314;
  assign n27607 = n25695 ^ n18706;
  assign n27608 = n27607 ^ n2174;
  assign n17459 = n15309 ^ x341;
  assign n17460 = n17459 ^ n2162;
  assign n17461 = n17460 ^ x277;
  assign n27609 = n27608 ^ n17461;
  assign n33735 = n27609 ^ n23847;
  assign n33736 = n33735 ^ n31212;
  assign n22440 = n20328 ^ n588;
  assign n22441 = n22440 ^ n17461;
  assign n12455 = x437 ^ x85;
  assign n12456 = n12455 ^ x277;
  assign n12457 = n12456 ^ x21;
  assign n22442 = n22441 ^ n12457;
  assign n33737 = n33736 ^ n22442;
  assign n39867 = n39866 ^ n33737;
  assign n27602 = n25701 ^ n590;
  assign n27603 = n27602 ^ n22442;
  assign n17454 = n15599 ^ x340;
  assign n17455 = n17454 ^ n12457;
  assign n17456 = n17455 ^ x276;
  assign n27604 = n27603 ^ n17456;
  assign n39868 = n39867 ^ n27604;
  assign n49915 = n47750 ^ n39868;
  assign n44304 = n42129 ^ n33737;
  assign n38233 = n35953 ^ n27609;
  assign n26201 = n24174 ^ n17461;
  assign n2212 = n2162 ^ n2107;
  assign n2213 = n2212 ^ n2206;
  assign n2214 = n2213 ^ x469;
  assign n26202 = n26201 ^ n2214;
  assign n15977 = n14147 ^ x277;
  assign n15978 = n15977 ^ x469;
  assign n15979 = n15978 ^ x213;
  assign n26203 = n26202 ^ n15979;
  assign n38234 = n38233 ^ n26203;
  assign n2210 = n2174 ^ n2110;
  assign n2202 = n2172 ^ n2102;
  assign n2197 = n2170 ^ n2094;
  assign n2061 = n1973 ^ x279;
  assign n2062 = n2061 ^ x471;
  assign n2063 = n2062 ^ x215;
  assign n2198 = n2197 ^ n2063;
  assign n2199 = n2198 ^ x470;
  assign n2203 = n2202 ^ n2199;
  assign n2207 = n2206 ^ n2203;
  assign n2211 = n2210 ^ n2207;
  assign n2215 = n2214 ^ n2211;
  assign n38235 = n38234 ^ n2215;
  assign n44305 = n44304 ^ n38235;
  assign n31869 = n26203 ^ n22442;
  assign n31870 = n31869 ^ n29646;
  assign n21153 = n19338 ^ n12457;
  assign n21154 = n21153 ^ n15979;
  assign n21155 = n21154 ^ x468;
  assign n31871 = n31870 ^ n21155;
  assign n44306 = n44305 ^ n31871;
  assign n49916 = n49915 ^ n44306;
  assign n38349 = n36040 ^ n27604;
  assign n38350 = n38349 ^ n31871;
  assign n26124 = n24249 ^ n17456;
  assign n26125 = n26124 ^ n21155;
  assign n16040 = n14095 ^ x276;
  assign n16041 = n16040 ^ x468;
  assign n16042 = n16041 ^ x212;
  assign n26126 = n26125 ^ n16042;
  assign n38351 = n38350 ^ n26126;
  assign n49917 = n49916 ^ n38351;
  assign n12818 = x468 ^ x116;
  assign n12819 = n12818 ^ x308;
  assign n12820 = n12819 ^ x52;
  assign n21536 = n19659 ^ n12820;
  assign n16768 = n14731 ^ x308;
  assign n16769 = n16768 ^ x500;
  assign n16770 = n16769 ^ x244;
  assign n21537 = n21536 ^ n16770;
  assign n21538 = n21537 ^ x499;
  assign n31200 = n29314 ^ n21538;
  assign n25707 = n23847 ^ n16770;
  assign n20615 = n18706 ^ x500;
  assign n20616 = n20615 ^ n15599;
  assign n20617 = n20616 ^ x436;
  assign n25708 = n25707 ^ n20617;
  assign n592 = n588 ^ x244;
  assign n593 = n592 ^ x436;
  assign n594 = n593 ^ x180;
  assign n25709 = n25708 ^ n594;
  assign n31201 = n31200 ^ n25709;
  assign n591 = n590 ^ x499;
  assign n595 = n594 ^ n591;
  assign n596 = n595 ^ x435;
  assign n31202 = n31201 ^ n596;
  assign n42122 = n39868 ^ n31202;
  assign n36471 = n33737 ^ n25709;
  assign n29639 = n27609 ^ n20617;
  assign n29640 = n29639 ^ n24249;
  assign n19331 = n17461 ^ x436;
  assign n19332 = n19331 ^ n14095;
  assign n19333 = n19332 ^ x372;
  assign n29641 = n29640 ^ n19333;
  assign n36472 = n36471 ^ n29641;
  assign n24167 = n22442 ^ n594;
  assign n24168 = n24167 ^ n19333;
  assign n14156 = n12457 ^ x180;
  assign n14157 = n14156 ^ x372;
  assign n14158 = n14157 ^ x116;
  assign n24169 = n24168 ^ n14158;
  assign n36473 = n36472 ^ n24169;
  assign n42123 = n42122 ^ n36473;
  assign n29733 = n27604 ^ n596;
  assign n29734 = n29733 ^ n24169;
  assign n19326 = n17456 ^ x435;
  assign n19327 = n19326 ^ n14158;
  assign n19328 = n19327 ^ x371;
  assign n29735 = n29734 ^ n19328;
  assign n42124 = n42123 ^ n29735;
  assign n52027 = n49917 ^ n42124;
  assign n46118 = n44306 ^ n36473;
  assign n40623 = n38235 ^ n29641;
  assign n34716 = n24249 ^ n2215;
  assign n28495 = n19338 ^ n2207;
  assign n23087 = n14147 ^ n2199;
  assign n2154 = n2063 ^ x374;
  assign n2155 = n2154 ^ n578;
  assign n2156 = n2155 ^ x310;
  assign n23088 = n23087 ^ n2156;
  assign n23089 = n23088 ^ n12792;
  assign n28496 = n28495 ^ n23089;
  assign n28497 = n28496 ^ n17818;
  assign n34717 = n34716 ^ n28497;
  assign n23082 = n14095 ^ n2214;
  assign n23083 = n23082 ^ n17818;
  assign n12735 = x469 ^ x117;
  assign n12736 = n12735 ^ x309;
  assign n12737 = n12736 ^ x53;
  assign n23084 = n23083 ^ n12737;
  assign n34718 = n34717 ^ n23084;
  assign n40624 = n40623 ^ n34718;
  assign n28490 = n26203 ^ n19333;
  assign n28491 = n28490 ^ n23084;
  assign n18078 = n15979 ^ x372;
  assign n18079 = n18078 ^ n12737;
  assign n18080 = n18079 ^ x308;
  assign n28492 = n28491 ^ n18080;
  assign n40625 = n40624 ^ n28492;
  assign n46119 = n46118 ^ n40625;
  assign n34711 = n31871 ^ n28492;
  assign n34712 = n34711 ^ n24169;
  assign n23077 = n21155 ^ n14158;
  assign n23078 = n23077 ^ n18080;
  assign n23079 = n23078 ^ n12820;
  assign n34713 = n34712 ^ n23079;
  assign n46120 = n46119 ^ n34713;
  assign n52028 = n52027 ^ n46120;
  assign n40515 = n38351 ^ n29735;
  assign n40516 = n40515 ^ n34713;
  assign n28485 = n26126 ^ n19328;
  assign n28486 = n28485 ^ n23079;
  assign n18073 = n16042 ^ x371;
  assign n18074 = n18073 ^ n12820;
  assign n18075 = n18074 ^ x307;
  assign n28487 = n28486 ^ n18075;
  assign n40517 = n40516 ^ n28487;
  assign n52029 = n52028 ^ n40517;
  assign n14719 = n12820 ^ x211;
  assign n14720 = n14719 ^ x403;
  assign n14721 = n14720 ^ x147;
  assign n23840 = n21538 ^ n14721;
  assign n18697 = n16770 ^ x403;
  assign n13797 = x500 ^ x148;
  assign n13798 = n13797 ^ x340;
  assign n13799 = n13798 ^ x84;
  assign n18698 = n18697 ^ n13799;
  assign n18699 = n18698 ^ x339;
  assign n23841 = n23840 ^ n18699;
  assign n513 = x499 ^ x147;
  assign n514 = n513 ^ x339;
  assign n515 = n514 ^ x83;
  assign n23842 = n23841 ^ n515;
  assign n33637 = n31202 ^ n23842;
  assign n27663 = n25709 ^ n18699;
  assign n22448 = n20617 ^ n13799;
  assign n22449 = n22448 ^ n17456;
  assign n599 = x436 ^ x84;
  assign n600 = n599 ^ x276;
  assign n601 = n600 ^ x20;
  assign n22450 = n22449 ^ n601;
  assign n27664 = n27663 ^ n22450;
  assign n598 = n594 ^ x339;
  assign n602 = n601 ^ n598;
  assign n603 = n602 ^ x275;
  assign n27665 = n27664 ^ n603;
  assign n33638 = n33637 ^ n27665;
  assign n597 = n596 ^ n515;
  assign n604 = n603 ^ n597;
  assign n570 = x435 ^ x83;
  assign n571 = n570 ^ x275;
  assign n572 = n571 ^ x19;
  assign n605 = n604 ^ n572;
  assign n33639 = n33638 ^ n605;
  assign n44294 = n42124 ^ n33639;
  assign n38372 = n36473 ^ n27665;
  assign n31978 = n29641 ^ n22450;
  assign n31979 = n31978 ^ n26126;
  assign n21148 = n19333 ^ n601;
  assign n21149 = n21148 ^ n16042;
  assign n21150 = n21149 ^ x467;
  assign n31980 = n31979 ^ n21150;
  assign n38373 = n38372 ^ n31980;
  assign n26119 = n24169 ^ n603;
  assign n26120 = n26119 ^ n21150;
  assign n15972 = n14158 ^ x275;
  assign n15973 = n15972 ^ x467;
  assign n15974 = n15973 ^ x211;
  assign n26121 = n26120 ^ n15974;
  assign n38374 = n38373 ^ n26121;
  assign n44295 = n44294 ^ n38374;
  assign n32372 = n29735 ^ n605;
  assign n32373 = n32372 ^ n26121;
  assign n21193 = n15974 ^ n572;
  assign n21194 = n21193 ^ n19328;
  assign n21195 = n21194 ^ x466;
  assign n32374 = n32373 ^ n21195;
  assign n44296 = n44295 ^ n32374;
  assign n54145 = n52029 ^ n44296;
  assign n48476 = n46120 ^ n38374;
  assign n42698 = n40625 ^ n31980;
  assign n37173 = n34718 ^ n26126;
  assign n30577 = n28497 ^ n21155;
  assign n24983 = n23089 ^ n15979;
  assign n2259 = n2156 ^ x469;
  assign n2260 = n2259 ^ n581;
  assign n2261 = n2260 ^ x405;
  assign n24984 = n24983 ^ n2261;
  assign n24985 = n24984 ^ n14731;
  assign n30578 = n30577 ^ n24985;
  assign n30579 = n30578 ^ n19659;
  assign n37174 = n37173 ^ n30579;
  assign n24978 = n19659 ^ n16042;
  assign n24979 = n24978 ^ n23084;
  assign n14724 = n12737 ^ x212;
  assign n14725 = n14724 ^ x404;
  assign n14726 = n14725 ^ x148;
  assign n24980 = n24979 ^ n14726;
  assign n37175 = n37174 ^ n24980;
  assign n42699 = n42698 ^ n37175;
  assign n30571 = n28492 ^ n21150;
  assign n30572 = n30571 ^ n24980;
  assign n19745 = n18080 ^ x467;
  assign n19746 = n19745 ^ n14726;
  assign n19747 = n19746 ^ x403;
  assign n30573 = n30572 ^ n19747;
  assign n42700 = n42699 ^ n30573;
  assign n48477 = n48476 ^ n42700;
  assign n37151 = n34713 ^ n26121;
  assign n37152 = n37151 ^ n30573;
  assign n24973 = n23079 ^ n15974;
  assign n24974 = n24973 ^ n19747;
  assign n24975 = n24974 ^ n14721;
  assign n37153 = n37152 ^ n24975;
  assign n48478 = n48477 ^ n37153;
  assign n54146 = n54145 ^ n48478;
  assign n42831 = n40517 ^ n32374;
  assign n42832 = n42831 ^ n37153;
  assign n30566 = n28487 ^ n21195;
  assign n30567 = n30566 ^ n24975;
  assign n19952 = n18075 ^ x466;
  assign n19953 = n19952 ^ n14721;
  assign n19954 = n19953 ^ x402;
  assign n30568 = n30567 ^ n19954;
  assign n42833 = n42832 ^ n30568;
  assign n54147 = n54146 ^ n42833;
  assign n16758 = n14721 ^ x306;
  assign n16759 = n16758 ^ x498;
  assign n16760 = n16759 ^ x242;
  assign n25725 = n23842 ^ n16760;
  assign n20630 = n18699 ^ x498;
  assign n15590 = n13799 ^ x243;
  assign n15591 = n15590 ^ x435;
  assign n15592 = n15591 ^ x179;
  assign n20631 = n20630 ^ n15592;
  assign n20632 = n20631 ^ x434;
  assign n25726 = n25725 ^ n20632;
  assign n516 = n515 ^ x242;
  assign n517 = n516 ^ x434;
  assign n518 = n517 ^ x178;
  assign n25727 = n25726 ^ n518;
  assign n36487 = n33639 ^ n25727;
  assign n29634 = n27665 ^ n20632;
  assign n24162 = n22450 ^ n15592;
  assign n24163 = n24162 ^ n19328;
  assign n608 = n601 ^ x179;
  assign n609 = n608 ^ x371;
  assign n610 = n609 ^ x115;
  assign n24164 = n24163 ^ n610;
  assign n29635 = n29634 ^ n24164;
  assign n607 = n603 ^ x434;
  assign n611 = n610 ^ n607;
  assign n612 = n611 ^ x370;
  assign n29636 = n29635 ^ n612;
  assign n36488 = n36487 ^ n29636;
  assign n606 = n605 ^ n518;
  assign n613 = n612 ^ n606;
  assign n573 = n572 ^ x178;
  assign n574 = n573 ^ x370;
  assign n575 = n574 ^ x114;
  assign n614 = n613 ^ n575;
  assign n36489 = n36488 ^ n614;
  assign n46113 = n44296 ^ n36489;
  assign n40510 = n38374 ^ n29636;
  assign n34706 = n31980 ^ n24164;
  assign n34707 = n34706 ^ n28487;
  assign n23160 = n18075 ^ n610;
  assign n23161 = n23160 ^ n21150;
  assign n12841 = x467 ^ x115;
  assign n12842 = n12841 ^ x307;
  assign n12843 = n12842 ^ x51;
  assign n23162 = n23161 ^ n12843;
  assign n34708 = n34707 ^ n23162;
  assign n40511 = n40510 ^ n34708;
  assign n28480 = n26121 ^ n612;
  assign n28481 = n28480 ^ n23162;
  assign n18068 = n15974 ^ x370;
  assign n18069 = n18068 ^ n12843;
  assign n18070 = n18069 ^ x306;
  assign n28482 = n28481 ^ n18070;
  assign n40512 = n40511 ^ n28482;
  assign n46114 = n46113 ^ n40512;
  assign n23072 = n21195 ^ n575;
  assign n23073 = n23072 ^ n18070;
  assign n630 = x466 ^ x114;
  assign n631 = n630 ^ x306;
  assign n632 = n631 ^ x50;
  assign n23074 = n23073 ^ n632;
  assign n34822 = n32374 ^ n23074;
  assign n34823 = n34822 ^ n28482;
  assign n34824 = n34823 ^ n614;
  assign n46115 = n46114 ^ n34824;
  assign n56234 = n54147 ^ n46115;
  assign n50563 = n48478 ^ n40512;
  assign n45074 = n42700 ^ n34708;
  assign n39166 = n37175 ^ n28487;
  assign n33203 = n30579 ^ n23079;
  assign n26938 = n24985 ^ n18080;
  assign n21541 = n12737 ^ n2261;
  assign n21542 = n21541 ^ n584;
  assign n21543 = n21542 ^ x500;
  assign n26939 = n26938 ^ n21543;
  assign n26940 = n26939 ^ n16770;
  assign n33204 = n33203 ^ n26940;
  assign n33205 = n33204 ^ n21538;
  assign n39167 = n39166 ^ n33205;
  assign n26933 = n24980 ^ n18075;
  assign n26934 = n26933 ^ n21538;
  assign n16763 = n14726 ^ x307;
  assign n16764 = n16763 ^ x499;
  assign n16765 = n16764 ^ x243;
  assign n26935 = n26934 ^ n16765;
  assign n39168 = n39167 ^ n26935;
  assign n45075 = n45074 ^ n39168;
  assign n33198 = n30573 ^ n23162;
  assign n33199 = n33198 ^ n26935;
  assign n21641 = n19747 ^ n12843;
  assign n21642 = n21641 ^ n16765;
  assign n21643 = n21642 ^ x498;
  assign n33200 = n33199 ^ n21643;
  assign n45076 = n45075 ^ n33200;
  assign n50564 = n50563 ^ n45076;
  assign n39161 = n37153 ^ n28482;
  assign n39162 = n39161 ^ n33200;
  assign n27038 = n24975 ^ n18070;
  assign n27039 = n27038 ^ n21643;
  assign n27040 = n27039 ^ n16760;
  assign n39163 = n39162 ^ n27040;
  assign n50565 = n50564 ^ n39163;
  assign n56235 = n56234 ^ n50565;
  assign n45118 = n42833 ^ n34824;
  assign n45119 = n45118 ^ n39163;
  assign n33258 = n30568 ^ n23074;
  assign n33259 = n33258 ^ n27040;
  assign n21857 = n19954 ^ n632;
  assign n21858 = n21857 ^ n16760;
  assign n21859 = n21858 ^ x497;
  assign n33260 = n33259 ^ n21859;
  assign n45120 = n45119 ^ n33260;
  assign n56236 = n56235 ^ n45120;
  assign n2474 = x484 ^ x132;
  assign n2475 = n2474 ^ x324;
  assign n2476 = n2475 ^ x68;
  assign n2549 = n2476 ^ x227;
  assign n2550 = n2549 ^ x419;
  assign n2551 = n2550 ^ x163;
  assign n2630 = n2551 ^ x322;
  assign n2631 = n2630 ^ n2538;
  assign n2632 = n2631 ^ x258;
  assign n2312 = x454 ^ x102;
  assign n2313 = n2312 ^ x38;
  assign n2314 = n2313 ^ x294;
  assign n2354 = n2314 ^ x197;
  assign n2355 = n2354 ^ x389;
  assign n2356 = n2355 ^ x133;
  assign n2407 = n2356 ^ x292;
  assign n2408 = n2407 ^ x484;
  assign n2409 = n2408 ^ x228;
  assign n2473 = n2409 ^ x387;
  assign n2477 = n2476 ^ n2473;
  assign n2478 = n2477 ^ x323;
  assign n2548 = n2478 ^ x482;
  assign n2552 = n2551 ^ n2548;
  assign n2553 = n2552 ^ x418;
  assign n1495 = x482 ^ x130;
  assign n1496 = n1495 ^ x322;
  assign n1497 = n1496 ^ x66;
  assign n2629 = n2553 ^ n1497;
  assign n2633 = n2632 ^ n2629;
  assign n2623 = x418 ^ x66;
  assign n2624 = n2623 ^ x258;
  assign n2625 = n2624 ^ x2;
  assign n2634 = n2633 ^ n2625;
  assign n1211 = x424 ^ x72;
  assign n1212 = n1211 ^ x264;
  assign n1213 = n1212 ^ x8;
  assign n1313 = n1213 ^ x167;
  assign n1314 = n1313 ^ x359;
  assign n1315 = n1314 ^ x103;
  assign n2279 = n1315 ^ x262;
  assign n2280 = n2279 ^ x454;
  assign n2281 = n2280 ^ x198;
  assign n2321 = n2281 ^ x357;
  assign n2322 = n2321 ^ n2314;
  assign n2323 = n2322 ^ x293;
  assign n2366 = n2323 ^ x452;
  assign n2367 = n2366 ^ n2356;
  assign n2368 = n2367 ^ x388;
  assign n1509 = x452 ^ x36;
  assign n1510 = n1509 ^ x100;
  assign n1511 = n1510 ^ x292;
  assign n2406 = n2368 ^ n1511;
  assign n2410 = n2409 ^ n2406;
  assign n2411 = n2410 ^ x483;
  assign n1512 = n1511 ^ x195;
  assign n1513 = n1512 ^ x387;
  assign n1514 = n1513 ^ x131;
  assign n2472 = n2411 ^ n1514;
  assign n2479 = n2478 ^ n2472;
  assign n2469 = x483 ^ x131;
  assign n2470 = n2469 ^ x323;
  assign n2471 = n2470 ^ x67;
  assign n2480 = n2479 ^ n2471;
  assign n1515 = n1514 ^ x290;
  assign n1516 = n1515 ^ x482;
  assign n1517 = n1516 ^ x226;
  assign n2547 = n2480 ^ n1517;
  assign n2554 = n2553 ^ n2547;
  assign n2544 = n2471 ^ x226;
  assign n2545 = n2544 ^ x418;
  assign n2546 = n2545 ^ x162;
  assign n2555 = n2554 ^ n2546;
  assign n1518 = n1517 ^ x385;
  assign n1519 = n1518 ^ n1497;
  assign n1520 = n1519 ^ x321;
  assign n2628 = n2555 ^ n1520;
  assign n2635 = n2634 ^ n2628;
  assign n2622 = n2546 ^ x321;
  assign n2626 = n2625 ^ n2622;
  assign n2627 = n2626 ^ x257;
  assign n2636 = n2635 ^ n2627;
  assign n1333 = x455 ^ x39;
  assign n1334 = n1333 ^ x295;
  assign n1335 = n1334 ^ x103;
  assign n2292 = n1335 ^ x198;
  assign n2293 = n2292 ^ x390;
  assign n2294 = n2293 ^ x134;
  assign n2341 = n2294 ^ x293;
  assign n2342 = n2341 ^ x485;
  assign n2343 = n2342 ^ x229;
  assign n2399 = n2343 ^ x388;
  assign n2393 = x485 ^ x133;
  assign n2394 = n2393 ^ x325;
  assign n2395 = n2394 ^ x69;
  assign n2400 = n2399 ^ n2395;
  assign n2401 = n2400 ^ x324;
  assign n2464 = n2401 ^ x483;
  assign n2443 = n2395 ^ x228;
  assign n2444 = n2443 ^ x420;
  assign n2445 = n2444 ^ x164;
  assign n2465 = n2464 ^ n2445;
  assign n2466 = n2465 ^ x419;
  assign n889 = x491 ^ x139;
  assign n890 = n889 ^ x331;
  assign n891 = n890 ^ x75;
  assign n953 = n891 ^ x234;
  assign n954 = n953 ^ x426;
  assign n955 = n954 ^ x170;
  assign n1040 = n955 ^ x329;
  assign n1035 = x426 ^ x74;
  assign n1036 = n1035 ^ x266;
  assign n1037 = n1036 ^ x10;
  assign n1041 = n1040 ^ n1037;
  assign n1042 = n1041 ^ x265;
  assign n1127 = n1042 ^ x424;
  assign n1122 = n1037 ^ x169;
  assign n1123 = n1122 ^ x361;
  assign n1124 = n1123 ^ x105;
  assign n1128 = n1127 ^ n1124;
  assign n1129 = n1128 ^ x360;
  assign n1226 = n1213 ^ n1129;
  assign n1221 = n1124 ^ x264;
  assign n1222 = n1221 ^ x456;
  assign n1223 = n1222 ^ x200;
  assign n1227 = n1226 ^ n1223;
  assign n1228 = n1227 ^ x455;
  assign n1331 = n1315 ^ n1228;
  assign n1326 = n1223 ^ x359;
  assign n1321 = x456 ^ x104;
  assign n1322 = n1321 ^ x296;
  assign n1323 = n1322 ^ x40;
  assign n1327 = n1326 ^ n1323;
  assign n1328 = n1327 ^ x295;
  assign n1332 = n1331 ^ n1328;
  assign n1336 = n1335 ^ n1332;
  assign n2290 = n2281 ^ n1336;
  assign n2287 = n1328 ^ x454;
  assign n2284 = n1323 ^ x199;
  assign n2285 = n2284 ^ x391;
  assign n2286 = n2285 ^ x135;
  assign n2288 = n2287 ^ n2286;
  assign n2289 = n2288 ^ x390;
  assign n2291 = n2290 ^ n2289;
  assign n2295 = n2294 ^ n2291;
  assign n2339 = n2323 ^ n2295;
  assign n2334 = n2314 ^ n2289;
  assign n2329 = n2286 ^ x294;
  assign n2330 = n2329 ^ x486;
  assign n2331 = n2330 ^ x230;
  assign n2335 = n2334 ^ n2331;
  assign n2336 = n2335 ^ x485;
  assign n2340 = n2339 ^ n2336;
  assign n2344 = n2343 ^ n2340;
  assign n2402 = n2368 ^ n2344;
  assign n2391 = n2356 ^ n2336;
  assign n2386 = n2331 ^ x389;
  assign n2381 = x486 ^ x134;
  assign n2382 = n2381 ^ x326;
  assign n2383 = n2382 ^ x70;
  assign n2387 = n2386 ^ n2383;
  assign n2388 = n2387 ^ x325;
  assign n2392 = n2391 ^ n2388;
  assign n2396 = n2395 ^ n2392;
  assign n2403 = n2402 ^ n2396;
  assign n2404 = n2403 ^ n2401;
  assign n2462 = n2411 ^ n2404;
  assign n2441 = n2409 ^ n2396;
  assign n2438 = n2388 ^ x484;
  assign n2435 = n2383 ^ x229;
  assign n2436 = n2435 ^ x421;
  assign n2437 = n2436 ^ x165;
  assign n2439 = n2438 ^ n2437;
  assign n2440 = n2439 ^ x420;
  assign n2442 = n2441 ^ n2440;
  assign n2446 = n2445 ^ n2442;
  assign n2463 = n2462 ^ n2446;
  assign n2467 = n2466 ^ n2463;
  assign n2540 = n2480 ^ n2467;
  assign n2528 = n2445 ^ x323;
  assign n2520 = x420 ^ x68;
  assign n2521 = n2520 ^ x260;
  assign n2522 = n2521 ^ x4;
  assign n2529 = n2528 ^ n2522;
  assign n2530 = n2529 ^ x259;
  assign n2526 = n2478 ^ n2446;
  assign n2518 = n2476 ^ n2440;
  assign n2513 = n2437 ^ x324;
  assign n2358 = x421 ^ x69;
  assign n2359 = n2358 ^ x261;
  assign n2360 = n2359 ^ x5;
  assign n2514 = n2513 ^ n2360;
  assign n2515 = n2514 ^ x260;
  assign n2519 = n2518 ^ n2515;
  assign n2523 = n2522 ^ n2519;
  assign n2527 = n2526 ^ n2523;
  assign n2531 = n2530 ^ n2527;
  assign n2541 = n2540 ^ n2531;
  assign n2534 = n2471 ^ n2466;
  assign n2535 = n2534 ^ n2530;
  assign n2539 = n2538 ^ n2535;
  assign n2542 = n2541 ^ n2539;
  assign n2618 = n2555 ^ n2542;
  assign n2606 = n2530 ^ x418;
  assign n2587 = n2522 ^ x163;
  assign n2588 = n2587 ^ x355;
  assign n2589 = n2588 ^ x99;
  assign n2607 = n2606 ^ n2589;
  assign n2608 = n2607 ^ x354;
  assign n2604 = n2553 ^ n2531;
  assign n2585 = n2551 ^ n2523;
  assign n2582 = n2515 ^ x419;
  assign n2424 = n2360 ^ x164;
  assign n2425 = n2424 ^ x356;
  assign n2426 = n2425 ^ x100;
  assign n2583 = n2582 ^ n2426;
  assign n2584 = n2583 ^ x355;
  assign n2586 = n2585 ^ n2584;
  assign n2590 = n2589 ^ n2586;
  assign n2605 = n2604 ^ n2590;
  assign n2609 = n2608 ^ n2605;
  assign n2619 = n2618 ^ n2609;
  assign n2612 = n2546 ^ n2539;
  assign n2613 = n2612 ^ n2608;
  assign n2617 = n2616 ^ n2613;
  assign n2620 = n2619 ^ n2617;
  assign n38275 = n2636 ^ n2620;
  assign n25795 = n2627 ^ n2617;
  assign n21368 = n2625 ^ n2608;
  assign n16337 = n2589 ^ x258;
  assign n16338 = n16337 ^ x450;
  assign n16339 = n16338 ^ x194;
  assign n21369 = n21368 ^ n16339;
  assign n21370 = n21369 ^ x449;
  assign n25796 = n25795 ^ n21370;
  assign n25797 = n25796 ^ n16401;
  assign n38276 = n38275 ^ n25797;
  assign n26588 = n2632 ^ n2590;
  assign n21355 = n2584 ^ n2538;
  assign n2487 = n2426 ^ x259;
  assign n2488 = n2487 ^ x451;
  assign n2489 = n2488 ^ x195;
  assign n21356 = n21355 ^ n2489;
  assign n21357 = n21356 ^ x450;
  assign n26589 = n26588 ^ n21357;
  assign n26590 = n26589 ^ n16339;
  assign n31912 = n26590 ^ n2609;
  assign n31913 = n31912 ^ n2634;
  assign n31914 = n31913 ^ n21370;
  assign n38277 = n38276 ^ n31914;
  assign n1494 = x417 ^ x225;
  assign n1498 = n1497 ^ n1494;
  assign n1499 = n1498 ^ x161;
  assign n24200 = n2634 ^ n1499;
  assign n19477 = n2632 ^ x417;
  assign n19478 = n19477 ^ n2616;
  assign n19479 = n19478 ^ x353;
  assign n24201 = n24200 ^ n19479;
  assign n14515 = n2625 ^ x161;
  assign n14516 = n14515 ^ x353;
  assign n14517 = n14516 ^ x97;
  assign n24202 = n24201 ^ n14517;
  assign n34770 = n31914 ^ n24202;
  assign n28518 = n26590 ^ n19479;
  assign n23278 = n21357 ^ n2616;
  assign n2557 = x451 ^ x99;
  assign n2558 = n2557 ^ x291;
  assign n2559 = n2558 ^ x35;
  assign n2556 = n2489 ^ x354;
  assign n2560 = n2559 ^ n2556;
  assign n2561 = n2560 ^ x290;
  assign n23279 = n23278 ^ n2561;
  assign n1422 = x450 ^ x98;
  assign n1423 = n1422 ^ x290;
  assign n1424 = n1423 ^ x34;
  assign n23280 = n23279 ^ n1424;
  assign n28519 = n28518 ^ n23280;
  assign n18237 = n16339 ^ x353;
  assign n18238 = n18237 ^ n1424;
  assign n18239 = n18238 ^ x289;
  assign n28520 = n28519 ^ n18239;
  assign n34771 = n34770 ^ n28520;
  assign n22535 = n21370 ^ n14517;
  assign n22536 = n22535 ^ n18239;
  assign n22537 = n22536 ^ n13254;
  assign n34772 = n34771 ^ n22537;
  assign n40556 = n38277 ^ n34772;
  assign n1521 = n1520 ^ x480;
  assign n1522 = n1521 ^ n1499;
  assign n1523 = n1522 ^ x416;
  assign n29677 = n2636 ^ n1523;
  assign n29678 = n29677 ^ n24202;
  assign n18849 = n2627 ^ x416;
  assign n18850 = n18849 ^ n14517;
  assign n18851 = n18850 ^ x352;
  assign n29679 = n29678 ^ n18851;
  assign n40557 = n40556 ^ n29679;
  assign n28523 = n25797 ^ n18851;
  assign n28524 = n28523 ^ n22537;
  assign n28525 = n28524 ^ n17764;
  assign n40558 = n40557 ^ n28525;
  assign n1410 = x480 ^ x128;
  assign n1411 = n1410 ^ x64;
  assign n1412 = n1411 ^ x320;
  assign n1524 = n1523 ^ n1412;
  assign n1500 = n1499 ^ x320;
  assign n1485 = x417 ^ x65;
  assign n1486 = n1485 ^ x257;
  assign n1487 = n1486 ^ x1;
  assign n1501 = n1500 ^ n1487;
  assign n1502 = n1501 ^ x256;
  assign n1525 = n1524 ^ n1502;
  assign n1468 = x416 ^ x64;
  assign n1469 = n1468 ^ x256;
  assign n1470 = n1469 ^ x0;
  assign n1526 = n1525 ^ n1470;
  assign n31908 = n29679 ^ n1526;
  assign n26152 = n24202 ^ n1502;
  assign n20790 = n19479 ^ n1487;
  assign n20791 = n20790 ^ n16401;
  assign n20792 = n20791 ^ x448;
  assign n26153 = n26152 ^ n20792;
  assign n15993 = n14517 ^ x256;
  assign n15994 = n15993 ^ x448;
  assign n15995 = n15994 ^ x192;
  assign n26154 = n26153 ^ n15995;
  assign n31909 = n31908 ^ n26154;
  assign n20794 = n18851 ^ n1470;
  assign n20795 = n20794 ^ n15995;
  assign n20796 = n20795 ^ x479;
  assign n31910 = n31909 ^ n20796;
  assign n42737 = n40558 ^ n31910;
  assign n25012 = n22537 ^ n15995;
  assign n19678 = n18239 ^ x448;
  assign n1425 = n1424 ^ x193;
  assign n1426 = n1425 ^ x385;
  assign n1427 = n1426 ^ x129;
  assign n19679 = n19678 ^ n1427;
  assign n19680 = n19679 ^ x384;
  assign n25013 = n25012 ^ n19680;
  assign n25014 = n25013 ^ n14747;
  assign n36709 = n34772 ^ n25014;
  assign n36710 = n36709 ^ n26154;
  assign n30624 = n28520 ^ n20792;
  assign n25008 = n23280 ^ n16401;
  assign n20095 = n2561 ^ x449;
  assign n2637 = n2559 ^ x194;
  assign n2638 = n2637 ^ x386;
  assign n2639 = n2638 ^ x130;
  assign n20096 = n20095 ^ n2639;
  assign n20097 = n20096 ^ x385;
  assign n25009 = n25008 ^ n20097;
  assign n25010 = n25009 ^ n1427;
  assign n30625 = n30624 ^ n25010;
  assign n30626 = n30625 ^ n19680;
  assign n36711 = n36710 ^ n30626;
  assign n42738 = n42737 ^ n36711;
  assign n30632 = n28525 ^ n20796;
  assign n30633 = n30632 ^ n25014;
  assign n30634 = n30633 ^ n19684;
  assign n42739 = n42738 ^ n30634;
  assign n1413 = n1412 ^ x255;
  assign n1414 = n1413 ^ x447;
  assign n1415 = n1414 ^ x191;
  assign n1527 = n1526 ^ n1415;
  assign n1503 = n1502 ^ x447;
  assign n1488 = n1487 ^ x160;
  assign n1489 = n1488 ^ x352;
  assign n1490 = n1489 ^ x96;
  assign n1504 = n1503 ^ n1490;
  assign n1505 = n1504 ^ x383;
  assign n1528 = n1527 ^ n1505;
  assign n1474 = n1470 ^ x191;
  assign n1475 = n1474 ^ x383;
  assign n1476 = n1475 ^ x127;
  assign n1529 = n1528 ^ n1476;
  assign n34756 = n31910 ^ n1529;
  assign n28532 = n26154 ^ n1505;
  assign n23106 = n20792 ^ n1490;
  assign n23107 = n23106 ^ n17764;
  assign n12751 = x448 ^ x96;
  assign n12752 = n12751 ^ x288;
  assign n12753 = n12752 ^ x32;
  assign n23108 = n23107 ^ n12753;
  assign n28533 = n28532 ^ n23108;
  assign n17759 = n15995 ^ x383;
  assign n17760 = n17759 ^ n12753;
  assign n17761 = n17760 ^ x319;
  assign n28534 = n28533 ^ n17761;
  assign n34757 = n34756 ^ n28534;
  assign n23117 = n20796 ^ n1476;
  assign n23118 = n23117 ^ n17761;
  assign n23119 = n23118 ^ n1572;
  assign n34758 = n34757 ^ n23119;
  assign n44658 = n42739 ^ n34758;
  assign n32689 = n30626 ^ n23108;
  assign n26969 = n25010 ^ n17764;
  assign n21566 = n20097 ^ n13254;
  assign n2640 = n2639 ^ x289;
  assign n2641 = n2640 ^ x481;
  assign n2642 = n2641 ^ x225;
  assign n21567 = n21566 ^ n2642;
  assign n21568 = n21567 ^ x480;
  assign n26970 = n26969 ^ n21568;
  assign n1428 = n1427 ^ x288;
  assign n1429 = n1428 ^ x480;
  assign n1430 = n1429 ^ x224;
  assign n26971 = n26970 ^ n1430;
  assign n32690 = n32689 ^ n26971;
  assign n21570 = n19680 ^ x511;
  assign n21571 = n21570 ^ n1430;
  assign n21572 = n21571 ^ n12753;
  assign n32691 = n32690 ^ n21572;
  assign n39234 = n32691 ^ n28534;
  assign n39235 = n39234 ^ n36711;
  assign n26961 = n25014 ^ n17761;
  assign n26962 = n26961 ^ n21572;
  assign n26963 = n26962 ^ n16789;
  assign n39236 = n39235 ^ n26963;
  assign n44659 = n44658 ^ n39236;
  assign n32685 = n30634 ^ n23119;
  assign n32686 = n32685 ^ n26963;
  assign n32687 = n32686 ^ n21564;
  assign n44660 = n44659 ^ n32687;
  assign n1417 = x447 ^ x95;
  assign n1418 = n1417 ^ x287;
  assign n1419 = n1418 ^ x31;
  assign n1416 = n1415 ^ x350;
  assign n1420 = n1419 ^ n1416;
  assign n1421 = n1420 ^ x286;
  assign n1530 = n1529 ^ n1421;
  assign n1506 = n1505 ^ n1419;
  assign n1491 = n1490 ^ x287;
  assign n1492 = n1491 ^ x479;
  assign n1493 = n1492 ^ x223;
  assign n1507 = n1506 ^ n1493;
  assign n1508 = n1507 ^ x478;
  assign n1531 = n1530 ^ n1508;
  assign n1480 = n1476 ^ x286;
  assign n1481 = n1480 ^ x478;
  assign n1482 = n1481 ^ x222;
  assign n1532 = n1531 ^ n1482;
  assign n36704 = n34758 ^ n1532;
  assign n30641 = n28534 ^ n1508;
  assign n25003 = n23108 ^ n1493;
  assign n25004 = n25003 ^ n19684;
  assign n14749 = n12753 ^ x223;
  assign n14750 = n14749 ^ x415;
  assign n14751 = n14750 ^ x159;
  assign n25005 = n25004 ^ n14751;
  assign n30642 = n30641 ^ n25005;
  assign n19673 = n17761 ^ x478;
  assign n19674 = n19673 ^ n14751;
  assign n19675 = n19674 ^ x414;
  assign n30643 = n30642 ^ n19675;
  assign n36705 = n36704 ^ n30643;
  assign n24998 = n23119 ^ n1482;
  assign n24999 = n24998 ^ n19675;
  assign n25000 = n24999 ^ n1607;
  assign n36706 = n36705 ^ n25000;
  assign n47027 = n44660 ^ n36706;
  assign n41452 = n39236 ^ n30643;
  assign n35059 = n32691 ^ n25005;
  assign n28805 = n26971 ^ n19684;
  assign n23395 = n21568 ^ n14747;
  assign n18357 = n2642 ^ x384;
  assign n1461 = x481 ^ x129;
  assign n1462 = n1461 ^ x321;
  assign n1463 = n1462 ^ x65;
  assign n18358 = n18357 ^ n1463;
  assign n18359 = n18358 ^ x320;
  assign n23396 = n23395 ^ n18359;
  assign n23397 = n23396 ^ n1412;
  assign n28806 = n28805 ^ n23397;
  assign n1431 = n1430 ^ x415;
  assign n1432 = n1431 ^ n1412;
  assign n1433 = n1432 ^ x351;
  assign n28807 = n28806 ^ n1433;
  assign n35060 = n35059 ^ n28807;
  assign n23403 = n21572 ^ n14751;
  assign n23404 = n23403 ^ n1433;
  assign n23405 = n23404 ^ n13343;
  assign n35061 = n35060 ^ n23405;
  assign n41453 = n41452 ^ n35061;
  assign n28801 = n26963 ^ n19675;
  assign n28802 = n28801 ^ n23405;
  assign n28803 = n28802 ^ n18370;
  assign n41454 = n41453 ^ n28803;
  assign n47028 = n47027 ^ n41454;
  assign n35054 = n32687 ^ n25000;
  assign n35055 = n35054 ^ n28803;
  assign n35056 = n35055 ^ n23392;
  assign n47029 = n47028 ^ n35056;
  assign n1581 = n1482 ^ x381;
  assign n1576 = x478 ^ x126;
  assign n1577 = n1576 ^ x318;
  assign n1578 = n1577 ^ x62;
  assign n1582 = n1581 ^ n1578;
  assign n1583 = n1582 ^ x317;
  assign n1569 = n1493 ^ x382;
  assign n1573 = n1572 ^ n1569;
  assign n1574 = n1573 ^ x318;
  assign n1451 = n1419 ^ x190;
  assign n1452 = n1451 ^ x382;
  assign n1453 = n1452 ^ x126;
  assign n1568 = n1508 ^ n1453;
  assign n1575 = n1574 ^ n1568;
  assign n1579 = n1578 ^ n1575;
  assign n1450 = n1421 ^ x445;
  assign n1454 = n1453 ^ n1450;
  assign n1455 = n1454 ^ x381;
  assign n1567 = n1532 ^ n1455;
  assign n1580 = n1579 ^ n1567;
  assign n1584 = n1583 ^ n1580;
  assign n39202 = n36706 ^ n1584;
  assign n32673 = n30643 ^ n1579;
  assign n26957 = n25005 ^ n1574;
  assign n26958 = n26957 ^ n21564;
  assign n16795 = n14751 ^ x318;
  assign n16796 = n16795 ^ x510;
  assign n16797 = n16796 ^ x254;
  assign n26959 = n26958 ^ n16797;
  assign n32674 = n32673 ^ n26959;
  assign n21556 = n19675 ^ n1578;
  assign n21557 = n21556 ^ n16797;
  assign n21558 = n21557 ^ x509;
  assign n32675 = n32674 ^ n21558;
  assign n39203 = n39202 ^ n32675;
  assign n26987 = n25000 ^ n1583;
  assign n26988 = n26987 ^ n21558;
  assign n26989 = n26988 ^ n1665;
  assign n39204 = n39203 ^ n26989;
  assign n49243 = n47029 ^ n39204;
  assign n43614 = n41454 ^ n32675;
  assign n37362 = n35061 ^ n26959;
  assign n31243 = n28807 ^ n21564;
  assign n25179 = n23397 ^ n16789;
  assign n20251 = n18359 ^ x511;
  assign n1464 = n1463 ^ x224;
  assign n1465 = n1464 ^ x416;
  assign n1466 = n1465 ^ x160;
  assign n20252 = n20251 ^ n1466;
  assign n20253 = n20252 ^ x447;
  assign n25180 = n25179 ^ n20253;
  assign n25181 = n25180 ^ n1415;
  assign n31244 = n31243 ^ n25181;
  assign n1434 = n1433 ^ x510;
  assign n1435 = n1434 ^ n1415;
  assign n1436 = n1435 ^ x446;
  assign n31245 = n31244 ^ n1436;
  assign n37363 = n37362 ^ n31245;
  assign n25649 = n23405 ^ n16797;
  assign n25650 = n25649 ^ n1436;
  assign n25651 = n25650 ^ n15255;
  assign n37364 = n37363 ^ n25651;
  assign n43615 = n43614 ^ n37364;
  assign n31238 = n28803 ^ n21558;
  assign n31239 = n31238 ^ n25651;
  assign n31240 = n31239 ^ n20266;
  assign n43616 = n43615 ^ n31240;
  assign n49244 = n49243 ^ n43616;
  assign n37357 = n35056 ^ n26989;
  assign n37358 = n37357 ^ n31240;
  assign n37359 = n37358 ^ n25646;
  assign n49245 = n49244 ^ n37359;
  assign n1616 = n1583 ^ x476;
  assign n1611 = n1578 ^ x221;
  assign n1612 = n1611 ^ x413;
  assign n1613 = n1612 ^ x157;
  assign n1617 = n1616 ^ n1613;
  assign n1618 = n1617 ^ x412;
  assign n1604 = n1574 ^ x477;
  assign n1608 = n1607 ^ n1604;
  assign n1609 = n1608 ^ x413;
  assign n1597 = n1453 ^ x285;
  assign n1598 = n1597 ^ x477;
  assign n1599 = n1598 ^ x221;
  assign n1603 = n1599 ^ n1579;
  assign n1610 = n1609 ^ n1603;
  assign n1614 = n1613 ^ n1610;
  assign n1596 = n1595 ^ n1455;
  assign n1600 = n1599 ^ n1596;
  assign n1601 = n1600 ^ x476;
  assign n1602 = n1601 ^ n1584;
  assign n1615 = n1614 ^ n1602;
  assign n1619 = n1618 ^ n1615;
  assign n41441 = n39204 ^ n1619;
  assign n35089 = n32675 ^ n1614;
  assign n28797 = n26959 ^ n1609;
  assign n28798 = n28797 ^ n23392;
  assign n18353 = n16797 ^ x413;
  assign n18354 = n18353 ^ n1439;
  assign n18355 = n18354 ^ x349;
  assign n28799 = n28798 ^ n18355;
  assign n35090 = n35089 ^ n28799;
  assign n23384 = n21558 ^ n1613;
  assign n23385 = n23384 ^ n18355;
  assign n23386 = n23385 ^ n1717;
  assign n35091 = n35090 ^ n23386;
  assign n41442 = n41441 ^ n35091;
  assign n28792 = n26989 ^ n1618;
  assign n28793 = n28792 ^ n23386;
  assign n28794 = n28793 ^ n1719;
  assign n41443 = n41442 ^ n28794;
  assign n51288 = n49245 ^ n41443;
  assign n45534 = n43616 ^ n35091;
  assign n39900 = n37364 ^ n28799;
  assign n33676 = n31245 ^ n23392;
  assign n27195 = n25181 ^ n18370;
  assign n22386 = n20253 ^ n13343;
  assign n1467 = n1466 ^ x351;
  assign n1471 = n1470 ^ n1467;
  assign n1472 = n1471 ^ x287;
  assign n22387 = n22386 ^ n1472;
  assign n22388 = n22387 ^ n1419;
  assign n27196 = n27195 ^ n22388;
  assign n27197 = n27196 ^ n1421;
  assign n33677 = n33676 ^ n27197;
  assign n1440 = n1439 ^ n1436;
  assign n1441 = n1440 ^ n1421;
  assign n1445 = n1444 ^ n1441;
  assign n33678 = n33677 ^ n1445;
  assign n39901 = n39900 ^ n33678;
  assign n27282 = n25651 ^ n18355;
  assign n27283 = n27282 ^ n1445;
  assign n27284 = n27283 ^ n17478;
  assign n39902 = n39901 ^ n27284;
  assign n45535 = n45534 ^ n39902;
  assign n33671 = n31240 ^ n23386;
  assign n33672 = n33671 ^ n27284;
  assign n33673 = n33672 ^ n22381;
  assign n45536 = n45535 ^ n33673;
  assign n51289 = n51288 ^ n45536;
  assign n39895 = n37359 ^ n28794;
  assign n39896 = n39895 ^ n33673;
  assign n39897 = n39896 ^ n27625;
  assign n51290 = n51289 ^ n39897;
  assign n1674 = n1652 ^ n1618;
  assign n1669 = n1613 ^ x316;
  assign n1670 = n1669 ^ x508;
  assign n1671 = n1670 ^ x252;
  assign n1675 = n1674 ^ n1671;
  assign n1676 = n1675 ^ x507;
  assign n1588 = x477 ^ x125;
  assign n1589 = n1588 ^ x317;
  assign n1590 = n1589 ^ x61;
  assign n1662 = n1609 ^ n1590;
  assign n1666 = n1665 ^ n1662;
  assign n1667 = n1666 ^ x508;
  assign n1646 = n1599 ^ x380;
  assign n1647 = n1646 ^ n1590;
  assign n1648 = n1647 ^ x316;
  assign n1661 = n1648 ^ n1614;
  assign n1668 = n1667 ^ n1661;
  assign n1672 = n1671 ^ n1668;
  assign n1645 = n1640 ^ n1601;
  assign n1649 = n1648 ^ n1645;
  assign n1653 = n1652 ^ n1649;
  assign n1660 = n1653 ^ n1619;
  assign n1673 = n1672 ^ n1660;
  assign n1677 = n1676 ^ n1673;
  assign n43625 = n41443 ^ n1677;
  assign n37397 = n35091 ^ n1672;
  assign n31232 = n28799 ^ n1667;
  assign n31233 = n31232 ^ n25646;
  assign n20243 = n18355 ^ x508;
  assign n20244 = n20243 ^ n1448;
  assign n20245 = n20244 ^ x444;
  assign n31234 = n31233 ^ n20245;
  assign n37398 = n37397 ^ n31234;
  assign n25664 = n23386 ^ n1671;
  assign n25665 = n25664 ^ n20245;
  assign n25666 = n25665 ^ n1783;
  assign n37399 = n37398 ^ n25666;
  assign n43626 = n43625 ^ n37399;
  assign n31227 = n28794 ^ n1676;
  assign n31228 = n31227 ^ n25666;
  assign n31229 = n31228 ^ n1785;
  assign n43627 = n43626 ^ n31229;
  assign n53399 = n51290 ^ n43627;
  assign n47773 = n45536 ^ n37399;
  assign n42149 = n39902 ^ n31234;
  assign n35977 = n33678 ^ n25646;
  assign n29664 = n27197 ^ n20266;
  assign n24193 = n22388 ^ n15255;
  assign n1473 = n1472 ^ x446;
  assign n1477 = n1476 ^ n1473;
  assign n1478 = n1477 ^ x382;
  assign n24194 = n24193 ^ n1478;
  assign n24195 = n24194 ^ n1453;
  assign n29665 = n29664 ^ n24195;
  assign n29666 = n29665 ^ n1455;
  assign n35978 = n35977 ^ n29666;
  assign n1449 = n1448 ^ n1445;
  assign n1456 = n1455 ^ n1449;
  assign n1460 = n1459 ^ n1456;
  assign n35979 = n35978 ^ n1460;
  assign n42150 = n42149 ^ n35979;
  assign n29660 = n27284 ^ n20245;
  assign n29661 = n29660 ^ n1460;
  assign n29662 = n29661 ^ n19351;
  assign n42151 = n42150 ^ n29662;
  assign n47774 = n47773 ^ n42151;
  assign n35972 = n33673 ^ n25666;
  assign n35973 = n35972 ^ n29662;
  assign n35974 = n35973 ^ n24188;
  assign n47775 = n47774 ^ n35974;
  assign n53400 = n53399 ^ n47775;
  assign n42144 = n39897 ^ n31229;
  assign n42145 = n42144 ^ n35974;
  assign n42146 = n42145 ^ n29704;
  assign n53401 = n53400 ^ n42146;
  assign n1731 = n1703 ^ n1676;
  assign n1726 = n1671 ^ x411;
  assign n1721 = x508 ^ x156;
  assign n1722 = n1721 ^ x348;
  assign n1723 = n1722 ^ x92;
  assign n1727 = n1726 ^ n1723;
  assign n1728 = n1727 ^ x347;
  assign n1732 = n1731 ^ n1728;
  assign n1736 = n1735 ^ n1732;
  assign n1633 = n1590 ^ x220;
  assign n1634 = n1633 ^ x412;
  assign n1635 = n1634 ^ x156;
  assign n1713 = n1667 ^ n1635;
  assign n1720 = n1719 ^ n1713;
  assign n1724 = n1723 ^ n1720;
  assign n1697 = n1648 ^ x475;
  assign n1698 = n1697 ^ n1635;
  assign n1699 = n1698 ^ x411;
  assign n1712 = n1699 ^ n1672;
  assign n1725 = n1724 ^ n1712;
  assign n1729 = n1728 ^ n1725;
  assign n1696 = n1688 ^ n1653;
  assign n1700 = n1699 ^ n1696;
  assign n1704 = n1703 ^ n1700;
  assign n1711 = n1704 ^ n1677;
  assign n1730 = n1729 ^ n1711;
  assign n1737 = n1736 ^ n1730;
  assign n45523 = n43627 ^ n1737;
  assign n39889 = n37399 ^ n1729;
  assign n33665 = n31234 ^ n1724;
  assign n33666 = n33665 ^ n27625;
  assign n22410 = n20245 ^ n1723;
  assign n22411 = n22410 ^ n1623;
  assign n22412 = n22411 ^ n1855;
  assign n33667 = n33666 ^ n22412;
  assign n39890 = n39889 ^ n33667;
  assign n27617 = n25666 ^ n1728;
  assign n27618 = n27617 ^ n22412;
  assign n27619 = n27618 ^ n1858;
  assign n39891 = n39890 ^ n27619;
  assign n45524 = n45523 ^ n39891;
  assign n33660 = n31229 ^ n1736;
  assign n33661 = n33660 ^ n27619;
  assign n33662 = n33661 ^ n1860;
  assign n45525 = n45524 ^ n33662;
  assign n55322 = n53401 ^ n45525;
  assign n49526 = n47775 ^ n39891;
  assign n44372 = n42151 ^ n33667;
  assign n38252 = n35979 ^ n27625;
  assign n31896 = n29666 ^ n22381;
  assign n26147 = n24195 ^ n17478;
  assign n1479 = n1478 ^ n1444;
  assign n1483 = n1482 ^ n1479;
  assign n1484 = n1483 ^ x477;
  assign n26148 = n26147 ^ n1484;
  assign n26149 = n26148 ^ n1599;
  assign n31897 = n31896 ^ n26149;
  assign n31898 = n31897 ^ n1601;
  assign n38253 = n38252 ^ n31898;
  assign n1624 = n1623 ^ n1460;
  assign n1625 = n1624 ^ n1601;
  assign n1629 = n1628 ^ n1625;
  assign n38254 = n38253 ^ n1629;
  assign n44373 = n44372 ^ n38254;
  assign n31892 = n29662 ^ n22412;
  assign n31893 = n31892 ^ n1629;
  assign n31894 = n31893 ^ n20829;
  assign n44374 = n44373 ^ n31894;
  assign n49527 = n49526 ^ n44374;
  assign n38247 = n35974 ^ n27619;
  assign n38248 = n38247 ^ n31894;
  assign n38249 = n38248 ^ n26142;
  assign n49528 = n49527 ^ n38249;
  assign n55323 = n55322 ^ n49528;
  assign n44380 = n42146 ^ n33662;
  assign n44381 = n44380 ^ n38249;
  assign n44382 = n44381 ^ n31889;
  assign n55324 = n55323 ^ n44382;
  assign n19943 = n18070 ^ x465;
  assign n14801 = n12843 ^ x210;
  assign n14802 = n14801 ^ x402;
  assign n14803 = n14802 ^ x146;
  assign n19944 = n19943 ^ n14803;
  assign n19945 = n19944 ^ x401;
  assign n29297 = n27040 ^ n19945;
  assign n23874 = n21643 ^ n14803;
  assign n18692 = n16765 ^ x402;
  assign n18693 = n18692 ^ n515;
  assign n18694 = n18693 ^ x338;
  assign n23875 = n23874 ^ n18694;
  assign n13808 = x498 ^ x146;
  assign n13809 = n13808 ^ x338;
  assign n13810 = n13809 ^ x82;
  assign n23876 = n23875 ^ n13810;
  assign n29298 = n29297 ^ n23876;
  assign n18687 = n16760 ^ x401;
  assign n18688 = n18687 ^ n13810;
  assign n18689 = n18688 ^ x337;
  assign n29299 = n29298 ^ n18689;
  assign n636 = x465 ^ x113;
  assign n637 = n636 ^ x305;
  assign n638 = n637 ^ x49;
  assign n21852 = n19945 ^ n638;
  assign n16848 = n14803 ^ x305;
  assign n16849 = n16848 ^ x497;
  assign n16850 = n16849 ^ x241;
  assign n21853 = n21852 ^ n16850;
  assign n21854 = n21853 ^ x496;
  assign n31632 = n29299 ^ n21854;
  assign n25635 = n23876 ^ n16850;
  assign n20608 = n18694 ^ x497;
  assign n20609 = n20608 ^ n518;
  assign n20610 = n20609 ^ x433;
  assign n25636 = n25635 ^ n20610;
  assign n15585 = n13810 ^ x241;
  assign n15586 = n15585 ^ x433;
  assign n15587 = n15586 ^ x177;
  assign n25637 = n25636 ^ n15587;
  assign n31633 = n31632 ^ n25637;
  assign n20603 = n18689 ^ x496;
  assign n20604 = n20603 ^ n15587;
  assign n20605 = n20604 ^ x432;
  assign n31634 = n31633 ^ n20605;
  assign n685 = x496 ^ x144;
  assign n686 = n685 ^ x336;
  assign n687 = n686 ^ x80;
  assign n22361 = n20605 ^ n687;
  assign n17442 = n15587 ^ x336;
  assign n12448 = x433 ^ x81;
  assign n12449 = n12448 ^ x273;
  assign n12450 = n12449 ^ x17;
  assign n17443 = n17442 ^ n12450;
  assign n17444 = n17443 ^ x272;
  assign n22362 = n22361 ^ n17444;
  assign n531 = x432 ^ x80;
  assign n532 = n531 ^ x272;
  assign n533 = n532 ^ x16;
  assign n22363 = n22362 ^ n533;
  assign n34157 = n31634 ^ n22363;
  assign n18682 = n16850 ^ x400;
  assign n13771 = x497 ^ x145;
  assign n13772 = n13771 ^ x337;
  assign n13773 = n13772 ^ x81;
  assign n18683 = n18682 ^ n13773;
  assign n18684 = n18683 ^ x336;
  assign n27587 = n25637 ^ n18684;
  assign n22366 = n20610 ^ n13773;
  assign n520 = x434 ^ x82;
  assign n521 = n520 ^ x274;
  assign n522 = n521 ^ x18;
  assign n519 = n518 ^ x337;
  assign n523 = n522 ^ n519;
  assign n524 = n523 ^ x273;
  assign n22367 = n22366 ^ n524;
  assign n22368 = n22367 ^ n12450;
  assign n27588 = n27587 ^ n22368;
  assign n27589 = n27588 ^ n17444;
  assign n34158 = n34157 ^ n27589;
  assign n654 = n638 ^ x208;
  assign n655 = n654 ^ x400;
  assign n656 = n655 ^ x144;
  assign n23830 = n21854 ^ n656;
  assign n23831 = n23830 ^ n18684;
  assign n23832 = n23831 ^ n687;
  assign n34159 = n34158 ^ n23832;
  assign n672 = n656 ^ x303;
  assign n673 = n672 ^ x495;
  assign n674 = n673 ^ x239;
  assign n25630 = n23832 ^ n674;
  assign n20598 = n18684 ^ x495;
  assign n15580 = n13773 ^ x240;
  assign n15581 = n15580 ^ x432;
  assign n15582 = n15581 ^ x176;
  assign n20599 = n20598 ^ n15582;
  assign n20600 = n20599 ^ x431;
  assign n25631 = n25630 ^ n20600;
  assign n743 = n687 ^ x239;
  assign n744 = n743 ^ x431;
  assign n745 = n744 ^ x175;
  assign n25632 = n25631 ^ n745;
  assign n36451 = n34159 ^ n25632;
  assign n30122 = n27589 ^ n20600;
  assign n24155 = n22368 ^ n15582;
  assign n526 = n522 ^ x177;
  assign n527 = n526 ^ x369;
  assign n528 = n527 ^ x113;
  assign n525 = n524 ^ x432;
  assign n529 = n528 ^ n525;
  assign n530 = n529 ^ x368;
  assign n24156 = n24155 ^ n530;
  assign n14190 = n12450 ^ x176;
  assign n14191 = n14190 ^ x368;
  assign n14192 = n14191 ^ x112;
  assign n24157 = n24156 ^ n14192;
  assign n30123 = n30122 ^ n24157;
  assign n19312 = n17444 ^ x431;
  assign n19313 = n19312 ^ n14192;
  assign n19314 = n19313 ^ x367;
  assign n30124 = n30123 ^ n19314;
  assign n36452 = n36451 ^ n30124;
  assign n24288 = n22363 ^ n745;
  assign n24289 = n24288 ^ n19314;
  assign n540 = n533 ^ x175;
  assign n541 = n540 ^ x367;
  assign n542 = n541 ^ x111;
  assign n24290 = n24289 ^ n542;
  assign n36453 = n36452 ^ n24290;
  assign n696 = n674 ^ x398;
  assign n691 = x495 ^ x143;
  assign n692 = n691 ^ x335;
  assign n693 = n692 ^ x79;
  assign n697 = n696 ^ n693;
  assign n698 = n697 ^ x334;
  assign n27577 = n25632 ^ n698;
  assign n22475 = n20600 ^ n693;
  assign n17536 = n15582 ^ x335;
  assign n17537 = n17536 ^ n533;
  assign n17538 = n17537 ^ x271;
  assign n22476 = n22475 ^ n17538;
  assign n779 = x431 ^ x79;
  assign n780 = n779 ^ x271;
  assign n781 = n780 ^ x15;
  assign n22477 = n22476 ^ n781;
  assign n27578 = n27577 ^ n22477;
  assign n778 = n745 ^ x334;
  assign n782 = n781 ^ n778;
  assign n783 = n782 ^ x270;
  assign n27579 = n27578 ^ n783;
  assign n38745 = n36453 ^ n27579;
  assign n32402 = n30124 ^ n22477;
  assign n25806 = n24157 ^ n17538;
  assign n535 = n528 ^ x272;
  assign n536 = n535 ^ x464;
  assign n537 = n536 ^ x208;
  assign n534 = n533 ^ n530;
  assign n538 = n537 ^ n534;
  assign n539 = n538 ^ x463;
  assign n25807 = n25806 ^ n539;
  assign n15961 = n14192 ^ x271;
  assign n15962 = n15961 ^ x463;
  assign n15963 = n15962 ^ x207;
  assign n25808 = n25807 ^ n15963;
  assign n32403 = n32402 ^ n25808;
  assign n21134 = n19314 ^ n781;
  assign n21135 = n21134 ^ n15963;
  assign n21136 = n21135 ^ x462;
  assign n32404 = n32403 ^ n21136;
  assign n38746 = n38745 ^ n32404;
  assign n26503 = n24290 ^ n783;
  assign n26504 = n26503 ^ n21136;
  assign n555 = n542 ^ x270;
  assign n556 = n555 ^ x462;
  assign n557 = n556 ^ x206;
  assign n26505 = n26504 ^ n557;
  assign n38747 = n38746 ^ n26505;
  assign n729 = n693 ^ x238;
  assign n730 = n729 ^ x430;
  assign n731 = n730 ^ x174;
  assign n728 = n698 ^ x493;
  assign n732 = n731 ^ n728;
  assign n733 = n732 ^ x429;
  assign n30117 = n27579 ^ n733;
  assign n24561 = n22477 ^ n731;
  assign n19405 = n17538 ^ x430;
  assign n19406 = n19405 ^ n542;
  assign n19407 = n19406 ^ x366;
  assign n24562 = n24561 ^ n19407;
  assign n839 = n781 ^ x174;
  assign n840 = n839 ^ x366;
  assign n841 = n840 ^ x110;
  assign n24563 = n24562 ^ n841;
  assign n30118 = n30117 ^ n24563;
  assign n838 = n783 ^ x429;
  assign n842 = n841 ^ n838;
  assign n843 = n842 ^ x365;
  assign n30119 = n30118 ^ n843;
  assign n41003 = n38747 ^ n30119;
  assign n23060 = n21136 ^ n841;
  assign n18105 = n15963 ^ x366;
  assign n551 = x463 ^ x111;
  assign n552 = n551 ^ x303;
  assign n553 = n552 ^ x47;
  assign n18106 = n18105 ^ n553;
  assign n18107 = n18106 ^ x302;
  assign n23061 = n23060 ^ n18107;
  assign n709 = x462 ^ x110;
  assign n710 = n709 ^ x302;
  assign n711 = n710 ^ x46;
  assign n23062 = n23061 ^ n711;
  assign n34685 = n32404 ^ n23062;
  assign n28462 = n25808 ^ n19407;
  assign n545 = x464 ^ x112;
  assign n546 = n545 ^ x304;
  assign n547 = n546 ^ x48;
  assign n544 = n537 ^ x367;
  assign n548 = n547 ^ n544;
  assign n549 = n548 ^ x303;
  assign n543 = n542 ^ n539;
  assign n550 = n549 ^ n543;
  assign n554 = n553 ^ n550;
  assign n28463 = n28462 ^ n554;
  assign n28464 = n28463 ^ n18107;
  assign n34686 = n34685 ^ n28464;
  assign n34687 = n34686 ^ n24563;
  assign n41004 = n41003 ^ n34687;
  assign n28458 = n26505 ^ n843;
  assign n28459 = n28458 ^ n23062;
  assign n708 = n557 ^ x365;
  assign n712 = n711 ^ n708;
  assign n713 = n712 ^ x301;
  assign n28460 = n28459 ^ n713;
  assign n41005 = n41004 ^ n28460;
  assign n797 = x429 ^ x77;
  assign n798 = n797 ^ x269;
  assign n799 = n798 ^ x13;
  assign n765 = x493 ^ x141;
  assign n766 = n765 ^ x333;
  assign n767 = n766 ^ x77;
  assign n795 = n767 ^ n733;
  assign n790 = n731 ^ x333;
  assign n785 = x430 ^ x78;
  assign n786 = n785 ^ x270;
  assign n787 = n786 ^ x14;
  assign n791 = n790 ^ n787;
  assign n792 = n791 ^ x269;
  assign n796 = n795 ^ n792;
  assign n800 = n799 ^ n796;
  assign n32413 = n30119 ^ n800;
  assign n26496 = n24563 ^ n792;
  assign n21213 = n19407 ^ n787;
  assign n21214 = n21213 ^ n557;
  assign n21215 = n21214 ^ x461;
  assign n26497 = n26496 ^ n21215;
  assign n924 = n841 ^ x269;
  assign n925 = n924 ^ x461;
  assign n926 = n925 ^ x205;
  assign n26498 = n26497 ^ n926;
  assign n32414 = n32413 ^ n26498;
  assign n923 = n843 ^ n799;
  assign n927 = n926 ^ n923;
  assign n928 = n927 ^ x460;
  assign n32415 = n32414 ^ n928;
  assign n43108 = n41005 ^ n32415;
  assign n37125 = n34687 ^ n26498;
  assign n30686 = n28464 ^ n21215;
  assign n566 = n553 ^ x206;
  assign n567 = n566 ^ x398;
  assign n568 = n567 ^ x142;
  assign n560 = n547 ^ x207;
  assign n561 = n560 ^ x399;
  assign n562 = n561 ^ x143;
  assign n559 = n549 ^ x462;
  assign n563 = n562 ^ n559;
  assign n564 = n563 ^ x398;
  assign n558 = n557 ^ n554;
  assign n565 = n564 ^ n558;
  assign n569 = n568 ^ n565;
  assign n30687 = n30686 ^ n569;
  assign n19972 = n18107 ^ x461;
  assign n19973 = n19972 ^ n568;
  assign n19974 = n19973 ^ x397;
  assign n30688 = n30687 ^ n19974;
  assign n37126 = n37125 ^ n30688;
  assign n24956 = n23062 ^ n926;
  assign n24957 = n24956 ^ n19974;
  assign n754 = n711 ^ x205;
  assign n755 = n754 ^ x397;
  assign n756 = n755 ^ x141;
  assign n24958 = n24957 ^ n756;
  assign n37127 = n37126 ^ n24958;
  assign n43109 = n43108 ^ n37127;
  assign n30691 = n28460 ^ n928;
  assign n30692 = n30691 ^ n24958;
  assign n753 = n713 ^ x460;
  assign n757 = n756 ^ n753;
  assign n758 = n757 ^ x396;
  assign n30693 = n30692 ^ n758;
  assign n43110 = n43109 ^ n30693;
  assign n857 = n799 ^ x172;
  assign n858 = n857 ^ x364;
  assign n859 = n858 ^ x108;
  assign n825 = n767 ^ x236;
  assign n826 = n825 ^ x428;
  assign n827 = n826 ^ x172;
  assign n855 = n827 ^ n800;
  assign n850 = n792 ^ x428;
  assign n845 = n787 ^ x173;
  assign n846 = n845 ^ x365;
  assign n847 = n846 ^ x109;
  assign n851 = n850 ^ n847;
  assign n852 = n851 ^ x364;
  assign n856 = n855 ^ n852;
  assign n860 = n859 ^ n856;
  assign n34676 = n32415 ^ n860;
  assign n28453 = n26498 ^ n852;
  assign n23055 = n21215 ^ n847;
  assign n23056 = n23055 ^ n713;
  assign n984 = x461 ^ x109;
  assign n985 = n984 ^ x301;
  assign n986 = n985 ^ x45;
  assign n23057 = n23056 ^ n986;
  assign n28454 = n28453 ^ n23057;
  assign n983 = n926 ^ x364;
  assign n987 = n986 ^ n983;
  assign n988 = n987 ^ x300;
  assign n28455 = n28454 ^ n988;
  assign n34677 = n34676 ^ n28455;
  assign n982 = n928 ^ n859;
  assign n989 = n988 ^ n982;
  assign n810 = x460 ^ x108;
  assign n811 = n810 ^ x300;
  assign n812 = n811 ^ x44;
  assign n990 = n989 ^ n812;
  assign n34678 = n34677 ^ n990;
  assign n45059 = n43110 ^ n34678;
  assign n39140 = n37127 ^ n28455;
  assign n33273 = n30688 ^ n23057;
  assign n722 = n568 ^ x301;
  assign n723 = n722 ^ x493;
  assign n724 = n723 ^ x237;
  assign n715 = n562 ^ x302;
  assign n716 = n715 ^ x494;
  assign n717 = n716 ^ x238;
  assign n718 = n717 ^ n564;
  assign n719 = n718 ^ n711;
  assign n720 = n719 ^ x493;
  assign n714 = n713 ^ n569;
  assign n721 = n720 ^ n714;
  assign n725 = n724 ^ n721;
  assign n33274 = n33273 ^ n725;
  assign n21843 = n19974 ^ n986;
  assign n21844 = n21843 ^ n724;
  assign n21845 = n21844 ^ x492;
  assign n33275 = n33274 ^ n21845;
  assign n39141 = n39140 ^ n33275;
  assign n27066 = n24958 ^ n988;
  assign n27067 = n27066 ^ n21845;
  assign n814 = x492 ^ x300;
  assign n815 = n814 ^ n756;
  assign n816 = n815 ^ x236;
  assign n27068 = n27067 ^ n816;
  assign n39142 = n39141 ^ n27068;
  assign n45060 = n45059 ^ n39142;
  assign n33268 = n30693 ^ n990;
  assign n33269 = n33268 ^ n27068;
  assign n813 = n812 ^ n758;
  assign n817 = n816 ^ n813;
  assign n818 = n817 ^ x491;
  assign n33270 = n33269 ^ n818;
  assign n45061 = n45060 ^ n33270;
  assign n916 = n859 ^ x267;
  assign n917 = n916 ^ x459;
  assign n918 = n917 ^ x203;
  assign n910 = n847 ^ x268;
  assign n911 = n910 ^ x460;
  assign n912 = n911 ^ x204;
  assign n879 = x428 ^ x76;
  assign n880 = n879 ^ x268;
  assign n881 = n880 ^ x12;
  assign n909 = n881 ^ n852;
  assign n913 = n912 ^ n909;
  assign n914 = n913 ^ x459;
  assign n884 = n827 ^ x331;
  assign n885 = n884 ^ n881;
  assign n886 = n885 ^ x267;
  assign n908 = n886 ^ n860;
  assign n915 = n914 ^ n908;
  assign n919 = n918 ^ n915;
  assign n37116 = n34678 ^ n919;
  assign n30697 = n28455 ^ n914;
  assign n25092 = n23057 ^ n912;
  assign n25093 = n25092 ^ n758;
  assign n1081 = n986 ^ x204;
  assign n1082 = n1081 ^ x396;
  assign n1083 = n1082 ^ x140;
  assign n25094 = n25093 ^ n1083;
  assign n30698 = n30697 ^ n25094;
  assign n1080 = n988 ^ x459;
  assign n1084 = n1083 ^ n1080;
  assign n1085 = n1084 ^ x395;
  assign n30699 = n30698 ^ n1085;
  assign n37117 = n37116 ^ n30699;
  assign n1079 = n990 ^ n918;
  assign n1086 = n1085 ^ n1079;
  assign n899 = n812 ^ x203;
  assign n900 = n899 ^ x395;
  assign n901 = n900 ^ x139;
  assign n1087 = n1086 ^ n901;
  assign n37118 = n37117 ^ n1087;
  assign n46947 = n45061 ^ n37118;
  assign n41386 = n39142 ^ n30699;
  assign n35611 = n33275 ^ n25094;
  assign n770 = n724 ^ x396;
  assign n771 = n770 ^ n767;
  assign n772 = n771 ^ x332;
  assign n761 = n717 ^ x397;
  assign n703 = x494 ^ x142;
  assign n704 = n703 ^ x334;
  assign n705 = n704 ^ x78;
  assign n762 = n761 ^ n705;
  assign n763 = n762 ^ x333;
  assign n760 = n756 ^ n720;
  assign n764 = n763 ^ n760;
  assign n768 = n767 ^ n764;
  assign n759 = n758 ^ n725;
  assign n769 = n768 ^ n759;
  assign n773 = n772 ^ n769;
  assign n35612 = n35611 ^ n773;
  assign n23819 = n21845 ^ n1083;
  assign n23820 = n23819 ^ n772;
  assign n871 = x492 ^ x140;
  assign n872 = n871 ^ x332;
  assign n873 = n872 ^ x76;
  assign n23821 = n23820 ^ n873;
  assign n35613 = n35612 ^ n23821;
  assign n41387 = n41386 ^ n35613;
  assign n29369 = n27068 ^ n1085;
  assign n29370 = n29369 ^ n23821;
  assign n870 = n816 ^ x395;
  assign n874 = n873 ^ n870;
  assign n875 = n874 ^ x331;
  assign n29371 = n29370 ^ n875;
  assign n41388 = n41387 ^ n29371;
  assign n46948 = n46947 ^ n41388;
  assign n35607 = n33270 ^ n1087;
  assign n35608 = n35607 ^ n29371;
  assign n902 = n901 ^ n818;
  assign n903 = n902 ^ n875;
  assign n904 = n903 ^ n891;
  assign n35609 = n35608 ^ n904;
  assign n46949 = n46948 ^ n35609;
  assign n1007 = n918 ^ x362;
  assign n999 = x459 ^ x107;
  assign n1000 = n999 ^ x299;
  assign n1001 = n1000 ^ x43;
  assign n1008 = n1007 ^ n1001;
  assign n1009 = n1008 ^ x298;
  assign n966 = n886 ^ x426;
  assign n961 = n881 ^ x171;
  assign n962 = n961 ^ x363;
  assign n963 = n962 ^ x107;
  assign n967 = n966 ^ n963;
  assign n968 = n967 ^ x362;
  assign n1005 = n968 ^ n919;
  assign n997 = n963 ^ n914;
  assign n992 = n912 ^ x363;
  assign n993 = n992 ^ n812;
  assign n994 = n993 ^ x299;
  assign n998 = n997 ^ n994;
  assign n1002 = n1001 ^ n998;
  assign n1006 = n1005 ^ n1002;
  assign n1010 = n1009 ^ n1006;
  assign n39337 = n37118 ^ n1010;
  assign n33284 = n30699 ^ n1002;
  assign n27074 = n25094 ^ n994;
  assign n27075 = n27074 ^ n818;
  assign n1160 = n1083 ^ x299;
  assign n1161 = n1160 ^ x491;
  assign n1162 = n1161 ^ x235;
  assign n27076 = n27075 ^ n1162;
  assign n33285 = n33284 ^ n27076;
  assign n1163 = n1162 ^ n1001;
  assign n1164 = n1163 ^ n1085;
  assign n1165 = n1164 ^ x490;
  assign n33286 = n33285 ^ n1165;
  assign n39338 = n39337 ^ n33286;
  assign n1159 = n1087 ^ n1009;
  assign n1166 = n1165 ^ n1159;
  assign n942 = n901 ^ x298;
  assign n943 = n942 ^ x490;
  assign n944 = n943 ^ x234;
  assign n1167 = n1166 ^ n944;
  assign n39339 = n39338 ^ n1167;
  assign n49158 = n46949 ^ n39339;
  assign n43511 = n41388 ^ n33286;
  assign n37890 = n35613 ^ n27076;
  assign n830 = n772 ^ x491;
  assign n831 = n830 ^ n827;
  assign n832 = n831 ^ x427;
  assign n821 = n763 ^ x492;
  assign n735 = n705 ^ x237;
  assign n736 = n735 ^ x429;
  assign n737 = n736 ^ x173;
  assign n822 = n821 ^ n737;
  assign n823 = n822 ^ x428;
  assign n820 = n816 ^ n768;
  assign n824 = n823 ^ n820;
  assign n828 = n827 ^ n824;
  assign n819 = n818 ^ n773;
  assign n829 = n828 ^ n819;
  assign n833 = n832 ^ n829;
  assign n37891 = n37890 ^ n833;
  assign n25619 = n23821 ^ n1162;
  assign n25620 = n25619 ^ n832;
  assign n947 = n873 ^ x235;
  assign n948 = n947 ^ x427;
  assign n949 = n948 ^ x171;
  assign n25621 = n25620 ^ n949;
  assign n37892 = n37891 ^ n25621;
  assign n43512 = n43511 ^ n37892;
  assign n31608 = n29371 ^ n1165;
  assign n31609 = n31608 ^ n25621;
  assign n946 = n875 ^ x490;
  assign n950 = n949 ^ n946;
  assign n951 = n950 ^ x426;
  assign n31610 = n31609 ^ n951;
  assign n43513 = n43512 ^ n31610;
  assign n49159 = n49158 ^ n43513;
  assign n37886 = n35609 ^ n1167;
  assign n37887 = n37886 ^ n31610;
  assign n945 = n944 ^ n904;
  assign n952 = n951 ^ n945;
  assign n956 = n955 ^ n952;
  assign n37888 = n37887 ^ n956;
  assign n49160 = n49159 ^ n37888;
  assign n1094 = n1009 ^ x457;
  assign n1073 = n1001 ^ x202;
  assign n1074 = n1073 ^ x394;
  assign n1075 = n1074 ^ x138;
  assign n1095 = n1094 ^ n1075;
  assign n1096 = n1095 ^ x393;
  assign n1047 = n963 ^ x266;
  assign n1048 = n1047 ^ x458;
  assign n1049 = n1048 ^ x202;
  assign n1046 = n1037 ^ n968;
  assign n1050 = n1049 ^ n1046;
  assign n1051 = n1050 ^ x457;
  assign n1092 = n1051 ^ n1010;
  assign n1069 = n994 ^ x458;
  assign n1070 = n1069 ^ n901;
  assign n1071 = n1070 ^ x394;
  assign n1068 = n1049 ^ n1002;
  assign n1072 = n1071 ^ n1068;
  assign n1076 = n1075 ^ n1072;
  assign n1093 = n1092 ^ n1076;
  assign n1097 = n1096 ^ n1093;
  assign n41593 = n39339 ^ n1097;
  assign n35602 = n33286 ^ n1076;
  assign n29273 = n27076 ^ n1071;
  assign n29274 = n29273 ^ n904;
  assign n1260 = n1162 ^ x394;
  assign n1261 = n1260 ^ n891;
  assign n1262 = n1261 ^ x330;
  assign n29275 = n29274 ^ n1262;
  assign n35603 = n35602 ^ n29275;
  assign n1259 = n1165 ^ n1075;
  assign n1263 = n1262 ^ n1259;
  assign n1024 = x490 ^ x138;
  assign n1025 = n1024 ^ x330;
  assign n1026 = n1025 ^ x74;
  assign n1264 = n1263 ^ n1026;
  assign n35604 = n35603 ^ n1264;
  assign n41594 = n41593 ^ n35604;
  assign n1258 = n1167 ^ n1096;
  assign n1265 = n1264 ^ n1258;
  assign n1023 = n944 ^ x393;
  assign n1027 = n1026 ^ n1023;
  assign n1028 = n1027 ^ x329;
  assign n1266 = n1265 ^ n1028;
  assign n41595 = n41594 ^ n1266;
  assign n51195 = n49160 ^ n41595;
  assign n40248 = n37892 ^ n29275;
  assign n894 = x427 ^ x267;
  assign n895 = n894 ^ x75;
  assign n896 = n895 ^ x11;
  assign n892 = n891 ^ n832;
  assign n893 = n892 ^ n886;
  assign n897 = n896 ^ n893;
  assign n877 = n873 ^ n823;
  assign n805 = n737 ^ x332;
  assign n806 = n805 ^ n799;
  assign n807 = n806 ^ x268;
  assign n878 = n877 ^ n807;
  assign n882 = n881 ^ n878;
  assign n876 = n875 ^ n828;
  assign n883 = n882 ^ n876;
  assign n887 = n886 ^ n883;
  assign n888 = n887 ^ n833;
  assign n898 = n897 ^ n888;
  assign n905 = n904 ^ n898;
  assign n40249 = n40248 ^ n905;
  assign n27988 = n25621 ^ n1262;
  assign n27989 = n27988 ^ n897;
  assign n1031 = n949 ^ x330;
  assign n1032 = n1031 ^ n896;
  assign n1033 = n1032 ^ x266;
  assign n27990 = n27989 ^ n1033;
  assign n40250 = n40249 ^ n27990;
  assign n45858 = n40250 ^ n35604;
  assign n45859 = n45858 ^ n43513;
  assign n1030 = n1026 ^ n951;
  assign n1034 = n1033 ^ n1030;
  assign n1038 = n1037 ^ n1034;
  assign n34214 = n31610 ^ n1038;
  assign n34215 = n34214 ^ n27990;
  assign n34216 = n34215 ^ n1264;
  assign n45860 = n45859 ^ n34216;
  assign n51196 = n51195 ^ n45860;
  assign n40269 = n37888 ^ n1266;
  assign n40270 = n40269 ^ n34216;
  assign n1029 = n1028 ^ n956;
  assign n1039 = n1038 ^ n1029;
  assign n1043 = n1042 ^ n1039;
  assign n40271 = n40270 ^ n1043;
  assign n51197 = n51196 ^ n40271;
  assign n1142 = x457 ^ x297;
  assign n1143 = n1142 ^ x105;
  assign n1144 = n1143 ^ x41;
  assign n1184 = n1144 ^ n1096;
  assign n1176 = n1075 ^ x297;
  assign n1177 = n1176 ^ x489;
  assign n1178 = n1177 ^ x233;
  assign n1185 = n1184 ^ n1178;
  assign n1186 = n1185 ^ x488;
  assign n1140 = n1124 ^ n1051;
  assign n1135 = n1049 ^ x361;
  assign n1017 = x458 ^ x106;
  assign n1018 = n1017 ^ x298;
  assign n1019 = n1018 ^ x42;
  assign n1136 = n1135 ^ n1019;
  assign n1137 = n1136 ^ x297;
  assign n1141 = n1140 ^ n1137;
  assign n1145 = n1144 ^ n1141;
  assign n1182 = n1145 ^ n1097;
  assign n1174 = n1137 ^ n1076;
  assign n1169 = n1071 ^ n1019;
  assign n1170 = n1169 ^ n944;
  assign n1171 = n1170 ^ x489;
  assign n1175 = n1174 ^ n1171;
  assign n1179 = n1178 ^ n1175;
  assign n1183 = n1182 ^ n1179;
  assign n1187 = n1186 ^ n1183;
  assign n43723 = n41595 ^ n1187;
  assign n38025 = n35604 ^ n1179;
  assign n31603 = n29275 ^ n1171;
  assign n31604 = n31603 ^ n956;
  assign n1368 = n1262 ^ x489;
  assign n1369 = n1368 ^ n955;
  assign n1370 = n1369 ^ x425;
  assign n31605 = n31604 ^ n1370;
  assign n38026 = n38025 ^ n31605;
  assign n1367 = n1264 ^ n1178;
  assign n1371 = n1370 ^ n1367;
  assign n1111 = n1026 ^ x233;
  assign n1112 = n1111 ^ x425;
  assign n1113 = n1112 ^ x169;
  assign n1372 = n1371 ^ n1113;
  assign n38027 = n38026 ^ n1372;
  assign n43724 = n43723 ^ n38027;
  assign n1366 = n1266 ^ n1186;
  assign n1373 = n1372 ^ n1366;
  assign n1110 = n1028 ^ x488;
  assign n1114 = n1113 ^ n1110;
  assign n1115 = n1114 ^ x424;
  assign n1374 = n1373 ^ n1115;
  assign n43725 = n43724 ^ n1374;
  assign n53314 = n51197 ^ n43725;
  assign n47717 = n45860 ^ n38027;
  assign n42447 = n40250 ^ n31605;
  assign n973 = n896 ^ x170;
  assign n974 = n973 ^ x362;
  assign n975 = n974 ^ x106;
  assign n971 = n955 ^ n897;
  assign n972 = n971 ^ n968;
  assign n976 = n975 ^ n972;
  assign n959 = n949 ^ n882;
  assign n865 = n807 ^ x427;
  assign n866 = n865 ^ n859;
  assign n867 = n866 ^ x363;
  assign n960 = n959 ^ n867;
  assign n964 = n963 ^ n960;
  assign n958 = n951 ^ n887;
  assign n965 = n964 ^ n958;
  assign n969 = n968 ^ n965;
  assign n957 = n956 ^ n905;
  assign n970 = n969 ^ n957;
  assign n977 = n976 ^ n970;
  assign n42448 = n42447 ^ n977;
  assign n30106 = n27990 ^ n1370;
  assign n30107 = n30106 ^ n976;
  assign n1118 = n1033 ^ x425;
  assign n1119 = n1118 ^ n975;
  assign n1120 = n1119 ^ x361;
  assign n30108 = n30107 ^ n1120;
  assign n42449 = n42448 ^ n30108;
  assign n47718 = n47717 ^ n42449;
  assign n36427 = n34216 ^ n1372;
  assign n36428 = n36427 ^ n30108;
  assign n1117 = n1113 ^ n1038;
  assign n1121 = n1120 ^ n1117;
  assign n1125 = n1124 ^ n1121;
  assign n36429 = n36428 ^ n1125;
  assign n47719 = n47718 ^ n36429;
  assign n53315 = n53314 ^ n47719;
  assign n42430 = n40271 ^ n1374;
  assign n42431 = n42430 ^ n36429;
  assign n1116 = n1115 ^ n1043;
  assign n1126 = n1125 ^ n1116;
  assign n1130 = n1129 ^ n1126;
  assign n42432 = n42431 ^ n1130;
  assign n53316 = n53315 ^ n42432;
  assign n623 = n575 ^ x273;
  assign n624 = n623 ^ x465;
  assign n625 = n624 ^ x209;
  assign n617 = n610 ^ x274;
  assign n618 = n617 ^ x466;
  assign n619 = n618 ^ x210;
  assign n616 = n612 ^ n522;
  assign n620 = n619 ^ n616;
  assign n621 = n620 ^ x465;
  assign n615 = n614 ^ n524;
  assign n622 = n621 ^ n615;
  assign n626 = n625 ^ n622;
  assign n37146 = n34824 ^ n626;
  assign n30704 = n28482 ^ n621;
  assign n24968 = n23162 ^ n619;
  assign n24969 = n24968 ^ n19954;
  assign n24970 = n24969 ^ n14803;
  assign n30705 = n30704 ^ n24970;
  assign n30706 = n30705 ^ n19945;
  assign n37147 = n37146 ^ n30706;
  assign n24963 = n23074 ^ n625;
  assign n24964 = n24963 ^ n19945;
  assign n648 = n632 ^ x209;
  assign n649 = n648 ^ x401;
  assign n650 = n649 ^ x145;
  assign n24965 = n24964 ^ n650;
  assign n37148 = n37147 ^ n24965;
  assign n46977 = n45120 ^ n37148;
  assign n41412 = n39163 ^ n30706;
  assign n35639 = n33200 ^ n24970;
  assign n29302 = n26935 ^ n19954;
  assign n29303 = n29302 ^ n23842;
  assign n29304 = n29303 ^ n18694;
  assign n35640 = n35639 ^ n29304;
  assign n35641 = n35640 ^ n23876;
  assign n41413 = n41412 ^ n35641;
  assign n41414 = n41413 ^ n29299;
  assign n46978 = n46977 ^ n41414;
  assign n35634 = n33260 ^ n24965;
  assign n35635 = n35634 ^ n29299;
  assign n23835 = n21859 ^ n650;
  assign n23836 = n23835 ^ n18689;
  assign n23837 = n23836 ^ n13773;
  assign n35636 = n35635 ^ n23837;
  assign n46979 = n46978 ^ n35636;
  assign n641 = n625 ^ x368;
  assign n642 = n641 ^ n638;
  assign n643 = n642 ^ x304;
  assign n629 = n619 ^ x369;
  assign n633 = n632 ^ n629;
  assign n634 = n633 ^ x305;
  assign n628 = n621 ^ n528;
  assign n635 = n634 ^ n628;
  assign n639 = n638 ^ n635;
  assign n627 = n626 ^ n530;
  assign n640 = n639 ^ n627;
  assign n644 = n643 ^ n640;
  assign n39294 = n37148 ^ n644;
  assign n33253 = n30706 ^ n639;
  assign n26928 = n24970 ^ n634;
  assign n26929 = n26928 ^ n21859;
  assign n26930 = n26929 ^ n16850;
  assign n33254 = n33253 ^ n26930;
  assign n33255 = n33254 ^ n21854;
  assign n39295 = n39294 ^ n33255;
  assign n26923 = n24965 ^ n643;
  assign n26924 = n26923 ^ n21854;
  assign n666 = n650 ^ x304;
  assign n667 = n666 ^ x496;
  assign n668 = n667 ^ x240;
  assign n26925 = n26924 ^ n668;
  assign n39296 = n39295 ^ n26925;
  assign n49188 = n46979 ^ n39296;
  assign n43537 = n41414 ^ n33255;
  assign n37918 = n35641 ^ n26930;
  assign n37919 = n37918 ^ n25637;
  assign n31190 = n29304 ^ n21859;
  assign n31191 = n31190 ^ n25727;
  assign n31192 = n31191 ^ n20610;
  assign n37920 = n37919 ^ n31192;
  assign n43538 = n43537 ^ n37920;
  assign n43539 = n43538 ^ n31634;
  assign n49189 = n49188 ^ n43539;
  assign n37913 = n35636 ^ n26925;
  assign n37914 = n37913 ^ n31634;
  assign n25736 = n23837 ^ n668;
  assign n25737 = n25736 ^ n20605;
  assign n25738 = n25737 ^ n15582;
  assign n37915 = n37914 ^ n25738;
  assign n49190 = n49189 ^ n37915;
  assign n1797 = n1769 ^ n1736;
  assign n1792 = n1728 ^ x506;
  assign n1787 = n1723 ^ x251;
  assign n1788 = n1787 ^ x443;
  assign n1789 = n1788 ^ x187;
  assign n1793 = n1792 ^ n1789;
  assign n1794 = n1793 ^ x442;
  assign n1798 = n1797 ^ n1794;
  assign n1802 = n1801 ^ n1798;
  assign n1875 = n1838 ^ n1802;
  assign n1862 = n1789 ^ x346;
  assign n1863 = n1862 ^ n1691;
  assign n1864 = n1863 ^ x282;
  assign n1867 = n1864 ^ n1794;
  assign n1868 = n1867 ^ n1833;
  assign n1872 = n1871 ^ n1868;
  assign n1876 = n1875 ^ n1872;
  assign n1880 = n1879 ^ n1876;
  assign n1959 = n1922 ^ n1880;
  assign n1951 = n1917 ^ n1872;
  assign n1946 = n1864 ^ x441;
  assign n1947 = n1946 ^ n1757;
  assign n1948 = n1947 ^ x377;
  assign n1952 = n1951 ^ n1948;
  assign n1956 = n1955 ^ n1952;
  assign n1960 = n1959 ^ n1956;
  assign n1964 = n1963 ^ n1960;
  assign n2049 = n2012 ^ n1964;
  assign n2041 = n2004 ^ n1956;
  assign n2036 = n1948 ^ n1889;
  assign n2037 = n2036 ^ n1823;
  assign n2038 = n2037 ^ x472;
  assign n2042 = n2041 ^ n2038;
  assign n2046 = n2045 ^ n2042;
  assign n2050 = n2049 ^ n2046;
  assign n2054 = n2053 ^ n2050;
  assign n2142 = n2102 ^ n2054;
  assign n2134 = n2094 ^ n2046;
  assign n2126 = n2038 ^ n1973;
  assign n2127 = n2126 ^ n1901;
  assign n2131 = n2130 ^ n2127;
  assign n2135 = n2134 ^ n2131;
  assign n2139 = n2138 ^ n2135;
  assign n2143 = n2142 ^ n2139;
  assign n2147 = n2146 ^ n2143;
  assign n2247 = n2207 ^ n2147;
  assign n2251 = n2250 ^ n2247;
  assign n2239 = n2199 ^ n2139;
  assign n2231 = n2131 ^ n2063;
  assign n2232 = n2231 ^ n1988;
  assign n2236 = n2235 ^ n2232;
  assign n2240 = n2239 ^ n2236;
  assign n2244 = n2243 ^ n2240;
  assign n2252 = n2251 ^ n2244;
  assign n39171 = n28497 ^ n2252;
  assign n33213 = n23089 ^ n2244;
  assign n26948 = n2236 ^ n2156;
  assign n26949 = n26948 ^ n2078;
  assign n26950 = n26949 ^ n16830;
  assign n33214 = n33213 ^ n26950;
  assign n33215 = n33214 ^ n21548;
  assign n39172 = n39171 ^ n33215;
  assign n39173 = n39172 ^ n26945;
  assign n41528 = n39173 ^ n30579;
  assign n35654 = n33215 ^ n24985;
  assign n29317 = n26950 ^ n2261;
  assign n29318 = n29317 ^ n2183;
  assign n29319 = n29318 ^ n18706;
  assign n35655 = n35654 ^ n29319;
  assign n35656 = n35655 ^ n23847;
  assign n41529 = n41528 ^ n35656;
  assign n41530 = n41529 ^ n29314;
  assign n43542 = n41530 ^ n33205;
  assign n37987 = n35656 ^ n26940;
  assign n31205 = n29319 ^ n21543;
  assign n31206 = n31205 ^ n25701;
  assign n31207 = n31206 ^ n20617;
  assign n37988 = n37987 ^ n31207;
  assign n37989 = n37988 ^ n25709;
  assign n43543 = n43542 ^ n37989;
  assign n43544 = n43543 ^ n31202;
  assign n35644 = n33205 ^ n24975;
  assign n29307 = n26940 ^ n19747;
  assign n23863 = n21543 ^ n14726;
  assign n23864 = n23863 ^ n590;
  assign n23865 = n23864 ^ n13799;
  assign n29308 = n29307 ^ n23865;
  assign n29309 = n29308 ^ n18699;
  assign n35645 = n35644 ^ n29309;
  assign n35646 = n35645 ^ n23842;
  assign n45499 = n43544 ^ n35646;
  assign n39861 = n37989 ^ n29309;
  assign n33642 = n31207 ^ n23865;
  assign n33643 = n33642 ^ n27604;
  assign n33644 = n33643 ^ n22450;
  assign n39862 = n39861 ^ n33644;
  assign n39863 = n39862 ^ n27665;
  assign n45500 = n45499 ^ n39863;
  assign n45501 = n45500 ^ n33639;
  assign n37923 = n35646 ^ n27040;
  assign n31195 = n29309 ^ n21643;
  assign n25717 = n23865 ^ n16765;
  assign n25718 = n25717 ^ n596;
  assign n25719 = n25718 ^ n15592;
  assign n31196 = n31195 ^ n25719;
  assign n31197 = n31196 ^ n20632;
  assign n37924 = n37923 ^ n31197;
  assign n37925 = n37924 ^ n25727;
  assign n47865 = n45501 ^ n37925;
  assign n42238 = n39863 ^ n31197;
  assign n36466 = n33644 ^ n25719;
  assign n36467 = n36466 ^ n29735;
  assign n36468 = n36467 ^ n24164;
  assign n42239 = n42238 ^ n36468;
  assign n42240 = n42239 ^ n29636;
  assign n47866 = n47865 ^ n42240;
  assign n47867 = n47866 ^ n36489;
  assign n1681 = n1635 ^ x315;
  assign n1682 = n1681 ^ x507;
  assign n1683 = n1682 ^ x251;
  assign n1741 = n1683 ^ x410;
  assign n1742 = n1741 ^ n1735;
  assign n1743 = n1742 ^ x346;
  assign n1807 = n1743 ^ x505;
  assign n1808 = n1807 ^ n1801;
  assign n1809 = n1808 ^ x441;
  assign n1586 = n1484 ^ n1459;
  assign n1587 = n1586 ^ n1583;
  assign n1591 = n1590 ^ n1587;
  assign n1631 = n1628 ^ n1591;
  assign n1632 = n1631 ^ n1618;
  assign n1636 = n1635 ^ n1632;
  assign n1679 = n1657 ^ n1636;
  assign n1680 = n1679 ^ n1676;
  assign n1684 = n1683 ^ n1680;
  assign n1739 = n1708 ^ n1684;
  assign n1740 = n1739 ^ n1736;
  assign n1744 = n1743 ^ n1740;
  assign n1805 = n1774 ^ n1744;
  assign n1806 = n1805 ^ n1802;
  assign n1810 = n1809 ^ n1806;
  assign n37942 = n27012 ^ n1810;
  assign n28508 = n26149 ^ n19351;
  assign n28509 = n28508 ^ n1591;
  assign n28510 = n28509 ^ n1648;
  assign n30606 = n28510 ^ n20829;
  assign n30607 = n30606 ^ n1636;
  assign n30608 = n30607 ^ n1699;
  assign n32666 = n30608 ^ n23100;
  assign n32667 = n32666 ^ n1684;
  assign n1763 = n1751 ^ n1699;
  assign n1764 = n1763 ^ n1683;
  assign n1765 = n1764 ^ x506;
  assign n32668 = n32667 ^ n1765;
  assign n35675 = n32668 ^ n24994;
  assign n35676 = n35675 ^ n1744;
  assign n1829 = n1817 ^ n1765;
  assign n1830 = n1829 ^ n1743;
  assign n1834 = n1833 ^ n1830;
  assign n35677 = n35676 ^ n1834;
  assign n37943 = n37942 ^ n35677;
  assign n1913 = n1906 ^ n1834;
  assign n1914 = n1913 ^ n1809;
  assign n1918 = n1917 ^ n1914;
  assign n37944 = n37943 ^ n1918;
  assign n39877 = n37944 ^ n28866;
  assign n1885 = n1843 ^ n1809;
  assign n1886 = n1885 ^ n1879;
  assign n1890 = n1889 ^ n1886;
  assign n1883 = n1846 ^ n1810;
  assign n1884 = n1883 ^ n1880;
  assign n1891 = n1890 ^ n1884;
  assign n39878 = n39877 ^ n1891;
  assign n2000 = n1993 ^ n1918;
  assign n2001 = n2000 ^ n1890;
  assign n2005 = n2004 ^ n2001;
  assign n39879 = n39878 ^ n2005;
  assign n42131 = n39879 ^ n31219;
  assign n1969 = n1927 ^ n1890;
  assign n1970 = n1969 ^ n1963;
  assign n1974 = n1973 ^ n1970;
  assign n1967 = n1930 ^ n1891;
  assign n1968 = n1967 ^ n1964;
  assign n1975 = n1974 ^ n1968;
  assign n42132 = n42131 ^ n1975;
  assign n2090 = n2083 ^ n2005;
  assign n2091 = n2090 ^ n1974;
  assign n2095 = n2094 ^ n2091;
  assign n42133 = n42132 ^ n2095;
  assign n44311 = n42133 ^ n33656;
  assign n2059 = n2017 ^ n1974;
  assign n2060 = n2059 ^ n2053;
  assign n2064 = n2063 ^ n2060;
  assign n2057 = n2020 ^ n1975;
  assign n2058 = n2057 ^ n2054;
  assign n2065 = n2064 ^ n2058;
  assign n44312 = n44311 ^ n2065;
  assign n2195 = n2188 ^ n2095;
  assign n2196 = n2195 ^ n2064;
  assign n2200 = n2199 ^ n2196;
  assign n44313 = n44312 ^ n2200;
  assign n46128 = n44313 ^ n35953;
  assign n2152 = n2107 ^ n2064;
  assign n2153 = n2152 ^ n2146;
  assign n2157 = n2156 ^ n2153;
  assign n2150 = n2110 ^ n2065;
  assign n2151 = n2150 ^ n2147;
  assign n2158 = n2157 ^ n2151;
  assign n46129 = n46128 ^ n2158;
  assign n34720 = n24174 ^ n2200;
  assign n34721 = n34720 ^ n2157;
  assign n34722 = n34721 ^ n23089;
  assign n46130 = n46129 ^ n34722;
  assign n1270 = x489 ^ x137;
  assign n1271 = n1270 ^ x329;
  assign n1272 = n1271 ^ x73;
  assign n1103 = n1019 ^ x201;
  assign n1104 = n1103 ^ x393;
  assign n1105 = n1104 ^ x137;
  assign n1268 = n1171 ^ n1105;
  assign n1269 = n1268 ^ n1028;
  assign n1273 = n1272 ^ n1269;
  assign n34219 = n31605 ^ n1273;
  assign n34220 = n34219 ^ n1043;
  assign n22352 = n1370 ^ n1272;
  assign n22353 = n22352 ^ n1042;
  assign n1205 = x425 ^ x73;
  assign n1206 = n1205 ^ x265;
  assign n1207 = n1206 ^ x9;
  assign n22354 = n22353 ^ n1207;
  assign n34221 = n34220 ^ n22354;
  assign n1378 = n1272 ^ x232;
  assign n1379 = n1378 ^ x424;
  assign n1380 = n1379 ^ x168;
  assign n1194 = n1105 ^ x296;
  assign n1195 = n1194 ^ x488;
  assign n1196 = n1195 ^ x232;
  assign n1376 = n1273 ^ n1196;
  assign n1377 = n1376 ^ n1115;
  assign n1381 = n1380 ^ n1377;
  assign n36422 = n34221 ^ n1381;
  assign n36423 = n36422 ^ n1130;
  assign n24548 = n22354 ^ n1380;
  assign n24549 = n24548 ^ n1129;
  assign n1307 = n1207 ^ x168;
  assign n1308 = n1307 ^ x360;
  assign n1309 = n1308 ^ x104;
  assign n24550 = n24549 ^ n1309;
  assign n36424 = n36423 ^ n24550;
  assign n2655 = ~x30 & ~x31;
  assign n2656 = x29 & ~n2655;
  assign n2657 = x28 & n2656;
  assign n2658 = ~x27 & ~n2657;
  assign n2659 = ~x26 & n2658;
  assign n2660 = x25 & ~n2659;
  assign n2661 = ~x24 & ~n2660;
  assign n2662 = x23 & ~n2661;
  assign n2663 = x22 & n2662;
  assign n2664 = x21 & n2663;
  assign n2665 = ~x20 & ~n2664;
  assign n2666 = ~x19 & n2665;
  assign n2667 = x18 & ~n2666;
  assign n2668 = x17 & n2667;
  assign n2669 = ~x16 & ~n2668;
  assign n2670 = x15 & ~n2669;
  assign n2671 = x14 & n2670;
  assign n2930 = n2671 ^ x13;
  assign n2733 = n2656 ^ x28;
  assign n2734 = n2655 ^ x29;
  assign n2735 = x31 ^ x30;
  assign n2672 = ~x13 & ~n2671;
  assign n2673 = x12 & ~n2672;
  assign n2674 = ~x11 & ~n2673;
  assign n2675 = ~x10 & n2674;
  assign n2676 = x9 & ~n2675;
  assign n2677 = ~x8 & ~n2676;
  assign n2678 = ~x7 & n2677;
  assign n2679 = ~x6 & n2678;
  assign n2680 = ~x5 & n2679;
  assign n2681 = ~x4 & n2680;
  assign n2683 = ~x3 & n2681;
  assign n2689 = x2 & ~n2683;
  assign n2710 = x1 & n2689;
  assign n2711 = n2710 ^ x0;
  assign n2682 = n2681 ^ x3;
  assign n2684 = n2683 ^ x2;
  assign n2688 = ~n2682 & n2684;
  assign n2690 = n2689 ^ x1;
  assign n2736 = n2688 & ~n2690;
  assign n2737 = n2711 & n2736;
  assign n2738 = x31 & n2737;
  assign n2739 = n2735 & n2738;
  assign n2740 = n2734 & n2739;
  assign n2741 = n2733 & ~n2740;
  assign n2732 = n2657 ^ x27;
  assign n2776 = n2741 ^ n2732;
  assign n2766 = n2740 ^ n2733;
  assign n2767 = n2739 ^ n2734;
  assign n2768 = n2737 ^ x31;
  assign n2685 = n2682 & n2684;
  assign n2691 = n2690 ^ n2688;
  assign n2769 = ~n2685 & n2691;
  assign n2770 = n2711 & ~n2769;
  assign n2771 = n2768 & n2770;
  assign n2772 = n2738 ^ n2735;
  assign n2773 = n2771 & n2772;
  assign n2774 = ~n2767 & ~n2773;
  assign n2775 = ~n2766 & n2774;
  assign n2800 = n2776 ^ n2775;
  assign n2801 = n2773 ^ n2767;
  assign n2802 = n2772 ^ n2771;
  assign n2803 = n2770 ^ n2768;
  assign n2709 = ~n2684 & n2690;
  assign n2712 = n2711 ^ n2709;
  assign n2686 = n2680 ^ x4;
  assign n2713 = n2691 ^ n2685;
  assign n2714 = ~n2691 & n2713;
  assign n2715 = n2686 & n2714;
  assign n2716 = n2715 ^ n2713;
  assign n2804 = ~n2712 & n2716;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = ~n2802 & n2805;
  assign n2807 = ~n2801 & ~n2806;
  assign n2808 = n2774 ^ n2766;
  assign n2809 = n2807 & n2808;
  assign n2810 = n2800 & ~n2809;
  assign n2777 = n2775 & n2776;
  assign n2742 = n2732 & ~n2741;
  assign n2725 = n2658 ^ x26;
  assign n2765 = n2742 ^ n2725;
  assign n2811 = n2777 ^ n2765;
  assign n2812 = n2810 & ~n2811;
  assign n2744 = n2659 ^ x25;
  assign n2743 = ~n2725 & n2742;
  assign n2779 = n2744 ^ n2743;
  assign n2778 = ~n2765 & ~n2777;
  assign n2813 = n2779 ^ n2778;
  assign n2814 = ~n2812 & ~n2813;
  assign n2746 = n2660 ^ x24;
  assign n2745 = n2743 & n2744;
  assign n2781 = n2746 ^ n2745;
  assign n2780 = ~n2778 & ~n2779;
  assign n2815 = n2781 ^ n2780;
  assign n2816 = n2814 & ~n2815;
  assign n2748 = n2661 ^ x23;
  assign n2747 = n2745 & n2746;
  assign n2783 = n2748 ^ n2747;
  assign n2782 = ~n2780 & n2781;
  assign n2817 = n2783 ^ n2782;
  assign n2818 = n2816 & ~n2817;
  assign n2749 = n2747 & n2748;
  assign n2720 = n2662 ^ x22;
  assign n2785 = n2749 ^ n2720;
  assign n2784 = ~n2782 & ~n2783;
  assign n2819 = n2785 ^ n2784;
  assign n2820 = n2818 & n2819;
  assign n2786 = ~n2784 & ~n2785;
  assign n2750 = ~n2720 & n2749;
  assign n2731 = n2663 ^ x21;
  assign n2764 = n2750 ^ n2731;
  assign n2799 = n2786 ^ n2764;
  assign n2885 = n2820 ^ n2799;
  assign n2880 = n2819 ^ n2818;
  assign n2875 = n2817 ^ n2816;
  assign n2870 = n2815 ^ n2814;
  assign n2865 = n2813 ^ n2812;
  assign n2860 = n2811 ^ n2810;
  assign n2832 = n2809 ^ n2800;
  assign n2833 = n2832 ^ x54;
  assign n2852 = n2808 ^ n2807;
  assign n2847 = n2806 ^ n2801;
  assign n2834 = n2805 ^ n2802;
  assign n2835 = n2834 ^ x57;
  assign n2836 = n2804 ^ n2803;
  assign n2837 = n2836 ^ x58;
  assign n2717 = n2716 ^ n2712;
  assign n2687 = n2685 & ~n2686;
  assign n2692 = n2691 ^ n2687;
  assign n2693 = n2692 ^ x60;
  assign n2694 = n2682 & n2686;
  assign n2695 = n2694 ^ n2684;
  assign n2696 = n2695 ^ x61;
  assign n2697 = x63 & ~n2686;
  assign n2698 = n2697 ^ x62;
  assign n2699 = n2686 ^ n2682;
  assign n2700 = n2699 ^ n2697;
  assign n2701 = n2698 & ~n2700;
  assign n2702 = n2701 ^ x62;
  assign n2703 = n2702 ^ n2695;
  assign n2704 = n2696 & ~n2703;
  assign n2705 = n2704 ^ x61;
  assign n2706 = n2705 ^ n2692;
  assign n2707 = n2693 & ~n2706;
  assign n2708 = n2707 ^ x60;
  assign n2718 = n2717 ^ n2708;
  assign n2838 = n2717 ^ x59;
  assign n2839 = ~n2718 & n2838;
  assign n2840 = n2839 ^ x59;
  assign n2841 = n2840 ^ n2836;
  assign n2842 = n2837 & ~n2841;
  assign n2843 = n2842 ^ x58;
  assign n2844 = n2843 ^ n2834;
  assign n2845 = ~n2835 & n2844;
  assign n2846 = n2845 ^ x57;
  assign n2848 = n2847 ^ n2846;
  assign n2849 = n2847 ^ x56;
  assign n2850 = n2848 & ~n2849;
  assign n2851 = n2850 ^ x56;
  assign n2853 = n2852 ^ n2851;
  assign n2854 = n2852 ^ x55;
  assign n2855 = n2853 & ~n2854;
  assign n2856 = n2855 ^ x55;
  assign n2857 = n2856 ^ n2832;
  assign n2858 = ~n2833 & n2857;
  assign n2859 = n2858 ^ x54;
  assign n2861 = n2860 ^ n2859;
  assign n2862 = n2860 ^ x53;
  assign n2863 = n2861 & ~n2862;
  assign n2864 = n2863 ^ x53;
  assign n2866 = n2865 ^ n2864;
  assign n2867 = n2865 ^ x52;
  assign n2868 = n2866 & ~n2867;
  assign n2869 = n2868 ^ x52;
  assign n2871 = n2870 ^ n2869;
  assign n2872 = n2870 ^ x51;
  assign n2873 = ~n2871 & n2872;
  assign n2874 = n2873 ^ x51;
  assign n2876 = n2875 ^ n2874;
  assign n2877 = n2875 ^ x50;
  assign n2878 = ~n2876 & n2877;
  assign n2879 = n2878 ^ x50;
  assign n2881 = n2880 ^ n2879;
  assign n2882 = n2880 ^ x49;
  assign n2883 = n2881 & ~n2882;
  assign n2884 = n2883 ^ x49;
  assign n2886 = n2885 ^ n2884;
  assign n2887 = n2885 ^ x48;
  assign n2888 = ~n2886 & n2887;
  assign n2889 = n2888 ^ x48;
  assign n2821 = ~n2799 & ~n2820;
  assign n2787 = n2764 & ~n2786;
  assign n2751 = ~n2731 & n2750;
  assign n2730 = n2664 ^ x20;
  assign n2763 = n2751 ^ n2730;
  assign n2798 = n2787 ^ n2763;
  assign n2830 = n2821 ^ n2798;
  assign n2831 = n2830 ^ x47;
  assign n3150 = n2889 ^ n2831;
  assign n3507 = n2930 & ~n3150;
  assign n3033 = n2699 ^ n2698;
  assign n2724 = n2686 ^ x63;
  assign n2726 = n2725 ^ n2724;
  assign n3007 = n2678 ^ x6;
  assign n2939 = n2672 ^ x12;
  assign n2727 = n2668 ^ x16;
  assign n2728 = n2666 ^ x18;
  assign n2729 = n2665 ^ x19;
  assign n2752 = n2730 & n2751;
  assign n2753 = ~n2729 & n2752;
  assign n2754 = ~n2728 & ~n2753;
  assign n2755 = n2667 ^ x17;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = n2727 & n2756;
  assign n2758 = n2669 ^ x15;
  assign n2918 = n2757 & n2758;
  assign n2919 = n2670 ^ x14;
  assign n2929 = n2918 & ~n2919;
  assign n2940 = n2929 & n2930;
  assign n2950 = n2939 & n2940;
  assign n2951 = n2673 ^ x11;
  assign n2962 = n2950 & n2951;
  assign n2963 = n2674 ^ x10;
  assign n2972 = ~n2962 & n2963;
  assign n2973 = n2675 ^ x9;
  assign n2983 = ~n2972 & n2973;
  assign n2984 = n2676 ^ x8;
  assign n2994 = n2983 & n2984;
  assign n2995 = n2677 ^ x7;
  assign n3006 = n2994 & ~n2995;
  assign n3008 = n3007 ^ n3006;
  assign n2996 = n2995 ^ n2994;
  assign n2985 = n2984 ^ n2983;
  assign n2952 = n2951 ^ n2950;
  assign n2941 = n2940 ^ n2939;
  assign n2759 = n2758 ^ n2757;
  assign n2760 = n2756 ^ n2727;
  assign n2761 = n2753 ^ n2728;
  assign n2762 = n2752 ^ n2729;
  assign n2788 = ~n2763 & n2787;
  assign n2789 = ~n2762 & ~n2788;
  assign n2790 = n2761 & ~n2789;
  assign n2791 = n2755 ^ n2754;
  assign n2792 = n2790 & ~n2791;
  assign n2793 = n2760 & ~n2792;
  assign n2917 = n2759 & n2793;
  assign n2920 = n2919 ^ n2918;
  assign n2928 = ~n2917 & n2920;
  assign n2931 = n2930 ^ n2929;
  assign n2942 = n2928 & ~n2931;
  assign n2953 = ~n2941 & n2942;
  assign n2961 = ~n2952 & n2953;
  assign n2964 = n2963 ^ n2962;
  assign n2971 = n2961 & ~n2964;
  assign n2974 = n2973 ^ n2972;
  assign n2986 = n2971 & n2974;
  assign n2997 = n2985 & ~n2986;
  assign n3005 = n2996 & ~n2997;
  assign n3009 = n3008 ^ n3005;
  assign n2975 = n2974 ^ n2971;
  assign n2794 = n2793 ^ n2759;
  assign n2795 = n2791 ^ n2790;
  assign n2796 = n2789 ^ n2761;
  assign n2797 = n2788 ^ n2762;
  assign n2822 = ~n2798 & n2821;
  assign n2823 = n2797 & ~n2822;
  assign n2824 = ~n2796 & ~n2823;
  assign n2825 = ~n2795 & n2824;
  assign n2826 = n2792 ^ n2760;
  assign n2827 = n2825 & n2826;
  assign n2916 = ~n2794 & n2827;
  assign n2921 = n2920 ^ n2917;
  assign n2927 = n2916 & ~n2921;
  assign n2932 = n2931 ^ n2928;
  assign n2938 = ~n2927 & n2932;
  assign n2943 = n2942 ^ n2941;
  assign n2949 = ~n2938 & ~n2943;
  assign n2954 = n2953 ^ n2952;
  assign n2960 = ~n2949 & n2954;
  assign n2965 = n2964 ^ n2961;
  assign n2976 = ~n2960 & ~n2965;
  assign n2982 = ~n2975 & ~n2976;
  assign n2987 = n2986 ^ n2985;
  assign n2993 = n2982 & ~n2987;
  assign n2998 = n2997 ^ n2996;
  assign n3004 = ~n2993 & ~n2998;
  assign n3010 = n3009 ^ n3004;
  assign n2999 = n2998 ^ n2993;
  assign n2988 = n2987 ^ n2982;
  assign n2977 = n2976 ^ n2975;
  assign n2966 = n2965 ^ n2960;
  assign n2955 = n2954 ^ n2949;
  assign n2944 = n2943 ^ n2938;
  assign n2933 = n2932 ^ n2927;
  assign n2922 = n2921 ^ n2916;
  assign n2828 = n2827 ^ n2794;
  assign n2829 = n2828 ^ x42;
  assign n2908 = n2826 ^ n2825;
  assign n2903 = n2824 ^ n2795;
  assign n2898 = n2823 ^ n2796;
  assign n2893 = n2822 ^ n2797;
  assign n2890 = n2889 ^ n2830;
  assign n2891 = ~n2831 & n2890;
  assign n2892 = n2891 ^ x47;
  assign n2894 = n2893 ^ n2892;
  assign n2895 = n2893 ^ x46;
  assign n2896 = ~n2894 & n2895;
  assign n2897 = n2896 ^ x46;
  assign n2899 = n2898 ^ n2897;
  assign n2900 = n2898 ^ x45;
  assign n2901 = ~n2899 & n2900;
  assign n2902 = n2901 ^ x45;
  assign n2904 = n2903 ^ n2902;
  assign n2905 = n2903 ^ x44;
  assign n2906 = n2904 & ~n2905;
  assign n2907 = n2906 ^ x44;
  assign n2909 = n2908 ^ n2907;
  assign n2910 = n2908 ^ x43;
  assign n2911 = ~n2909 & n2910;
  assign n2912 = n2911 ^ x43;
  assign n2913 = n2912 ^ n2828;
  assign n2914 = ~n2829 & n2913;
  assign n2915 = n2914 ^ x42;
  assign n2923 = n2922 ^ n2915;
  assign n2924 = n2922 ^ x41;
  assign n2925 = n2923 & ~n2924;
  assign n2926 = n2925 ^ x41;
  assign n2934 = n2933 ^ n2926;
  assign n2935 = n2933 ^ x40;
  assign n2936 = ~n2934 & n2935;
  assign n2937 = n2936 ^ x40;
  assign n2945 = n2944 ^ n2937;
  assign n2946 = n2944 ^ x39;
  assign n2947 = ~n2945 & n2946;
  assign n2948 = n2947 ^ x39;
  assign n2956 = n2955 ^ n2948;
  assign n2957 = n2955 ^ x38;
  assign n2958 = ~n2956 & n2957;
  assign n2959 = n2958 ^ x38;
  assign n2967 = n2966 ^ n2959;
  assign n2968 = n2966 ^ x37;
  assign n2969 = ~n2967 & n2968;
  assign n2970 = n2969 ^ x37;
  assign n2978 = n2977 ^ n2970;
  assign n2979 = n2977 ^ x36;
  assign n2980 = n2978 & ~n2979;
  assign n2981 = n2980 ^ x36;
  assign n2989 = n2988 ^ n2981;
  assign n2990 = n2988 ^ x35;
  assign n2991 = ~n2989 & n2990;
  assign n2992 = n2991 ^ x35;
  assign n3000 = n2999 ^ n2992;
  assign n3001 = n2999 ^ x34;
  assign n3002 = ~n3000 & n3001;
  assign n3003 = n3002 ^ x34;
  assign n3011 = n3010 ^ n3003;
  assign n3012 = n3011 ^ x33;
  assign n3013 = n2989 ^ x35;
  assign n3014 = n2735 & n3013;
  assign n3015 = n3000 ^ x34;
  assign n3016 = n3014 & n3015;
  assign n3017 = ~n3012 & n3016;
  assign n3025 = n2679 ^ x5;
  assign n3021 = ~n3004 & ~n3009;
  assign n3022 = n3021 ^ n3006;
  assign n3023 = ~n3008 & ~n3022;
  assign n3024 = n3023 ^ n3007;
  assign n3026 = n3025 ^ n3024;
  assign n3018 = n3010 ^ x33;
  assign n3019 = n3011 & ~n3018;
  assign n3020 = n3019 ^ x33;
  assign n3027 = n3026 ^ n3020;
  assign n3028 = n3027 ^ x32;
  assign n3029 = n3017 & n3028;
  assign n3030 = n3029 ^ n2724;
  assign n3031 = n2726 & n3030;
  assign n3032 = n3031 ^ n2725;
  assign n3050 = n3033 ^ n3032;
  assign n3051 = n3029 ^ n2726;
  assign n3052 = n3015 ^ n3014;
  assign n3053 = n3013 ^ n2735;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = n3016 ^ n3012;
  assign n3056 = n3054 & n3055;
  assign n3057 = n3028 ^ n3017;
  assign n3058 = n3056 & ~n3057;
  assign n3059 = ~n3051 & n3058;
  assign n3060 = ~n3050 & n3059;
  assign n3034 = n3032 & ~n3033;
  assign n2722 = n2702 ^ x61;
  assign n2723 = n2722 ^ n2695;
  assign n3061 = n3034 ^ n2723;
  assign n3062 = n3060 & ~n3061;
  assign n3036 = n2705 ^ n2693;
  assign n3035 = ~n2723 & n3034;
  assign n3063 = n3036 ^ n3035;
  assign n3064 = ~n3062 & ~n3063;
  assign n3037 = ~n3035 & n3036;
  assign n2719 = n2718 ^ x59;
  assign n2721 = n2720 ^ n2719;
  assign n3065 = n3037 ^ n2721;
  assign n3066 = n3064 & ~n3065;
  assign n3041 = n2840 ^ x58;
  assign n3042 = n3041 ^ n2836;
  assign n3038 = n3037 ^ n2719;
  assign n3039 = ~n2721 & ~n3038;
  assign n3040 = n3039 ^ n2720;
  assign n3049 = n3042 ^ n3040;
  assign n3072 = n3066 ^ n3049;
  assign n3073 = n3061 ^ n3060;
  assign n3074 = n3059 ^ n3050;
  assign n3075 = n3058 ^ n3051;
  assign n3076 = n3057 ^ n3056;
  assign n3077 = n3053 ^ n3052;
  assign n3078 = n2978 ^ x36;
  assign n3079 = ~n3053 & ~n3078;
  assign n3080 = ~n3077 & n3079;
  assign n3081 = n3055 ^ n3054;
  assign n3082 = ~n3080 & n3081;
  assign n3083 = ~n3076 & n3082;
  assign n3084 = n3075 & ~n3083;
  assign n3085 = n3074 & n3084;
  assign n3086 = ~n3073 & ~n3085;
  assign n3087 = n3063 ^ n3062;
  assign n3088 = n3086 & ~n3087;
  assign n3089 = n3065 ^ n3064;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = n3072 & n3090;
  assign n3044 = n2843 ^ x57;
  assign n3045 = n3044 ^ n2834;
  assign n3043 = ~n3040 & n3042;
  assign n3068 = n3045 ^ n3043;
  assign n3067 = n3049 & ~n3066;
  assign n3071 = n3068 ^ n3067;
  assign n3212 = n3091 ^ n3071;
  assign n3207 = n3090 ^ n3072;
  assign n3202 = n3089 ^ n3088;
  assign n3197 = n3087 ^ n3086;
  assign n3192 = n3085 ^ n3073;
  assign n3187 = n3084 ^ n3074;
  assign n3161 = n3083 ^ n3075;
  assign n3162 = n3161 ^ x90;
  assign n3179 = n3082 ^ n3076;
  assign n3174 = n3081 ^ n3080;
  assign n3169 = n3079 ^ n3077;
  assign n3163 = x95 & n3078;
  assign n3164 = n3163 ^ x94;
  assign n3165 = n3078 ^ n3053;
  assign n3166 = n3165 ^ n3163;
  assign n3167 = n3164 & ~n3166;
  assign n3168 = n3167 ^ x94;
  assign n3170 = n3169 ^ n3168;
  assign n3171 = n3169 ^ x93;
  assign n3172 = n3170 & ~n3171;
  assign n3173 = n3172 ^ x93;
  assign n3175 = n3174 ^ n3173;
  assign n3176 = n3174 ^ x92;
  assign n3177 = ~n3175 & n3176;
  assign n3178 = n3177 ^ x92;
  assign n3180 = n3179 ^ n3178;
  assign n3181 = n3179 ^ x91;
  assign n3182 = ~n3180 & n3181;
  assign n3183 = n3182 ^ x91;
  assign n3184 = n3183 ^ n3161;
  assign n3185 = ~n3162 & n3184;
  assign n3186 = n3185 ^ x90;
  assign n3188 = n3187 ^ n3186;
  assign n3189 = n3187 ^ x89;
  assign n3190 = ~n3188 & n3189;
  assign n3191 = n3190 ^ x89;
  assign n3193 = n3192 ^ n3191;
  assign n3194 = n3192 ^ x88;
  assign n3195 = n3193 & ~n3194;
  assign n3196 = n3195 ^ x88;
  assign n3198 = n3197 ^ n3196;
  assign n3199 = n3197 ^ x87;
  assign n3200 = ~n3198 & n3199;
  assign n3201 = n3200 ^ x87;
  assign n3203 = n3202 ^ n3201;
  assign n3204 = n3202 ^ x86;
  assign n3205 = ~n3203 & n3204;
  assign n3206 = n3205 ^ x86;
  assign n3208 = n3207 ^ n3206;
  assign n3209 = n3207 ^ x85;
  assign n3210 = ~n3208 & n3209;
  assign n3211 = n3210 ^ x85;
  assign n3213 = n3212 ^ n3211;
  assign n3506 = n3213 ^ x84;
  assign n3508 = n3507 ^ n3506;
  assign n3472 = n3208 ^ x85;
  assign n3144 = n2886 ^ x48;
  assign n3471 = n2919 & n3144;
  assign n3473 = n3472 ^ n3471;
  assign n3299 = n3203 ^ x86;
  assign n3139 = n2881 ^ x49;
  assign n3298 = n2758 & ~n3139;
  assign n3300 = n3299 ^ n3298;
  assign n3130 = n2876 ^ x50;
  assign n3302 = ~n2727 & n3130;
  assign n3301 = n3198 ^ x87;
  assign n3303 = n3302 ^ n3301;
  assign n3124 = n2871 ^ x51;
  assign n3305 = n2755 & n3124;
  assign n3304 = n3193 ^ x88;
  assign n3306 = n3305 ^ n3304;
  assign n3116 = n2866 ^ x52;
  assign n3308 = n2728 & ~n3116;
  assign n3307 = n3188 ^ x89;
  assign n3309 = n3308 ^ n3307;
  assign n3111 = n2861 ^ x53;
  assign n3312 = n2729 & ~n3111;
  assign n3310 = n3183 ^ x90;
  assign n3311 = n3310 ^ n3161;
  assign n3313 = n3312 ^ n3311;
  assign n3104 = n2856 ^ x54;
  assign n3105 = n3104 ^ n2832;
  assign n3315 = ~n2730 & ~n3105;
  assign n3314 = n3180 ^ x91;
  assign n3316 = n3315 ^ n3314;
  assign n3095 = n2853 ^ x55;
  assign n3318 = n2731 & ~n3095;
  assign n3317 = n3175 ^ x92;
  assign n3319 = n3318 ^ n3317;
  assign n3321 = n3170 ^ x93;
  assign n3047 = n2848 ^ x56;
  assign n3320 = ~n2720 & ~n3047;
  assign n3322 = n3321 ^ n3320;
  assign n3324 = n2748 & ~n3045;
  assign n3323 = n3165 ^ n3164;
  assign n3325 = n3324 ^ n3323;
  assign n3327 = n3078 ^ x95;
  assign n3326 = ~n2746 & n3042;
  assign n3328 = n3327 ^ n3326;
  assign n3414 = n2719 & ~n2744;
  assign n3396 = n2956 ^ x38;
  assign n3383 = n2945 ^ x39;
  assign n3384 = n3383 ^ n2684;
  assign n3329 = n2912 ^ x42;
  assign n3330 = n3329 ^ n2828;
  assign n3331 = n2909 ^ x43;
  assign n3332 = n3331 ^ n3007;
  assign n3263 = n2894 ^ x46;
  assign n3151 = n3150 ^ n2963;
  assign n3125 = n3124 ^ n2919;
  assign n3096 = n3095 ^ n2728;
  assign n3046 = ~n3043 & n3045;
  assign n3094 = ~n3046 & ~n3047;
  assign n3101 = n3095 ^ n3094;
  assign n3102 = ~n3096 & n3101;
  assign n3103 = n3102 ^ n2728;
  assign n3110 = ~n3103 & n3105;
  assign n3117 = ~n3110 & ~n3111;
  assign n3123 = n3116 & ~n3117;
  assign n3131 = n3124 ^ n3123;
  assign n3132 = ~n3125 & n3131;
  assign n3133 = n3132 ^ n2919;
  assign n3138 = n3130 & ~n3133;
  assign n3143 = n3138 & ~n3139;
  assign n3149 = ~n3143 & ~n3144;
  assign n3264 = n3150 ^ n3149;
  assign n3265 = n3151 & ~n3264;
  assign n3266 = n3265 ^ n2963;
  assign n3275 = ~n3263 & n3266;
  assign n3276 = n2899 ^ x45;
  assign n3286 = n3275 & ~n3276;
  assign n3287 = n2904 ^ x44;
  assign n3333 = n3286 & n3287;
  assign n3334 = n3333 ^ n3331;
  assign n3335 = ~n3332 & n3334;
  assign n3336 = n3335 ^ n3007;
  assign n3337 = ~n3330 & ~n3336;
  assign n3338 = n2923 ^ x41;
  assign n3354 = ~n3337 & n3338;
  assign n3355 = n2934 ^ x40;
  assign n3382 = n3354 & ~n3355;
  assign n3393 = n3383 ^ n3382;
  assign n3394 = n3384 & n3393;
  assign n3395 = n3394 ^ n2684;
  assign n3397 = n3396 ^ n3395;
  assign n3339 = n3338 ^ n3337;
  assign n3340 = n3336 ^ n3330;
  assign n3288 = n3287 ^ n3286;
  assign n3277 = n3276 ^ n3275;
  assign n3152 = n3151 ^ n3149;
  assign n3145 = n3144 ^ n3143;
  assign n3118 = n3117 ^ n3116;
  assign n3112 = n3111 ^ n3110;
  assign n3106 = n3105 ^ n3103;
  assign n3097 = n3096 ^ n3094;
  assign n3048 = n3047 ^ n3046;
  assign n3069 = n3067 & ~n3068;
  assign n3098 = ~n3048 & n3069;
  assign n3107 = ~n3097 & ~n3098;
  assign n3113 = ~n3106 & ~n3107;
  assign n3119 = ~n3112 & n3113;
  assign n3122 = n3118 & ~n3119;
  assign n3126 = n3125 ^ n3123;
  assign n3129 = ~n3122 & ~n3126;
  assign n3134 = n3133 ^ n3130;
  assign n3137 = ~n3129 & ~n3134;
  assign n3140 = n3139 ^ n3138;
  assign n3146 = ~n3137 & n3140;
  assign n3153 = n3145 & n3146;
  assign n3262 = n3152 & n3153;
  assign n3267 = n3266 ^ n3263;
  assign n3278 = ~n3262 & n3267;
  assign n3289 = ~n3277 & ~n3278;
  assign n3341 = ~n3288 & ~n3289;
  assign n3342 = n3333 ^ n3007;
  assign n3343 = n3342 ^ n3331;
  assign n3344 = n3341 & n3343;
  assign n3345 = n3340 & n3344;
  assign n3353 = ~n3339 & ~n3345;
  assign n3356 = n3355 ^ n3354;
  assign n3381 = n3353 & ~n3356;
  assign n3385 = n3384 ^ n3382;
  assign n3398 = ~n3381 & ~n3385;
  assign n3410 = ~n3397 & n3398;
  assign n3294 = n2967 ^ x37;
  assign n3411 = n3410 ^ n3294;
  assign n3407 = ~n3395 & ~n3396;
  assign n3399 = n3398 ^ n3397;
  assign n3386 = n3385 ^ n3381;
  assign n3346 = n3345 ^ n3339;
  assign n3347 = n3344 ^ n3340;
  assign n3348 = n3343 ^ n3341;
  assign n3070 = n3069 ^ n3048;
  assign n3092 = ~n3071 & ~n3091;
  assign n3093 = ~n3070 & n3092;
  assign n3099 = n3098 ^ n3097;
  assign n3100 = n3093 & ~n3099;
  assign n3108 = n3107 ^ n3106;
  assign n3109 = n3100 & n3108;
  assign n3114 = n3113 ^ n3112;
  assign n3115 = ~n3109 & n3114;
  assign n3120 = n3119 ^ n3118;
  assign n3121 = n3115 & ~n3120;
  assign n3127 = n3126 ^ n3122;
  assign n3128 = ~n3121 & n3127;
  assign n3135 = n3134 ^ n3129;
  assign n3136 = ~n3128 & n3135;
  assign n3141 = n3140 ^ n3137;
  assign n3142 = n3136 & n3141;
  assign n3147 = n3146 ^ n3145;
  assign n3148 = n3142 & ~n3147;
  assign n3154 = n3153 ^ n3152;
  assign n3261 = n3148 & ~n3154;
  assign n3268 = n3267 ^ n3262;
  assign n3274 = n3261 & ~n3268;
  assign n3279 = n3278 ^ n3277;
  assign n3285 = ~n3274 & n3279;
  assign n3290 = n3289 ^ n3288;
  assign n3349 = ~n3285 & n3290;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = n3347 & ~n3350;
  assign n3352 = n3346 & ~n3351;
  assign n3357 = n3356 ^ n3353;
  assign n3387 = n3352 & ~n3357;
  assign n3400 = n3386 & ~n3387;
  assign n3406 = n3399 & ~n3400;
  assign n3408 = n3407 ^ n3406;
  assign n3409 = n3408 ^ x64;
  assign n3412 = n3411 ^ n3409;
  assign n3401 = n3400 ^ n3399;
  assign n3388 = n3387 ^ n3386;
  assign n3358 = n3357 ^ n3352;
  assign n3359 = n3358 ^ x67;
  assign n3373 = n3351 ^ n3346;
  assign n3368 = n3350 ^ n3347;
  assign n3360 = n3349 ^ n3348;
  assign n3361 = n3360 ^ x70;
  assign n3291 = n3290 ^ n3285;
  assign n3280 = n3279 ^ n3274;
  assign n3269 = n3268 ^ n3261;
  assign n3155 = n3154 ^ n3148;
  assign n3156 = n3155 ^ x74;
  assign n3157 = n3147 ^ n3142;
  assign n3158 = n3157 ^ x75;
  assign n3250 = n3141 ^ n3136;
  assign n3245 = n3135 ^ n3128;
  assign n3240 = n3127 ^ n3121;
  assign n3159 = n3120 ^ n3115;
  assign n3160 = n3159 ^ x79;
  assign n3232 = n3114 ^ n3109;
  assign n3227 = n3108 ^ n3100;
  assign n3222 = n3099 ^ n3093;
  assign n3217 = n3092 ^ n3070;
  assign n3214 = n3212 ^ x84;
  assign n3215 = n3213 & ~n3214;
  assign n3216 = n3215 ^ x84;
  assign n3218 = n3217 ^ n3216;
  assign n3219 = n3217 ^ x83;
  assign n3220 = ~n3218 & n3219;
  assign n3221 = n3220 ^ x83;
  assign n3223 = n3222 ^ n3221;
  assign n3224 = n3222 ^ x82;
  assign n3225 = ~n3223 & n3224;
  assign n3226 = n3225 ^ x82;
  assign n3228 = n3227 ^ n3226;
  assign n3229 = n3227 ^ x81;
  assign n3230 = n3228 & ~n3229;
  assign n3231 = n3230 ^ x81;
  assign n3233 = n3232 ^ n3231;
  assign n3234 = n3232 ^ x80;
  assign n3235 = n3233 & ~n3234;
  assign n3236 = n3235 ^ x80;
  assign n3237 = n3236 ^ n3159;
  assign n3238 = ~n3160 & n3237;
  assign n3239 = n3238 ^ x79;
  assign n3241 = n3240 ^ n3239;
  assign n3242 = n3240 ^ x78;
  assign n3243 = ~n3241 & n3242;
  assign n3244 = n3243 ^ x78;
  assign n3246 = n3245 ^ n3244;
  assign n3247 = n3245 ^ x77;
  assign n3248 = n3246 & ~n3247;
  assign n3249 = n3248 ^ x77;
  assign n3251 = n3250 ^ n3249;
  assign n3252 = n3250 ^ x76;
  assign n3253 = ~n3251 & n3252;
  assign n3254 = n3253 ^ x76;
  assign n3255 = n3254 ^ n3157;
  assign n3256 = ~n3158 & n3255;
  assign n3257 = n3256 ^ x75;
  assign n3258 = n3257 ^ n3155;
  assign n3259 = ~n3156 & n3258;
  assign n3260 = n3259 ^ x74;
  assign n3270 = n3269 ^ n3260;
  assign n3271 = n3269 ^ x73;
  assign n3272 = n3270 & ~n3271;
  assign n3273 = n3272 ^ x73;
  assign n3281 = n3280 ^ n3273;
  assign n3282 = n3280 ^ x72;
  assign n3283 = ~n3281 & n3282;
  assign n3284 = n3283 ^ x72;
  assign n3292 = n3291 ^ n3284;
  assign n3362 = n3291 ^ x71;
  assign n3363 = n3292 & ~n3362;
  assign n3364 = n3363 ^ x71;
  assign n3365 = n3364 ^ n3360;
  assign n3366 = ~n3361 & n3365;
  assign n3367 = n3366 ^ x70;
  assign n3369 = n3368 ^ n3367;
  assign n3370 = n3368 ^ x69;
  assign n3371 = n3369 & ~n3370;
  assign n3372 = n3371 ^ x69;
  assign n3374 = n3373 ^ n3372;
  assign n3375 = n3373 ^ x68;
  assign n3376 = ~n3374 & n3375;
  assign n3377 = n3376 ^ x68;
  assign n3378 = n3377 ^ n3358;
  assign n3379 = n3359 & ~n3378;
  assign n3380 = n3379 ^ x67;
  assign n3389 = n3388 ^ n3380;
  assign n3390 = n3388 ^ x66;
  assign n3391 = n3389 & ~n3390;
  assign n3392 = n3391 ^ x66;
  assign n3402 = n3401 ^ n3392;
  assign n3403 = n3401 ^ x65;
  assign n3404 = ~n3402 & n3403;
  assign n3405 = n3404 ^ x65;
  assign n3413 = n3412 ^ n3405;
  assign n3415 = n3414 ^ n3413;
  assign n3417 = n2725 & n3036;
  assign n3416 = n3402 ^ x65;
  assign n3418 = n3417 ^ n3416;
  assign n3420 = n3389 ^ x66;
  assign n3419 = n2723 & ~n2732;
  assign n3421 = n3420 ^ n3419;
  assign n3423 = n3374 ^ x68;
  assign n3424 = ~n2724 & ~n2734;
  assign n3425 = n3423 & n3424;
  assign n3422 = n2733 & n3033;
  assign n3426 = n3425 ^ n3422;
  assign n3427 = n3377 ^ x67;
  assign n3428 = n3427 ^ n3358;
  assign n3429 = n3428 ^ n3422;
  assign n3430 = n3426 & ~n3429;
  assign n3431 = n3430 ^ n3425;
  assign n3432 = n3431 ^ n3420;
  assign n3433 = ~n3421 & n3432;
  assign n3434 = n3433 ^ n3419;
  assign n3435 = n3434 ^ n3416;
  assign n3436 = n3418 & ~n3435;
  assign n3437 = n3436 ^ n3417;
  assign n3438 = n3437 ^ n3413;
  assign n3439 = ~n3415 & n3438;
  assign n3440 = n3439 ^ n3414;
  assign n3441 = n3440 ^ n3327;
  assign n3442 = n3328 & ~n3441;
  assign n3443 = n3442 ^ n3326;
  assign n3444 = n3443 ^ n3323;
  assign n3445 = ~n3325 & ~n3444;
  assign n3446 = n3445 ^ n3324;
  assign n3447 = n3446 ^ n3321;
  assign n3448 = n3322 & ~n3447;
  assign n3449 = n3448 ^ n3320;
  assign n3450 = n3449 ^ n3317;
  assign n3451 = n3319 & n3450;
  assign n3452 = n3451 ^ n3318;
  assign n3453 = n3452 ^ n3314;
  assign n3454 = n3316 & ~n3453;
  assign n3455 = n3454 ^ n3315;
  assign n3456 = n3455 ^ n3311;
  assign n3457 = ~n3313 & n3456;
  assign n3458 = n3457 ^ n3312;
  assign n3459 = n3458 ^ n3307;
  assign n3460 = ~n3309 & ~n3459;
  assign n3461 = n3460 ^ n3308;
  assign n3462 = n3461 ^ n3304;
  assign n3463 = ~n3306 & ~n3462;
  assign n3464 = n3463 ^ n3305;
  assign n3465 = n3464 ^ n3301;
  assign n3466 = n3303 & ~n3465;
  assign n3467 = n3466 ^ n3302;
  assign n3468 = n3467 ^ n3298;
  assign n3469 = ~n3300 & n3468;
  assign n3470 = n3469 ^ n3299;
  assign n3503 = n3472 ^ n3470;
  assign n3504 = n3473 & ~n3503;
  assign n3505 = n3504 ^ n3471;
  assign n3509 = n3508 ^ n3505;
  assign n3474 = n3473 ^ n3470;
  assign n3475 = n3467 ^ n3300;
  assign n3476 = n3461 ^ n3306;
  assign n3477 = n3458 ^ n3309;
  assign n3478 = n3440 ^ n3328;
  assign n3479 = n3428 ^ n3426;
  assign n3480 = n3431 ^ n3421;
  assign n3481 = n3479 & ~n3480;
  assign n3482 = n3434 ^ n3418;
  assign n3483 = n3481 & n3482;
  assign n3484 = n3437 ^ n3415;
  assign n3485 = n3483 & ~n3484;
  assign n3486 = ~n3478 & ~n3485;
  assign n3487 = n3443 ^ n3325;
  assign n3488 = n3486 & n3487;
  assign n3489 = n3446 ^ n3322;
  assign n3490 = n3488 & n3489;
  assign n3491 = n3449 ^ n3319;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = n3452 ^ n3316;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = n3455 ^ n3313;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = n3477 & ~n3496;
  assign n3498 = n3476 & ~n3497;
  assign n3499 = n3464 ^ n3303;
  assign n3500 = ~n3498 & ~n3499;
  assign n3501 = n3475 & n3500;
  assign n3502 = n3474 & ~n3501;
  assign n3510 = n3509 ^ n3502;
  assign n3511 = n3501 ^ n3474;
  assign n3512 = n3499 ^ n3498;
  assign n3513 = n3497 ^ n3476;
  assign n3514 = n3485 ^ n3478;
  assign n3515 = n3484 ^ n3483;
  assign n3516 = n3424 ^ n3423;
  assign n3517 = ~n3479 & n3516;
  assign n3518 = n3480 ^ n3479;
  assign n3519 = n3517 & ~n3518;
  assign n3520 = n3482 ^ n3481;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = n3515 & n3521;
  assign n3523 = ~n3514 & ~n3522;
  assign n3524 = n3487 ^ n3486;
  assign n3525 = n3523 & ~n3524;
  assign n3526 = n3489 ^ n3488;
  assign n3527 = ~n3525 & n3526;
  assign n3528 = n3491 ^ n3490;
  assign n3529 = n3527 & ~n3528;
  assign n3530 = n3493 ^ n3492;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = n3495 ^ n3494;
  assign n3533 = n3531 & n3532;
  assign n3534 = n3496 ^ n3477;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = n3513 & n3535;
  assign n3537 = n3512 & n3536;
  assign n3538 = n3500 ^ n3475;
  assign n3539 = n3537 & n3538;
  assign n3540 = ~n3511 & ~n3539;
  assign n3541 = ~n3510 & n3540;
  assign n3549 = ~n3502 & ~n3509;
  assign n3546 = n3218 ^ x83;
  assign n3545 = ~n2939 & n3263;
  assign n3547 = n3546 ^ n3545;
  assign n3542 = n3506 ^ n3505;
  assign n3543 = n3508 & n3542;
  assign n3544 = n3543 ^ n3507;
  assign n3548 = n3547 ^ n3544;
  assign n3550 = n3549 ^ n3548;
  assign n3551 = ~n3541 & n3550;
  assign n3557 = n3223 ^ x82;
  assign n3556 = ~n2951 & n3276;
  assign n3558 = n3557 ^ n3556;
  assign n3553 = n3546 ^ n3544;
  assign n3554 = n3547 & n3553;
  assign n3555 = n3554 ^ n3545;
  assign n3559 = n3558 ^ n3555;
  assign n3552 = n3548 & n3549;
  assign n3560 = n3559 ^ n3552;
  assign n3661 = ~n3551 & ~n3560;
  assign n3667 = n3228 ^ x81;
  assign n3666 = n2963 & ~n3287;
  assign n3668 = n3667 ^ n3666;
  assign n3663 = n3557 ^ n3555;
  assign n3664 = n3558 & ~n3663;
  assign n3665 = n3664 ^ n3556;
  assign n3669 = n3668 ^ n3665;
  assign n3662 = ~n3552 & n3559;
  assign n3670 = n3669 ^ n3662;
  assign n3872 = n3661 & ~n3670;
  assign n3831 = n3662 & ~n3669;
  assign n3799 = n3667 ^ n3665;
  assign n3800 = ~n3668 & n3799;
  assign n3801 = n3800 ^ n3666;
  assign n3797 = n2973 & n3331;
  assign n3829 = n3801 ^ n3797;
  assign n3728 = n3233 ^ x80;
  assign n3830 = n3829 ^ n3728;
  assign n3871 = n3831 ^ n3830;
  assign n3898 = n3872 ^ n3871;
  assign n3914 = x107 & ~n3898;
  assign n3798 = n3797 ^ n3728;
  assign n3802 = n3801 ^ n3728;
  assign n3803 = n3798 & n3802;
  assign n3804 = n3803 ^ n3797;
  assign n3795 = ~n2984 & ~n3330;
  assign n3723 = n3236 ^ n3160;
  assign n3796 = n3795 ^ n3723;
  assign n3833 = n3804 ^ n3796;
  assign n3832 = ~n3830 & ~n3831;
  assign n3874 = n3833 ^ n3832;
  assign n3873 = ~n3871 & n3872;
  assign n3896 = n3874 ^ n3873;
  assign n3915 = n3896 ^ x106;
  assign n3916 = ~n3914 & n3915;
  assign n3897 = ~x106 & ~n3896;
  assign n3917 = n3916 ^ n3897;
  assign n3899 = ~x107 & n3898;
  assign n3900 = ~n3897 & ~n3899;
  assign n3671 = n3670 ^ n3661;
  assign n3672 = n3671 ^ x108;
  assign n3561 = n3560 ^ n3551;
  assign n3562 = n3561 ^ x109;
  assign n3565 = n3550 ^ n3541;
  assign n3568 = ~x110 & ~n3565;
  assign n3563 = n3540 ^ n3510;
  assign n3564 = x111 & ~n3563;
  assign n3566 = n3565 ^ x110;
  assign n3567 = ~n3564 & n3566;
  assign n3569 = n3568 ^ n3567;
  assign n3918 = n3562 & n3569;
  assign n3901 = ~x109 & ~n3561;
  assign n3919 = n3918 ^ n3901;
  assign n3920 = n3919 ^ n3671;
  assign n3921 = ~n3672 & ~n3920;
  assign n3922 = n3921 ^ x108;
  assign n3570 = n3539 ^ n3511;
  assign n3571 = n3570 ^ x112;
  assign n3572 = n3538 ^ n3537;
  assign n3573 = n3572 ^ x113;
  assign n3574 = n3526 ^ n3525;
  assign n3575 = n3574 ^ x120;
  assign n3576 = n3524 ^ n3523;
  assign n3577 = n3576 ^ x121;
  assign n3578 = ~n3481 & ~n3519;
  assign n3579 = n3578 ^ n3482;
  assign n3580 = n3579 ^ x124;
  assign n3581 = n3518 ^ n3517;
  assign n3582 = n3581 ^ x125;
  assign n3583 = x127 & ~n3516;
  assign n3584 = n3583 ^ x126;
  assign n3585 = n3516 ^ n3479;
  assign n3586 = n3585 ^ n3583;
  assign n3587 = n3584 & n3586;
  assign n3588 = n3587 ^ x126;
  assign n3589 = n3588 ^ n3581;
  assign n3590 = ~n3582 & n3589;
  assign n3591 = n3590 ^ x125;
  assign n3592 = n3591 ^ n3579;
  assign n3593 = n3580 & ~n3592;
  assign n3594 = n3593 ^ x124;
  assign n3595 = n3521 ^ n3515;
  assign n3596 = ~x123 & n3595;
  assign n3597 = n3522 ^ n3514;
  assign n3598 = ~x122 & ~n3597;
  assign n3599 = ~n3596 & ~n3598;
  assign n3600 = n3594 & n3599;
  assign n3601 = x123 & ~n3595;
  assign n3602 = n3597 ^ x122;
  assign n3603 = ~n3601 & n3602;
  assign n3604 = n3603 ^ n3598;
  assign n3605 = ~n3600 & n3604;
  assign n3606 = n3605 ^ n3576;
  assign n3607 = ~n3577 & ~n3606;
  assign n3608 = n3607 ^ x121;
  assign n3609 = n3608 ^ n3574;
  assign n3610 = n3575 & ~n3609;
  assign n3611 = n3610 ^ x120;
  assign n3612 = n3532 ^ n3531;
  assign n3613 = ~x117 & ~n3612;
  assign n3614 = n3530 ^ n3529;
  assign n3615 = ~x118 & ~n3614;
  assign n3616 = n3528 ^ n3527;
  assign n3617 = ~x119 & ~n3616;
  assign n3618 = ~n3615 & ~n3617;
  assign n3619 = n3534 ^ n3533;
  assign n3620 = ~x116 & n3619;
  assign n3621 = n3618 & ~n3620;
  assign n3622 = ~n3613 & n3621;
  assign n3623 = n3611 & n3622;
  assign n3624 = n3619 ^ x116;
  assign n3625 = n3612 ^ x117;
  assign n3626 = x119 & n3616;
  assign n3627 = n3614 ^ x118;
  assign n3628 = ~n3626 & n3627;
  assign n3629 = n3628 ^ n3615;
  assign n3630 = n3629 ^ n3612;
  assign n3631 = n3625 & n3630;
  assign n3632 = n3631 ^ x117;
  assign n3633 = ~n3624 & n3632;
  assign n3634 = n3633 ^ n3624;
  assign n3635 = n3634 ^ n3620;
  assign n3636 = ~n3623 & ~n3635;
  assign n3637 = n3535 ^ n3513;
  assign n3638 = ~x115 & n3637;
  assign n3639 = n3536 ^ n3512;
  assign n3640 = ~x114 & n3639;
  assign n3641 = ~n3638 & ~n3640;
  assign n3642 = ~n3636 & n3641;
  assign n3643 = x115 & ~n3637;
  assign n3644 = n3639 ^ x114;
  assign n3645 = ~n3643 & ~n3644;
  assign n3646 = n3645 ^ n3640;
  assign n3647 = ~n3642 & n3646;
  assign n3648 = n3647 ^ n3572;
  assign n3649 = ~n3573 & ~n3648;
  assign n3650 = n3649 ^ x113;
  assign n3651 = n3650 ^ n3570;
  assign n3652 = n3571 & ~n3651;
  assign n3653 = n3652 ^ x112;
  assign n3654 = ~x111 & n3563;
  assign n3655 = ~n3568 & ~n3654;
  assign n3902 = ~x108 & n3671;
  assign n3903 = n3655 & ~n3902;
  assign n3904 = ~n3901 & n3903;
  assign n4098 = n3653 & n3904;
  assign n4099 = ~n3922 & ~n4098;
  assign n4402 = n3900 & ~n4099;
  assign n4403 = n3917 & ~n4402;
  assign n3805 = n3804 ^ n3723;
  assign n3806 = ~n3796 & ~n3805;
  assign n3807 = n3806 ^ n3795;
  assign n3793 = ~n2995 & ~n3338;
  assign n3712 = n3241 ^ x78;
  assign n3794 = n3793 ^ n3712;
  assign n3835 = n3807 ^ n3794;
  assign n3834 = n3832 & ~n3833;
  assign n3876 = n3835 ^ n3834;
  assign n3875 = n3873 & n3874;
  assign n3905 = n3876 ^ n3875;
  assign n4401 = n3905 ^ x105;
  assign n4404 = n4403 ^ n4401;
  assign n4097 = n3898 ^ x107;
  assign n4112 = n4099 ^ n3898;
  assign n4113 = ~n4097 & ~n4112;
  assign n4114 = n4113 ^ x107;
  assign n4115 = n4114 ^ n3915;
  assign n3973 = n3369 ^ x69;
  assign n4108 = n3013 ^ n2682;
  assign n4109 = ~n3973 & n4108;
  assign n4110 = n4109 ^ n2682;
  assign n4397 = n4115 ^ n4110;
  assign n4100 = n4099 ^ n4097;
  assign n3656 = n3653 & n3655;
  assign n3657 = n3569 & ~n3656;
  assign n3658 = n3657 ^ n3561;
  assign n3659 = n3562 & n3658;
  assign n3660 = n3659 ^ x109;
  assign n3673 = n3672 ^ n3660;
  assign n3293 = n3292 ^ x71;
  assign n3295 = n3294 ^ n3025;
  assign n3296 = ~n3293 & n3295;
  assign n3297 = n3296 ^ n3025;
  assign n3674 = n3673 ^ n3297;
  assign n3679 = n3657 ^ n3562;
  assign n3675 = n3281 ^ x72;
  assign n3676 = n3396 ^ n3007;
  assign n3677 = n3675 & n3676;
  assign n3678 = n3677 ^ n3007;
  assign n3680 = n3679 ^ n3678;
  assign n3685 = n3563 ^ x111;
  assign n4079 = n3653 ^ n3563;
  assign n4080 = ~n3685 & n4079;
  assign n4081 = n4080 ^ x111;
  assign n4082 = n4081 ^ x110;
  assign n4083 = n4082 ^ n3565;
  assign n3686 = n3685 ^ n3653;
  assign n3681 = n3257 ^ n3156;
  assign n3682 = n3355 ^ n2984;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = n3683 ^ n2984;
  assign n3687 = n3686 ^ n3684;
  assign n3692 = n3650 ^ n3571;
  assign n3688 = n3254 ^ n3158;
  assign n3689 = n3338 ^ n2973;
  assign n3690 = ~n3688 & n3689;
  assign n3691 = n3690 ^ n2973;
  assign n3693 = n3692 ^ n3691;
  assign n3698 = n3647 ^ n3573;
  assign n3694 = n3251 ^ x76;
  assign n3695 = n3330 ^ n2963;
  assign n3696 = n3694 & ~n3695;
  assign n3697 = n3696 ^ n2963;
  assign n3699 = n3698 ^ n3697;
  assign n3704 = n3637 ^ x115;
  assign n3705 = n3637 ^ n3636;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = n3706 ^ x115;
  assign n3708 = n3707 ^ n3644;
  assign n3700 = n3246 ^ x77;
  assign n3701 = n3331 ^ n2951;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = n3702 ^ n2951;
  assign n3709 = n3708 ^ n3703;
  assign n3713 = n3287 ^ n2939;
  assign n3714 = n3712 & n3713;
  assign n3715 = n3714 ^ n2939;
  assign n3710 = n3636 ^ x115;
  assign n3711 = n3710 ^ n3637;
  assign n3716 = n3715 ^ n3711;
  assign n3724 = n3276 ^ n2930;
  assign n3725 = ~n3723 & ~n3724;
  assign n3726 = n3725 ^ n2930;
  assign n3717 = n3611 & n3618;
  assign n3718 = n3629 & ~n3717;
  assign n3719 = n3718 ^ n3612;
  assign n3720 = n3625 & n3719;
  assign n3721 = n3720 ^ x117;
  assign n3722 = n3721 ^ n3624;
  assign n3727 = n3726 ^ n3722;
  assign n3732 = n3718 ^ n3625;
  assign n3729 = n3263 ^ n2919;
  assign n3730 = ~n3728 & n3729;
  assign n3731 = n3730 ^ n2919;
  assign n3733 = n3732 ^ n3731;
  assign n3738 = n3150 ^ n2758;
  assign n3739 = ~n3667 & n3738;
  assign n3740 = n3739 ^ n2758;
  assign n3734 = n3616 ^ x119;
  assign n3735 = n3611 & n3734;
  assign n3736 = n3735 ^ n3626;
  assign n3737 = n3736 ^ n3627;
  assign n3741 = n3740 ^ n3737;
  assign n3743 = n3144 ^ n2727;
  assign n3744 = n3557 & ~n3743;
  assign n3745 = n3744 ^ n2727;
  assign n3742 = n3734 ^ n3611;
  assign n3746 = n3745 ^ n3742;
  assign n3750 = n3608 ^ n3575;
  assign n3747 = n3139 ^ n2755;
  assign n3748 = n3546 & ~n3747;
  assign n3749 = n3748 ^ n2755;
  assign n3751 = n3750 ^ n3749;
  assign n4041 = n3605 ^ n3577;
  assign n3755 = ~n3596 & ~n3601;
  assign n3756 = n3594 & n3755;
  assign n3757 = n3756 ^ n3601;
  assign n3758 = n3757 ^ n3602;
  assign n3752 = n3124 ^ n2729;
  assign n3753 = n3472 & n3752;
  assign n3754 = n3753 ^ n2729;
  assign n3759 = n3758 ^ n3754;
  assign n4030 = n3755 ^ n3594;
  assign n3762 = n3111 ^ n2731;
  assign n3763 = n3301 & ~n3762;
  assign n3764 = n3763 ^ n2731;
  assign n3760 = n3591 ^ x124;
  assign n3761 = n3760 ^ n3579;
  assign n3765 = n3764 ^ n3761;
  assign n3769 = n3588 ^ x125;
  assign n3770 = n3769 ^ n3581;
  assign n3766 = n3105 ^ n2720;
  assign n3767 = ~n3304 & ~n3766;
  assign n3768 = n3767 ^ n2720;
  assign n3771 = n3770 ^ n3768;
  assign n3773 = n3095 ^ n2748;
  assign n3774 = n3307 & n3773;
  assign n3775 = n3774 ^ n2748;
  assign n3772 = n3585 ^ n3584;
  assign n3776 = n3775 ^ n3772;
  assign n3778 = n3047 ^ n2746;
  assign n3779 = ~n3311 & n3778;
  assign n3780 = n3779 ^ n2746;
  assign n3777 = n3516 ^ x127;
  assign n3781 = n3780 ^ n3777;
  assign n3782 = n3045 ^ n2744;
  assign n3783 = n3314 & n3782;
  assign n3784 = n3783 ^ n2744;
  assign n3972 = ~n2735 & n3028;
  assign n3974 = n3973 ^ n3972;
  assign n3863 = x31 & ~n3012;
  assign n3862 = n3364 ^ n3361;
  assign n3864 = n3863 ^ n3862;
  assign n3855 = ~n2711 & n3015;
  assign n3856 = n3855 ^ n3293;
  assign n3848 = ~n2690 & n3013;
  assign n3849 = n3848 ^ n3675;
  assign n3824 = n2684 & ~n3078;
  assign n3823 = n3270 ^ x73;
  assign n3825 = n3824 ^ n3823;
  assign n3785 = n2682 & n3294;
  assign n3786 = n3785 ^ n3681;
  assign n3787 = n2686 & n3396;
  assign n3788 = n3787 ^ n3688;
  assign n3789 = ~n3025 & n3383;
  assign n3790 = n3789 ^ n3694;
  assign n3791 = ~n3007 & n3355;
  assign n3792 = n3791 ^ n3700;
  assign n3808 = n3807 ^ n3712;
  assign n3809 = ~n3794 & ~n3808;
  assign n3810 = n3809 ^ n3793;
  assign n3811 = n3810 ^ n3700;
  assign n3812 = n3792 & ~n3811;
  assign n3813 = n3812 ^ n3791;
  assign n3814 = n3813 ^ n3694;
  assign n3815 = ~n3790 & n3814;
  assign n3816 = n3815 ^ n3789;
  assign n3817 = n3816 ^ n3688;
  assign n3818 = ~n3788 & ~n3817;
  assign n3819 = n3818 ^ n3787;
  assign n3820 = n3819 ^ n3681;
  assign n3821 = ~n3786 & n3820;
  assign n3822 = n3821 ^ n3785;
  assign n3845 = n3823 ^ n3822;
  assign n3846 = n3825 & n3845;
  assign n3847 = n3846 ^ n3824;
  assign n3852 = n3847 ^ n3675;
  assign n3853 = ~n3849 & n3852;
  assign n3854 = n3853 ^ n3848;
  assign n3859 = n3855 ^ n3854;
  assign n3860 = n3856 & ~n3859;
  assign n3861 = n3860 ^ n3854;
  assign n3969 = n3862 ^ n3861;
  assign n3970 = n3864 & ~n3969;
  assign n3971 = n3970 ^ n3863;
  assign n3975 = n3974 ^ n3971;
  assign n3850 = n3849 ^ n3847;
  assign n3826 = n3825 ^ n3822;
  assign n3827 = n3819 ^ n3786;
  assign n3828 = n3816 ^ n3788;
  assign n3836 = n3834 & n3835;
  assign n3837 = n3810 ^ n3791;
  assign n3838 = n3837 ^ n3700;
  assign n3839 = n3836 & n3838;
  assign n3840 = n3813 ^ n3790;
  assign n3841 = n3839 & ~n3840;
  assign n3842 = ~n3828 & n3841;
  assign n3843 = ~n3827 & ~n3842;
  assign n3844 = ~n3826 & ~n3843;
  assign n3867 = n3850 ^ n3844;
  assign n3868 = n3843 ^ n3826;
  assign n3869 = n3840 ^ n3839;
  assign n3870 = n3838 ^ n3836;
  assign n3877 = n3875 & ~n3876;
  assign n3878 = n3870 & ~n3877;
  assign n3879 = n3869 & ~n3878;
  assign n3880 = n3841 ^ n3828;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = n3842 ^ n3827;
  assign n3883 = ~n3881 & n3882;
  assign n3884 = n3868 & ~n3883;
  assign n3885 = ~n3867 & n3884;
  assign n3857 = n3856 ^ n3854;
  assign n3851 = n3844 & ~n3850;
  assign n3886 = n3857 ^ n3851;
  assign n3887 = ~n3885 & n3886;
  assign n3865 = n3864 ^ n3861;
  assign n3964 = n3887 ^ n3865;
  assign n3858 = n3851 & ~n3857;
  assign n3965 = n3887 ^ n3858;
  assign n3966 = ~n3964 & n3965;
  assign n3967 = n3966 ^ n3865;
  assign n3968 = n3967 ^ x96;
  assign n3976 = n3975 ^ n3968;
  assign n3866 = n3865 ^ n3858;
  assign n3888 = n3887 ^ n3866;
  assign n3889 = n3888 ^ x97;
  assign n3890 = n3886 ^ n3885;
  assign n3891 = n3890 ^ x98;
  assign n3892 = n3884 ^ n3867;
  assign n3893 = n3892 ^ x99;
  assign n3950 = n3883 ^ n3868;
  assign n3894 = n3882 ^ n3881;
  assign n3895 = n3894 ^ x101;
  assign n3906 = ~x105 & n3905;
  assign n3907 = n3877 ^ n3870;
  assign n3908 = ~x104 & ~n3907;
  assign n3909 = ~n3906 & ~n3908;
  assign n3910 = n3904 & n3909;
  assign n3911 = n3900 & n3910;
  assign n3912 = n3653 & n3911;
  assign n3913 = n3907 ^ x104;
  assign n3923 = n3900 & n3922;
  assign n3924 = x105 & ~n3905;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = n3917 & n3925;
  assign n3927 = n3926 ^ n3907;
  assign n3928 = n3927 ^ n3907;
  assign n3929 = n3907 ^ n3906;
  assign n3930 = n3929 ^ n3907;
  assign n3931 = ~n3928 & ~n3930;
  assign n3932 = n3931 ^ n3907;
  assign n3933 = n3913 & ~n3932;
  assign n3934 = n3933 ^ x104;
  assign n3935 = ~n3912 & ~n3934;
  assign n3936 = n3878 ^ n3869;
  assign n3937 = ~x103 & n3936;
  assign n3938 = n3880 ^ n3879;
  assign n3939 = ~x102 & n3938;
  assign n3940 = ~n3937 & ~n3939;
  assign n3941 = ~n3935 & n3940;
  assign n3942 = x103 & ~n3936;
  assign n3943 = n3938 ^ x102;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = n3944 ^ n3939;
  assign n3946 = ~n3941 & n3945;
  assign n3947 = n3946 ^ n3894;
  assign n3948 = ~n3895 & ~n3947;
  assign n3949 = n3948 ^ x101;
  assign n3951 = n3950 ^ n3949;
  assign n3952 = n3950 ^ x100;
  assign n3953 = ~n3951 & n3952;
  assign n3954 = n3953 ^ x100;
  assign n3955 = n3954 ^ n3892;
  assign n3956 = n3893 & ~n3955;
  assign n3957 = n3956 ^ x99;
  assign n3958 = n3957 ^ n3890;
  assign n3959 = ~n3891 & n3958;
  assign n3960 = n3959 ^ x98;
  assign n3961 = n3960 ^ n3888;
  assign n3962 = n3889 & ~n3961;
  assign n3963 = n3962 ^ x97;
  assign n3977 = n3976 ^ n3963;
  assign n3978 = ~n3784 & n3977;
  assign n3979 = n3978 ^ n3780;
  assign n3980 = n3781 & n3979;
  assign n3981 = n3980 ^ n3777;
  assign n3982 = n3981 ^ n3772;
  assign n3983 = n3982 ^ n3772;
  assign n3987 = n3960 ^ n3889;
  assign n3984 = n3042 ^ n2725;
  assign n3985 = n3317 & n3984;
  assign n3986 = n3985 ^ n2725;
  assign n3988 = n3987 ^ n3986;
  assign n4003 = n2732 ^ n2719;
  assign n4004 = ~n3321 & ~n4003;
  assign n4005 = n4004 ^ n2732;
  assign n3991 = n3036 ^ n2733;
  assign n3992 = n3323 & n3991;
  assign n3993 = n3992 ^ n2733;
  assign n3989 = n3954 ^ x99;
  assign n3990 = n3989 ^ n3892;
  assign n3994 = n3993 ^ n3990;
  assign n3995 = n2734 ^ n2723;
  assign n3996 = n3327 & ~n3995;
  assign n3997 = n3996 ^ n2734;
  assign n3998 = n3951 ^ x100;
  assign n3999 = ~n3997 & n3998;
  assign n4000 = n3999 ^ n3990;
  assign n4001 = ~n3994 & n4000;
  assign n4002 = n4001 ^ n3999;
  assign n4006 = n4005 ^ n4002;
  assign n4007 = n3957 ^ n3891;
  assign n4008 = n4007 ^ n4002;
  assign n4009 = ~n4006 & n4008;
  assign n4010 = n4009 ^ n4005;
  assign n4011 = n4010 ^ n3986;
  assign n4012 = n3988 & n4011;
  assign n4013 = n4012 ^ n3987;
  assign n4014 = n3784 & ~n3977;
  assign n4015 = n4013 & ~n4014;
  assign n4016 = n3777 & n3780;
  assign n4017 = n4015 & ~n4016;
  assign n4018 = n4017 ^ n3772;
  assign n4019 = n4018 ^ n3772;
  assign n4020 = n3983 & ~n4019;
  assign n4021 = n4020 ^ n3772;
  assign n4022 = n3776 & ~n4021;
  assign n4023 = n4022 ^ n3775;
  assign n4024 = n4023 ^ n3770;
  assign n4025 = ~n3771 & ~n4024;
  assign n4026 = n4025 ^ n3768;
  assign n4027 = n4026 ^ n3761;
  assign n4028 = n3765 & ~n4027;
  assign n4029 = n4028 ^ n3764;
  assign n4031 = n4030 ^ n4029;
  assign n4032 = n3116 ^ n2730;
  assign n4033 = n3299 & n4032;
  assign n4034 = n4033 ^ n2730;
  assign n4035 = n4034 ^ n4030;
  assign n4036 = ~n4031 & ~n4035;
  assign n4037 = n4036 ^ n4034;
  assign n4038 = n4037 ^ n3758;
  assign n4039 = n3759 & n4038;
  assign n4040 = n4039 ^ n3754;
  assign n4042 = n4041 ^ n4040;
  assign n4043 = n3130 ^ n2728;
  assign n4044 = ~n3506 & ~n4043;
  assign n4045 = n4044 ^ n2728;
  assign n4046 = n4045 ^ n4041;
  assign n4047 = ~n4042 & ~n4046;
  assign n4048 = n4047 ^ n4045;
  assign n4049 = n4048 ^ n3750;
  assign n4050 = n3751 & n4049;
  assign n4051 = n4050 ^ n3749;
  assign n4052 = n4051 ^ n3742;
  assign n4053 = ~n3746 & ~n4052;
  assign n4054 = n4053 ^ n3745;
  assign n4055 = n4054 ^ n3737;
  assign n4056 = ~n3741 & n4055;
  assign n4057 = n4056 ^ n3740;
  assign n4058 = n4057 ^ n3732;
  assign n4059 = ~n3733 & ~n4058;
  assign n4060 = n4059 ^ n3731;
  assign n4061 = n4060 ^ n3722;
  assign n4062 = n3727 & n4061;
  assign n4063 = n4062 ^ n3726;
  assign n4064 = n4063 ^ n3711;
  assign n4065 = ~n3716 & n4064;
  assign n4066 = n4065 ^ n3715;
  assign n4067 = n4066 ^ n3708;
  assign n4068 = n3709 & ~n4067;
  assign n4069 = n4068 ^ n3703;
  assign n4070 = n4069 ^ n3698;
  assign n4071 = n3699 & n4070;
  assign n4072 = n4071 ^ n3697;
  assign n4073 = n4072 ^ n3692;
  assign n4074 = ~n3693 & ~n4073;
  assign n4075 = n4074 ^ n3691;
  assign n4076 = n4075 ^ n3684;
  assign n4077 = n3687 & ~n4076;
  assign n4078 = n4077 ^ n3686;
  assign n4084 = n4083 ^ n4078;
  assign n4085 = n3383 ^ n2995;
  assign n4086 = ~n3823 & n4085;
  assign n4087 = n4086 ^ n2995;
  assign n4088 = n4087 ^ n4083;
  assign n4089 = n4084 & n4088;
  assign n4090 = n4089 ^ n4087;
  assign n4091 = n4090 ^ n3678;
  assign n4092 = ~n3680 & ~n4091;
  assign n4093 = n4092 ^ n3679;
  assign n4094 = n4093 ^ n3673;
  assign n4095 = ~n3674 & ~n4094;
  assign n4096 = n4095 ^ n3297;
  assign n4101 = n4100 ^ n4096;
  assign n4102 = n3078 ^ n2686;
  assign n4103 = ~n3862 & ~n4102;
  assign n4104 = n4103 ^ n2686;
  assign n4105 = n4104 ^ n4100;
  assign n4106 = ~n4101 & n4105;
  assign n4107 = n4106 ^ n4104;
  assign n4398 = n4115 ^ n4107;
  assign n4399 = n4397 & ~n4398;
  assign n4400 = n4399 ^ n4110;
  assign n4405 = n4404 ^ n4400;
  assign n4394 = n3015 ^ n2684;
  assign n4395 = n3423 & ~n4394;
  assign n4396 = n4395 ^ n2684;
  assign n4406 = n4405 ^ n4396;
  assign n4111 = n4110 ^ n4107;
  assign n4116 = n4115 ^ n4111;
  assign n4117 = n4104 ^ n4101;
  assign n4118 = n4093 ^ n3297;
  assign n4119 = n4118 ^ n3673;
  assign n4120 = n4090 ^ n3680;
  assign n4121 = n4072 ^ n3693;
  assign n4122 = n4075 ^ n3687;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = n4087 ^ n4084;
  assign n4125 = ~n4123 & n4124;
  assign n4126 = n4120 & n4125;
  assign n4127 = ~n4119 & n4126;
  assign n4128 = n4117 & ~n4127;
  assign n4407 = n4116 & n4128;
  assign n4441 = n4406 & ~n4407;
  assign n4436 = ~n4401 & ~n4403;
  assign n4437 = n4436 ^ n3924;
  assign n4438 = n4437 ^ n3913;
  assign n4433 = n4404 ^ n4396;
  assign n4434 = ~n4405 & ~n4433;
  assign n4435 = n4434 ^ n4396;
  assign n4439 = n4438 ^ n4435;
  assign n4430 = n3012 ^ n2690;
  assign n4431 = n3428 & ~n4430;
  assign n4432 = n4431 ^ n2690;
  assign n4440 = n4439 ^ n4432;
  assign n4442 = n4441 ^ n4440;
  assign n4129 = n4128 ^ n4116;
  assign n4130 = n4127 ^ n4117;
  assign n4131 = n4126 ^ n4119;
  assign n4132 = n4125 ^ n4120;
  assign n4133 = n4060 ^ n3726;
  assign n4134 = n4133 ^ n3722;
  assign n4136 = n4054 ^ n3741;
  assign n4137 = n4051 ^ n3746;
  assign n4138 = n4026 ^ n3765;
  assign n4139 = ~n3978 & ~n4015;
  assign n4140 = n4139 ^ n3780;
  assign n4141 = n3781 & ~n4140;
  assign n4142 = n4141 ^ n3777;
  assign n4143 = n4142 ^ n3776;
  assign n4144 = n4142 ^ n3775;
  assign n4145 = n3776 & ~n4144;
  assign n4146 = n4145 ^ n3772;
  assign n4147 = n4146 ^ n3771;
  assign n4148 = n4143 & ~n4147;
  assign n4149 = n4138 & ~n4148;
  assign n4150 = n4034 ^ n4031;
  assign n4151 = n4149 & ~n4150;
  assign n4152 = n4037 ^ n3759;
  assign n4153 = n4151 & ~n4152;
  assign n4154 = n4045 ^ n4042;
  assign n4155 = ~n4153 & n4154;
  assign n4156 = n4048 ^ n3751;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4137 & n4157;
  assign n4159 = ~n4136 & ~n4158;
  assign n4135 = n4057 ^ n3733;
  assign n4160 = n4159 ^ n4135;
  assign n4161 = n4158 ^ n4136;
  assign n4162 = n4156 ^ n4155;
  assign n4163 = n4148 ^ n4138;
  assign n4164 = n4139 ^ n3781;
  assign n4168 = n3998 ^ n3997;
  assign n4169 = n3999 ^ n3993;
  assign n4170 = n4169 ^ n3990;
  assign n4171 = ~n4168 & n4170;
  assign n4172 = n4007 ^ n4006;
  assign n4173 = n4171 & n4172;
  assign n4174 = n4010 ^ n3988;
  assign n4175 = ~n4173 & n4174;
  assign n4176 = ~n4164 & ~n4175;
  assign n4165 = n3977 ^ n3784;
  assign n4166 = n4165 ^ n4013;
  assign n4167 = ~n4164 & ~n4166;
  assign n4177 = n4176 ^ n4167;
  assign n4178 = n4147 ^ n4143;
  assign n4179 = n4178 ^ n4167;
  assign n4180 = ~n4167 & n4179;
  assign n4181 = n4180 ^ n4167;
  assign n4182 = n4177 & ~n4181;
  assign n4183 = n4182 ^ n4180;
  assign n4184 = n4183 ^ n4167;
  assign n4185 = n4184 ^ n4178;
  assign n4186 = n4147 & n4185;
  assign n4187 = n4186 ^ n4178;
  assign n4188 = n4163 & ~n4187;
  assign n4189 = n4150 ^ n4149;
  assign n4190 = ~n4188 & ~n4189;
  assign n4191 = n4152 ^ n4151;
  assign n4192 = n4190 & ~n4191;
  assign n4193 = n4154 ^ n4153;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n4162 & n4194;
  assign n4196 = n4157 ^ n4137;
  assign n4197 = n4195 & n4196;
  assign n4198 = n4161 & n4197;
  assign n4199 = n4198 ^ n4159;
  assign n4200 = ~n4160 & n4199;
  assign n4201 = n4200 ^ n4159;
  assign n4202 = ~n4134 & n4201;
  assign n4203 = n4063 ^ n3716;
  assign n4204 = n4202 & ~n4203;
  assign n4205 = n4066 ^ n3709;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = n4069 ^ n3699;
  assign n4208 = n4206 & ~n4207;
  assign n4209 = n4121 & n4208;
  assign n4210 = n4122 ^ n4121;
  assign n4211 = n4209 & n4210;
  assign n4212 = n4124 ^ n4123;
  assign n4213 = n4211 & n4212;
  assign n4214 = n4132 & ~n4213;
  assign n4215 = n4131 & ~n4214;
  assign n4216 = n4130 & ~n4215;
  assign n4393 = n4129 & ~n4216;
  assign n4408 = n4407 ^ n4406;
  assign n4429 = ~n4393 & ~n4408;
  assign n4443 = n4442 ^ n4429;
  assign n4444 = n4443 ^ x131;
  assign n4409 = n4408 ^ n4393;
  assign n4410 = n4409 ^ x132;
  assign n4217 = n4216 ^ n4129;
  assign n4218 = n4217 ^ x133;
  assign n4219 = n4213 ^ n4132;
  assign n4220 = n4219 ^ x136;
  assign n4223 = n4210 ^ n4209;
  assign n4226 = ~x138 & ~n4223;
  assign n4221 = n4208 ^ n4121;
  assign n4222 = x139 & n4221;
  assign n4224 = n4223 ^ x138;
  assign n4225 = ~n4222 & n4224;
  assign n4227 = n4226 ^ n4225;
  assign n4228 = ~x139 & ~n4221;
  assign n4229 = ~n4226 & ~n4228;
  assign n4230 = n4207 ^ n4206;
  assign n4232 = n4230 ^ x140;
  assign n4233 = n4205 ^ n4204;
  assign n4234 = n4233 ^ x141;
  assign n4235 = n4203 ^ n4202;
  assign n4236 = n4235 ^ x142;
  assign n4237 = n4198 ^ n4135;
  assign n4238 = n4159 ^ n4134;
  assign n4239 = n4238 ^ n4198;
  assign n4240 = n4239 ^ n4134;
  assign n4241 = n4237 & n4240;
  assign n4242 = n4241 ^ n4238;
  assign n4243 = x143 & n4242;
  assign n4244 = n4243 ^ n4235;
  assign n4245 = n4236 & ~n4244;
  assign n4246 = n4245 ^ x142;
  assign n4247 = n4246 ^ n4233;
  assign n4248 = n4234 & ~n4247;
  assign n4249 = n4248 ^ x141;
  assign n4250 = ~n4232 & n4249;
  assign n4251 = n4250 ^ n4232;
  assign n4231 = ~x140 & n4230;
  assign n4252 = n4251 ^ n4231;
  assign n4253 = n4229 & n4252;
  assign n4254 = n4212 ^ n4211;
  assign n4255 = x137 & n4254;
  assign n4256 = ~n4253 & ~n4255;
  assign n4257 = n4227 & n4256;
  assign n4258 = n4257 ^ n4219;
  assign n4259 = n4258 ^ n4219;
  assign n4260 = ~x137 & ~n4254;
  assign n4261 = n4260 ^ n4219;
  assign n4262 = n4261 ^ n4219;
  assign n4263 = ~n4259 & ~n4262;
  assign n4264 = n4263 ^ n4219;
  assign n4265 = n4220 & ~n4264;
  assign n4266 = n4265 ^ x136;
  assign n4267 = n4215 ^ n4130;
  assign n4268 = ~x134 & ~n4267;
  assign n4269 = n4214 ^ n4131;
  assign n4270 = ~x135 & n4269;
  assign n4271 = ~n4268 & ~n4270;
  assign n4272 = n4266 & n4271;
  assign n4273 = n4272 ^ n4217;
  assign n4274 = n4273 ^ n4217;
  assign n4275 = x135 & ~n4269;
  assign n4276 = n4267 ^ x134;
  assign n4277 = ~n4275 & n4276;
  assign n4278 = n4277 ^ n4268;
  assign n4279 = n4278 ^ n4217;
  assign n4280 = n4279 ^ n4217;
  assign n4281 = ~n4274 & n4280;
  assign n4282 = n4281 ^ n4217;
  assign n4283 = ~n4218 & ~n4282;
  assign n4284 = n4283 ^ x133;
  assign n4422 = n4409 ^ n4284;
  assign n4423 = ~n4410 & n4422;
  assign n4424 = n4423 ^ x132;
  assign n4285 = n4166 & n4175;
  assign n4286 = ~n4164 & ~n4285;
  assign n4287 = n4143 & n4286;
  assign n4288 = n4287 ^ n4178;
  assign n4289 = n4288 ^ x152;
  assign n4290 = n4286 ^ n4143;
  assign n4291 = n4290 ^ x153;
  assign n4292 = n4285 ^ n4164;
  assign n4293 = n4292 ^ x154;
  assign n4294 = n4175 ^ n4166;
  assign n4295 = n4294 ^ x155;
  assign n4296 = n4174 ^ n4173;
  assign n4297 = n4296 ^ x156;
  assign n4298 = n4172 ^ n4171;
  assign n4299 = n4298 ^ x157;
  assign n4300 = x159 & n4168;
  assign n4301 = n4300 ^ x158;
  assign n4302 = n4170 ^ n4168;
  assign n4303 = n4302 ^ n4300;
  assign n4304 = n4301 & n4303;
  assign n4305 = n4304 ^ x158;
  assign n4306 = n4305 ^ n4298;
  assign n4307 = n4299 & ~n4306;
  assign n4308 = n4307 ^ x157;
  assign n4309 = n4308 ^ n4296;
  assign n4310 = n4297 & ~n4309;
  assign n4311 = n4310 ^ x156;
  assign n4312 = n4311 ^ n4294;
  assign n4313 = ~n4295 & n4312;
  assign n4314 = n4313 ^ x155;
  assign n4315 = n4314 ^ n4292;
  assign n4316 = n4293 & ~n4315;
  assign n4317 = n4316 ^ x154;
  assign n4318 = n4317 ^ n4290;
  assign n4319 = n4291 & ~n4318;
  assign n4320 = n4319 ^ x153;
  assign n4321 = n4320 ^ n4288;
  assign n4322 = ~n4289 & n4321;
  assign n4323 = n4322 ^ x152;
  assign n4324 = n4196 ^ n4195;
  assign n4325 = ~x146 & n4324;
  assign n4326 = n4194 ^ n4162;
  assign n4327 = ~x147 & ~n4326;
  assign n4328 = ~n4325 & ~n4327;
  assign n4329 = n4191 ^ n4190;
  assign n4330 = ~x149 & n4329;
  assign n4331 = n4193 ^ n4192;
  assign n4332 = ~x148 & n4331;
  assign n4333 = n4189 ^ n4188;
  assign n4334 = ~x150 & ~n4333;
  assign n4335 = n4187 ^ n4163;
  assign n4336 = ~x151 & ~n4335;
  assign n4337 = ~n4334 & ~n4336;
  assign n4338 = ~n4332 & n4337;
  assign n4339 = ~n4330 & n4338;
  assign n4340 = n4197 ^ n4161;
  assign n4341 = ~x145 & n4340;
  assign n4342 = n4198 ^ n4160;
  assign n4343 = ~x144 & ~n4342;
  assign n4344 = ~n4341 & ~n4343;
  assign n4345 = n4339 & n4344;
  assign n4346 = n4328 & n4345;
  assign n4347 = n4323 & n4346;
  assign n4348 = n4342 ^ x144;
  assign n4349 = x147 & n4326;
  assign n4350 = n4324 ^ x146;
  assign n4351 = ~n4349 & ~n4350;
  assign n4352 = n4351 ^ n4325;
  assign n4353 = x145 & ~n4340;
  assign n4354 = n4331 ^ x148;
  assign n4355 = n4329 ^ x149;
  assign n4356 = x151 & n4335;
  assign n4357 = n4333 ^ x150;
  assign n4358 = ~n4356 & n4357;
  assign n4359 = n4358 ^ n4334;
  assign n4360 = n4359 ^ n4329;
  assign n4361 = ~n4355 & ~n4360;
  assign n4362 = n4361 ^ x149;
  assign n4363 = ~n4354 & n4362;
  assign n4364 = n4363 ^ n4354;
  assign n4365 = n4364 ^ n4332;
  assign n4366 = n4328 & n4365;
  assign n4367 = ~n4353 & ~n4366;
  assign n4368 = n4352 & n4367;
  assign n4369 = n4368 ^ n4342;
  assign n4370 = n4369 ^ n4342;
  assign n4371 = n4342 ^ n4341;
  assign n4372 = n4371 ^ n4342;
  assign n4373 = ~n4370 & ~n4372;
  assign n4374 = n4373 ^ n4342;
  assign n4375 = n4348 & ~n4374;
  assign n4376 = n4375 ^ x144;
  assign n4377 = ~n4347 & ~n4376;
  assign n4378 = ~x141 & ~n4233;
  assign n4379 = ~x143 & ~n4242;
  assign n4380 = ~x142 & ~n4235;
  assign n4381 = ~n4379 & ~n4380;
  assign n4382 = ~n4231 & n4381;
  assign n4383 = ~n4378 & n4382;
  assign n4384 = ~x136 & ~n4219;
  assign n4385 = ~n4260 & ~n4384;
  assign n4386 = n4383 & n4385;
  assign n4387 = n4229 & n4386;
  assign n4388 = ~x133 & n4217;
  assign n4389 = n4387 & ~n4388;
  assign n4390 = n4271 & n4389;
  assign n4425 = ~x132 & n4409;
  assign n4426 = n4390 & ~n4425;
  assign n4427 = ~n4377 & n4426;
  assign n4428 = ~n4424 & ~n4427;
  assign n4445 = n4444 ^ n4428;
  assign n5890 = n3987 ^ n3416;
  assign n5891 = n4445 & n5890;
  assign n5892 = n5891 ^ n3416;
  assign n4757 = n4340 ^ x145;
  assign n4729 = n4323 & n4339;
  assign n4730 = ~n4365 & ~n4729;
  assign n4755 = n4328 & ~n4730;
  assign n4756 = n4352 & ~n4755;
  assign n4758 = n4757 ^ n4756;
  assign n4752 = n3681 ^ n3330;
  assign n4753 = ~n3673 & n4752;
  assign n4754 = n4753 ^ n3330;
  assign n4796 = n4758 ^ n4754;
  assign n4735 = n3688 ^ n3331;
  assign n4736 = ~n3679 & ~n4735;
  assign n4737 = n4736 ^ n3331;
  assign n4728 = n4326 ^ x147;
  assign n4731 = n4730 ^ n4326;
  assign n4732 = n4728 & n4731;
  assign n4733 = n4732 ^ x147;
  assign n4734 = n4733 ^ n4350;
  assign n4797 = n4737 ^ n4734;
  assign n4744 = n3700 ^ n3276;
  assign n4745 = ~n3686 & ~n4744;
  assign n4746 = n4745 ^ n3276;
  assign n4643 = n4323 & n4337;
  assign n4644 = n4359 & ~n4643;
  assign n4747 = n4644 ^ n4329;
  assign n4748 = ~n4355 & ~n4747;
  assign n4749 = n4748 ^ x149;
  assign n4750 = n4749 ^ n4354;
  assign n4798 = n4746 & ~n4750;
  assign n4740 = n3694 ^ n3287;
  assign n4741 = n4083 & ~n4740;
  assign n4742 = n4741 ^ n3287;
  assign n4739 = n4730 ^ n4728;
  assign n4799 = n4742 ^ n4739;
  assign n4800 = ~n4798 & n4799;
  assign n4743 = n4739 & n4742;
  assign n4801 = n4800 ^ n4743;
  assign n4802 = n4801 ^ n4734;
  assign n4803 = ~n4797 & ~n4802;
  assign n4804 = n4803 ^ n4737;
  assign n4805 = n4804 ^ n4754;
  assign n4806 = ~n4796 & n4805;
  assign n4807 = n4806 ^ n4758;
  assign n4645 = n4644 ^ n4355;
  assign n4640 = n3712 ^ n3263;
  assign n4641 = n3692 & n4640;
  assign n4642 = n4641 ^ n3263;
  assign n4646 = n4645 ^ n4642;
  assign n4647 = n3723 ^ n3150;
  assign n4648 = n3698 & n4647;
  assign n4649 = n4648 ^ n3150;
  assign n4589 = n4335 ^ x151;
  assign n4590 = n4335 ^ n4323;
  assign n4591 = n4589 & ~n4590;
  assign n4592 = n4591 ^ x151;
  assign n4593 = n4592 ^ n4357;
  assign n4650 = n4649 ^ n4593;
  assign n4651 = n3728 ^ n3144;
  assign n4652 = ~n3708 & ~n4651;
  assign n4653 = n4652 ^ n3144;
  assign n4599 = n4589 ^ n4323;
  assign n4654 = n4653 ^ n4599;
  assign n4655 = n3667 ^ n3139;
  assign n4656 = n3711 & n4655;
  assign n4657 = n4656 ^ n3139;
  assign n4604 = n4320 ^ n4289;
  assign n4658 = n4657 ^ n4604;
  assign n4659 = n3557 ^ n3130;
  assign n4660 = ~n3722 & n4659;
  assign n4661 = n4660 ^ n3130;
  assign n4612 = n4317 ^ n4291;
  assign n4662 = n4661 ^ n4612;
  assign n4663 = n3546 ^ n3124;
  assign n4664 = ~n3732 & n4663;
  assign n4665 = n4664 ^ n3124;
  assign n4618 = n4314 ^ n4293;
  assign n4666 = n4665 ^ n4618;
  assign n4668 = n3299 ^ n3105;
  assign n4669 = n3750 & ~n4668;
  assign n4670 = n4669 ^ n3105;
  assign n4667 = n4305 ^ n4299;
  assign n4671 = n4670 ^ n4667;
  assign n4673 = n3301 ^ n3095;
  assign n4674 = n4041 & ~n4673;
  assign n4675 = n4674 ^ n3095;
  assign n4672 = n4302 ^ n4301;
  assign n4676 = n4675 ^ n4672;
  assign n4680 = n4168 ^ x159;
  assign n4677 = n3304 ^ n3047;
  assign n4678 = n3758 & n4677;
  assign n4679 = n4678 ^ n3047;
  assign n4681 = n4680 ^ n4679;
  assign n4502 = n3936 ^ x103;
  assign n4503 = n3936 ^ n3935;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = n4504 ^ x103;
  assign n4506 = n4505 ^ n3943;
  assign n4471 = n3028 ^ n2711;
  assign n4472 = ~n3420 & ~n4471;
  assign n4473 = n4472 ^ n2711;
  assign n4469 = n3935 ^ x103;
  assign n4470 = n4469 ^ n3936;
  assign n4474 = n4473 ^ n4470;
  assign n4466 = n4438 ^ n4432;
  assign n4467 = n4439 & n4466;
  assign n4468 = n4467 ^ n4432;
  assign n4499 = n4470 ^ n4468;
  assign n4500 = ~n4474 & ~n4499;
  assign n4501 = n4500 ^ n4473;
  assign n4507 = n4506 ^ n4501;
  assign n4496 = n2724 ^ x31;
  assign n4497 = n3416 & n4496;
  assign n4498 = n4497 ^ x31;
  assign n4559 = n4506 ^ n4498;
  assign n4560 = ~n4507 & n4559;
  assign n4561 = n4560 ^ n4498;
  assign n4555 = n3033 ^ n2735;
  assign n4556 = ~n3413 & ~n4555;
  assign n4557 = n4556 ^ n2735;
  assign n4554 = n3946 ^ n3895;
  assign n4558 = n4557 ^ n4554;
  assign n4562 = n4561 ^ n4558;
  assign n4475 = n4474 ^ n4468;
  assign n4476 = n4440 & n4441;
  assign n4509 = ~n4475 & ~n4476;
  assign n4508 = n4507 ^ n4498;
  assign n4510 = n4509 ^ n4508;
  assign n4465 = n4429 & n4442;
  assign n4477 = n4476 ^ n4475;
  assign n4495 = ~n4465 & n4477;
  assign n4551 = n4509 ^ n4495;
  assign n4552 = n4510 & n4551;
  assign n4553 = n4552 ^ n4495;
  assign n4563 = n4562 ^ n4553;
  assign n4564 = n4563 ^ x128;
  assign n4478 = n4477 ^ n4465;
  assign n4479 = n4478 ^ x130;
  assign n4458 = n4443 ^ n4424;
  assign n4459 = ~n4444 & n4458;
  assign n4460 = n4459 ^ x131;
  assign n4513 = n4478 ^ n4460;
  assign n4514 = ~n4479 & n4513;
  assign n4515 = n4514 ^ x130;
  assign n4511 = n4510 ^ n4495;
  assign n4538 = x129 & ~n4511;
  assign n4539 = ~n4515 & ~n4538;
  assign n4461 = ~x131 & n4443;
  assign n4462 = n4426 & ~n4461;
  assign n4516 = ~x130 & n4478;
  assign n4517 = n4462 & ~n4516;
  assign n4540 = n4517 ^ n4377;
  assign n4541 = ~x129 & n4511;
  assign n4542 = n4541 ^ n4517;
  assign n4543 = n4517 & ~n4542;
  assign n4544 = n4543 ^ n4517;
  assign n4545 = ~n4540 & n4544;
  assign n4546 = n4545 ^ n4543;
  assign n4547 = n4546 ^ n4517;
  assign n4548 = n4547 ^ n4541;
  assign n4549 = n4539 & ~n4548;
  assign n4550 = n4549 ^ n4541;
  assign n4565 = n4564 ^ n4550;
  assign n4535 = n3307 ^ n3045;
  assign n4536 = n4030 & ~n4535;
  assign n4537 = n4536 ^ n3045;
  assign n4566 = n4565 ^ n4537;
  assign n4521 = n3311 ^ n3042;
  assign n4522 = n3761 & ~n4521;
  assign n4523 = n4522 ^ n3042;
  assign n4518 = ~n4377 & n4517;
  assign n4519 = ~n4515 & ~n4518;
  assign n4512 = n4511 ^ x129;
  assign n4520 = n4519 ^ n4512;
  assign n4524 = n4523 ^ n4520;
  assign n4481 = n3314 ^ n2719;
  assign n4482 = ~n3770 & n4481;
  assign n4483 = n4482 ^ n2719;
  assign n4463 = ~n4377 & n4462;
  assign n4464 = ~n4460 & ~n4463;
  assign n4480 = n4479 ^ n4464;
  assign n4484 = n4483 ^ n4480;
  assign n4418 = n3317 ^ n3036;
  assign n4419 = ~n3772 & n4418;
  assign n4420 = n4419 ^ n3036;
  assign n4454 = n4445 ^ n4420;
  assign n4391 = ~n4377 & n4390;
  assign n4392 = ~n4284 & ~n4391;
  assign n4411 = n4410 ^ n4392;
  assign n4412 = n3321 ^ n2723;
  assign n4413 = ~n3777 & ~n4412;
  assign n4414 = n4413 ^ n2723;
  assign n4417 = n4411 & n4414;
  assign n4455 = n4445 ^ n4417;
  assign n4456 = ~n4454 & n4455;
  assign n4457 = n4456 ^ n4417;
  assign n4492 = n4483 ^ n4457;
  assign n4493 = ~n4484 & n4492;
  assign n4494 = n4493 ^ n4457;
  assign n4532 = n4520 ^ n4494;
  assign n4533 = n4524 & ~n4532;
  assign n4534 = n4533 ^ n4523;
  assign n4682 = n4537 ^ n4534;
  assign n4683 = ~n4566 & n4682;
  assign n4684 = n4683 ^ n4565;
  assign n4685 = n4684 ^ n4680;
  assign n4686 = ~n4681 & ~n4685;
  assign n4687 = n4686 ^ n4679;
  assign n4688 = n4687 ^ n4672;
  assign n4689 = n4676 & ~n4688;
  assign n4690 = n4689 ^ n4675;
  assign n4691 = n4690 ^ n4667;
  assign n4692 = ~n4671 & n4691;
  assign n4693 = n4692 ^ n4670;
  assign n4694 = n4308 ^ n4297;
  assign n4695 = n3472 ^ n3111;
  assign n4696 = n3742 & ~n4695;
  assign n4697 = n4696 ^ n3111;
  assign n4698 = ~n4694 & n4697;
  assign n4623 = n4311 ^ n4295;
  assign n4699 = n3506 ^ n3116;
  assign n4700 = n3737 & n4699;
  assign n4701 = n4700 ^ n3116;
  assign n4702 = n4623 & n4701;
  assign n4703 = ~n4698 & ~n4702;
  assign n4704 = ~n4693 & n4703;
  assign n4705 = n4701 ^ n4623;
  assign n4706 = n4694 & ~n4697;
  assign n4707 = n4705 & ~n4706;
  assign n4708 = n4707 ^ n4702;
  assign n4709 = ~n4704 & n4708;
  assign n4710 = n4709 ^ n4618;
  assign n4711 = n4666 & n4710;
  assign n4712 = n4711 ^ n4665;
  assign n4713 = n4712 ^ n4612;
  assign n4714 = n4662 & ~n4713;
  assign n4715 = n4714 ^ n4661;
  assign n4716 = n4715 ^ n4604;
  assign n4717 = n4658 & n4716;
  assign n4718 = n4717 ^ n4657;
  assign n4719 = n4718 ^ n4599;
  assign n4720 = n4654 & n4719;
  assign n4721 = n4720 ^ n4653;
  assign n4722 = n4721 ^ n4593;
  assign n4723 = ~n4650 & ~n4722;
  assign n4724 = n4723 ^ n4649;
  assign n4725 = n4724 ^ n4645;
  assign n4726 = n4646 & n4725;
  assign n4727 = n4726 ^ n4642;
  assign n4738 = n4734 & ~n4737;
  assign n4751 = ~n4746 & n4750;
  assign n4759 = n4754 & ~n4758;
  assign n4760 = ~n4751 & ~n4759;
  assign n4761 = ~n4743 & n4760;
  assign n4762 = ~n4738 & n4761;
  assign n4966 = n4727 & n4762;
  assign n4967 = ~n4807 & ~n4966;
  assign n4767 = n3823 ^ n3338;
  assign n4768 = n4100 & n4767;
  assign n4769 = n4768 ^ n3338;
  assign n4763 = n4756 ^ n4340;
  assign n4764 = ~n4757 & ~n4763;
  assign n4765 = n4764 ^ x145;
  assign n4766 = n4765 ^ n4348;
  assign n4965 = n4769 ^ n4766;
  assign n4968 = n4967 ^ n4965;
  assign n5110 = n4968 ^ n2973;
  assign n4946 = n4727 & ~n4751;
  assign n4947 = ~n4743 & n4946;
  assign n4948 = n4801 & ~n4947;
  assign n4957 = n4948 ^ n4734;
  assign n4958 = ~n4797 & ~n4957;
  assign n4959 = n4958 ^ n4737;
  assign n4960 = n4959 ^ n4796;
  assign n4988 = n4960 ^ n2963;
  assign n4949 = n4948 ^ n4797;
  assign n4989 = n4949 ^ n2951;
  assign n4951 = ~n4798 & ~n4946;
  assign n4952 = n4951 ^ n4799;
  assign n4990 = n4952 ^ n2939;
  assign n4954 = n4750 ^ n4746;
  assign n4955 = n4954 ^ n4727;
  assign n4991 = ~n2930 & ~n4955;
  assign n4992 = n4991 ^ n4952;
  assign n4993 = n4990 & n4992;
  assign n4994 = n4993 ^ n2939;
  assign n4995 = n4994 ^ n4949;
  assign n4996 = ~n4989 & n4995;
  assign n4997 = n4996 ^ n2951;
  assign n4998 = n4997 ^ n4960;
  assign n4999 = ~n4988 & ~n4998;
  assign n5000 = n4999 ^ n2963;
  assign n4882 = n4724 ^ n4646;
  assign n4883 = n4882 ^ n2919;
  assign n4884 = n4721 ^ n4650;
  assign n4885 = n4884 ^ n2758;
  assign n4886 = n4718 ^ n4654;
  assign n4887 = n4886 ^ n2727;
  assign n4888 = n4715 ^ n4658;
  assign n4889 = n4888 ^ n2755;
  assign n4890 = n4712 ^ n4662;
  assign n4891 = n4890 ^ n2728;
  assign n4892 = n4709 ^ n4666;
  assign n4893 = n4892 ^ n2729;
  assign n4894 = n4690 ^ n4671;
  assign n4895 = n4894 ^ n2720;
  assign n4896 = n4687 ^ n4676;
  assign n4897 = n4896 ^ n2748;
  assign n4898 = n4684 ^ n4681;
  assign n4899 = n4898 ^ n2746;
  assign n4567 = n4566 ^ n4534;
  assign n4568 = n4567 ^ n2744;
  assign n4525 = n4524 ^ n4494;
  assign n4526 = n4525 ^ n2725;
  assign n4485 = n4484 ^ n4457;
  assign n4486 = n4485 ^ n2732;
  assign n4415 = n4414 ^ n4411;
  assign n4447 = ~n2734 & n4415;
  assign n4448 = n4447 ^ n2733;
  assign n4421 = n4420 ^ n4417;
  assign n4446 = n4445 ^ n4421;
  assign n4451 = n4447 ^ n4446;
  assign n4452 = n4448 & ~n4451;
  assign n4453 = n4452 ^ n2733;
  assign n4489 = n4485 ^ n4453;
  assign n4490 = ~n4486 & ~n4489;
  assign n4491 = n4490 ^ n2732;
  assign n4529 = n4525 ^ n4491;
  assign n4530 = n4526 & n4529;
  assign n4531 = n4530 ^ n2725;
  assign n4900 = n4567 ^ n4531;
  assign n4901 = n4568 & n4900;
  assign n4902 = n4901 ^ n2744;
  assign n4903 = n4902 ^ n4898;
  assign n4904 = n4899 & ~n4903;
  assign n4905 = n4904 ^ n2746;
  assign n4906 = n4905 ^ n4896;
  assign n4907 = n4897 & ~n4906;
  assign n4908 = n4907 ^ n2748;
  assign n4909 = n4908 ^ n4894;
  assign n4910 = n4895 & n4909;
  assign n4911 = n4910 ^ n2720;
  assign n4912 = n4697 ^ n4694;
  assign n4913 = n4912 ^ n4693;
  assign n4914 = ~n2731 & ~n4913;
  assign n4915 = n4694 ^ n4693;
  assign n4916 = ~n4912 & n4915;
  assign n4917 = n4916 ^ n4697;
  assign n4918 = n4917 ^ n4705;
  assign n4919 = n2730 & n4918;
  assign n4920 = ~n4914 & ~n4919;
  assign n4921 = n4911 & n4920;
  assign n4922 = n4918 ^ n2730;
  assign n4923 = n2731 & n4913;
  assign n4924 = n4923 ^ n4918;
  assign n4925 = n4922 & n4924;
  assign n4926 = n4925 ^ n2730;
  assign n4927 = ~n4921 & n4926;
  assign n4928 = n4927 ^ n4892;
  assign n4929 = ~n4893 & ~n4928;
  assign n4930 = n4929 ^ n2729;
  assign n4931 = n4930 ^ n4890;
  assign n4932 = ~n4891 & ~n4931;
  assign n4933 = n4932 ^ n2728;
  assign n4934 = n4933 ^ n4888;
  assign n4935 = n4889 & n4934;
  assign n4936 = n4935 ^ n2755;
  assign n4937 = n4936 ^ n4886;
  assign n4938 = n4887 & n4937;
  assign n4939 = n4938 ^ n2727;
  assign n4940 = n4939 ^ n4884;
  assign n4941 = n4885 & ~n4940;
  assign n4942 = n4941 ^ n2758;
  assign n4943 = n4942 ^ n4882;
  assign n4944 = ~n4883 & ~n4943;
  assign n4945 = n4944 ^ n2919;
  assign n4950 = n2951 & ~n4949;
  assign n4953 = n2939 & n4952;
  assign n4956 = n2930 & n4955;
  assign n4961 = ~n2963 & n4960;
  assign n4962 = ~n4956 & ~n4961;
  assign n4963 = ~n4953 & n4962;
  assign n4964 = ~n4950 & n4963;
  assign n5104 = n4945 & n4964;
  assign n5105 = ~n5000 & ~n5104;
  assign n5111 = n5110 ^ n5105;
  assign n5005 = ~n2973 & n4968;
  assign n4969 = n2973 & ~n4968;
  assign n5106 = ~n4969 & ~n5105;
  assign n5112 = ~n5005 & ~n5106;
  assign n4811 = n4766 & ~n4769;
  assign n4770 = ~n4766 & n4769;
  assign n4970 = ~n4770 & ~n4967;
  assign n4971 = ~n4811 & ~n4970;
  assign n4774 = ~n4243 & ~n4379;
  assign n4775 = n4774 ^ n4377;
  assign n4771 = n3675 ^ n3355;
  assign n4772 = n4115 & n4771;
  assign n4773 = n4772 ^ n3355;
  assign n4812 = n4775 ^ n4773;
  assign n4972 = n4971 ^ n4812;
  assign n5004 = n4972 ^ n2984;
  assign n5113 = n5112 ^ n5004;
  assign n5114 = n5111 & n5113;
  assign n5115 = n4945 & ~n4956;
  assign n5116 = ~n4953 & n5115;
  assign n5117 = n4994 & ~n5116;
  assign n5118 = n5117 ^ n4949;
  assign n5119 = ~n4989 & n5118;
  assign n5120 = n5119 ^ n2951;
  assign n5121 = n5120 ^ n4988;
  assign n5124 = n5117 ^ n4989;
  assign n5140 = ~n4991 & ~n5115;
  assign n5141 = n5140 ^ n4990;
  assign n5142 = n5124 & ~n5141;
  assign n5143 = n5121 & n5142;
  assign n5144 = n5114 & n5143;
  assign n5071 = n4905 ^ n4897;
  assign n4569 = n4568 ^ n4531;
  assign n5072 = n4902 ^ n4899;
  assign n5073 = n4569 & ~n5072;
  assign n5074 = ~n5071 & n5073;
  assign n4416 = n4415 ^ n2734;
  assign n4449 = n4448 ^ n4446;
  assign n4450 = ~n4416 & n4449;
  assign n4487 = n4486 ^ n4453;
  assign n4488 = n4450 & ~n4487;
  assign n4527 = n4526 ^ n4491;
  assign n4528 = ~n4488 & n4527;
  assign n5075 = ~n4528 & ~n5072;
  assign n5076 = ~n5071 & n5075;
  assign n5077 = n4908 ^ n4895;
  assign n5078 = ~n5076 & n5077;
  assign n5079 = ~n5074 & n5078;
  assign n5080 = n4911 ^ n2731;
  assign n5081 = n4913 ^ n4911;
  assign n5082 = n5080 & ~n5081;
  assign n5083 = n5082 ^ n2731;
  assign n5084 = n5083 ^ n4922;
  assign n5085 = n4927 ^ n4893;
  assign n5086 = n5084 & n5085;
  assign n5087 = n4942 ^ n4883;
  assign n5088 = n5086 & n5087;
  assign n5089 = ~n5079 & n5088;
  assign n5090 = n4913 ^ n2731;
  assign n5091 = n5090 ^ n4911;
  assign n5092 = n5086 & n5091;
  assign n5093 = n4930 ^ n4891;
  assign n5094 = ~n5092 & n5093;
  assign n5095 = n4933 ^ n4889;
  assign n5096 = n4936 ^ n4887;
  assign n5097 = n5095 & ~n5096;
  assign n5098 = n4939 ^ n4885;
  assign n5099 = n5097 & n5098;
  assign n5100 = n5087 & n5099;
  assign n5101 = n5094 & n5100;
  assign n5102 = n5101 ^ n5087;
  assign n5103 = ~n5089 & ~n5102;
  assign n5122 = n4955 ^ n2930;
  assign n5123 = n5122 ^ n4945;
  assign n5125 = n5123 & n5124;
  assign n5126 = n5121 & n5125;
  assign n5127 = n5114 & n5126;
  assign n5188 = ~n5103 & n5127;
  assign n5189 = ~n5144 & ~n5188;
  assign n5006 = n5005 ^ n4972;
  assign n5007 = ~n5004 & ~n5006;
  assign n5008 = n5007 ^ n2984;
  assign n4973 = n2984 & ~n4972;
  assign n5107 = ~n4973 & n5106;
  assign n5108 = n5008 & ~n5107;
  assign n4813 = ~n4811 & ~n4812;
  assign n4776 = ~n4773 & n4775;
  assign n4814 = n4813 ^ n4776;
  assign n4974 = ~n4776 & n4970;
  assign n4975 = n4814 & ~n4974;
  assign n4780 = n3383 ^ n3293;
  assign n4781 = n4404 & ~n4780;
  assign n4782 = n4781 ^ n3383;
  assign n4777 = ~n4377 & n4774;
  assign n4778 = n4777 ^ n4243;
  assign n4779 = n4778 ^ n4236;
  assign n4810 = n4782 ^ n4779;
  assign n4976 = n4975 ^ n4810;
  assign n5003 = n4976 ^ n2995;
  assign n5109 = n5108 ^ n5003;
  assign n5190 = n5189 ^ n5109;
  assign n5191 = n5190 ^ x169;
  assign n5192 = ~n5103 & n5126;
  assign n5193 = ~n5143 & n5192;
  assign n5194 = n5193 ^ n5103;
  assign n5195 = n5194 ^ n5103;
  assign n5196 = n5195 ^ n5143;
  assign n5197 = n5111 & ~n5196;
  assign n5198 = n5197 ^ n5111;
  assign n5199 = n5198 ^ n5113;
  assign n5200 = n5199 ^ x170;
  assign n5201 = n5143 ^ n5111;
  assign n5202 = n5201 ^ n5193;
  assign n5203 = n5202 ^ x171;
  assign n5204 = ~n5103 & n5125;
  assign n5205 = ~n5142 & ~n5204;
  assign n5206 = n5205 ^ n5121;
  assign n5207 = n5206 ^ x172;
  assign n5208 = ~n5103 & n5123;
  assign n5209 = n5141 & ~n5208;
  assign n5210 = n5209 ^ n5124;
  assign n5211 = n5210 ^ x173;
  assign n5212 = n5208 ^ n5141;
  assign n5213 = n5212 ^ x174;
  assign n5214 = n5123 ^ n5103;
  assign n5215 = n5214 ^ x175;
  assign n5216 = ~n5079 & n5086;
  assign n5217 = n5094 & ~n5216;
  assign n5218 = n5099 & n5217;
  assign n5219 = n5218 ^ n5087;
  assign n5220 = n5219 ^ x176;
  assign n5221 = n5097 & n5217;
  assign n5222 = n5221 ^ n5098;
  assign n5223 = n5222 ^ x177;
  assign n5224 = ~n5074 & ~n5076;
  assign n5225 = n5224 ^ n5077;
  assign n5226 = n5225 ^ x184;
  assign n4572 = n4527 ^ n4488;
  assign n4573 = n4572 ^ x188;
  assign n4574 = x191 & n4416;
  assign n4575 = n4574 ^ x190;
  assign n4576 = n4449 ^ n4416;
  assign n4577 = n4576 ^ n4574;
  assign n4578 = n4575 & n4577;
  assign n4579 = n4578 ^ x190;
  assign n4580 = n4579 ^ x189;
  assign n4581 = n4487 ^ n4450;
  assign n4582 = n4581 ^ n4579;
  assign n4583 = n4580 & n4582;
  assign n4584 = n4583 ^ x189;
  assign n4585 = n4584 ^ n4572;
  assign n4586 = n4573 & ~n4585;
  assign n4587 = n4586 ^ x188;
  assign n4570 = n4569 ^ n4528;
  assign n5227 = ~x187 & ~n4570;
  assign n5228 = n4528 & ~n4569;
  assign n5229 = n5228 ^ n5072;
  assign n5230 = ~x186 & ~n5229;
  assign n5231 = ~n5227 & ~n5230;
  assign n5232 = n4587 & n5231;
  assign n5233 = n5229 ^ x186;
  assign n5234 = x187 & n4570;
  assign n5235 = n5234 ^ n5229;
  assign n5236 = n5233 & ~n5235;
  assign n5237 = n5236 ^ x186;
  assign n5238 = ~n5232 & ~n5237;
  assign n5239 = n5238 ^ x185;
  assign n5240 = ~n5072 & n5228;
  assign n5241 = n5240 ^ n5072;
  assign n5242 = n5241 ^ n5071;
  assign n5243 = n5242 ^ n5238;
  assign n5244 = ~n5239 & n5243;
  assign n5245 = n5244 ^ x185;
  assign n5246 = n5245 ^ n5225;
  assign n5247 = ~n5226 & n5246;
  assign n5248 = n5247 ^ x184;
  assign n5249 = n5079 & ~n5091;
  assign n5250 = n5249 ^ n5084;
  assign n5251 = ~x182 & n5250;
  assign n5252 = n5091 ^ n5079;
  assign n5253 = ~x183 & ~n5252;
  assign n5254 = ~n5251 & ~n5253;
  assign n5255 = n5084 & n5249;
  assign n5256 = n5255 ^ n5084;
  assign n5257 = n5256 ^ n5085;
  assign n5258 = ~x181 & ~n5257;
  assign n5259 = n5254 & ~n5258;
  assign n5260 = ~n5092 & ~n5216;
  assign n5261 = n5260 ^ n5093;
  assign n5262 = ~x180 & n5261;
  assign n5263 = n5259 & ~n5262;
  assign n5264 = n5248 & n5263;
  assign n5265 = n5261 ^ x180;
  assign n5266 = n5257 ^ x181;
  assign n5267 = x183 & n5252;
  assign n5268 = n5267 ^ x182;
  assign n5269 = n5267 ^ n5250;
  assign n5270 = n5268 & n5269;
  assign n5271 = n5270 ^ x182;
  assign n5272 = n5271 ^ n5257;
  assign n5273 = n5266 & ~n5272;
  assign n5274 = n5273 ^ x181;
  assign n5275 = n5274 ^ n5261;
  assign n5276 = ~n5265 & n5275;
  assign n5277 = n5276 ^ x180;
  assign n5278 = ~n5264 & ~n5277;
  assign n5279 = n5217 ^ n5095;
  assign n5280 = ~x179 & n5279;
  assign n5281 = n5095 & n5217;
  assign n5282 = n5281 ^ n5096;
  assign n5283 = ~x178 & ~n5282;
  assign n5284 = ~n5280 & ~n5283;
  assign n5285 = ~n5278 & n5284;
  assign n5286 = n5282 ^ x178;
  assign n5287 = x179 & ~n5279;
  assign n5288 = n5287 ^ n5282;
  assign n5289 = n5286 & ~n5288;
  assign n5290 = n5289 ^ x178;
  assign n5291 = ~n5285 & ~n5290;
  assign n5292 = n5291 ^ n5222;
  assign n5293 = ~n5223 & ~n5292;
  assign n5294 = n5293 ^ x177;
  assign n5295 = n5294 ^ n5219;
  assign n5296 = ~n5220 & n5295;
  assign n5297 = n5296 ^ x176;
  assign n5298 = n5297 ^ n5214;
  assign n5299 = ~n5215 & n5298;
  assign n5300 = n5299 ^ x175;
  assign n5301 = n5300 ^ n5212;
  assign n5302 = n5213 & ~n5301;
  assign n5303 = n5302 ^ x174;
  assign n5304 = n5303 ^ n5210;
  assign n5305 = ~n5211 & n5304;
  assign n5306 = n5305 ^ x173;
  assign n5307 = n5306 ^ n5206;
  assign n5308 = ~n5207 & n5307;
  assign n5309 = n5308 ^ x172;
  assign n5310 = n5309 ^ n5202;
  assign n5311 = n5203 & ~n5310;
  assign n5312 = n5311 ^ x171;
  assign n5313 = n5312 ^ n5199;
  assign n5314 = n5200 & ~n5313;
  assign n5315 = n5314 ^ x170;
  assign n5316 = n5315 ^ n5190;
  assign n5317 = ~n5191 & n5316;
  assign n5318 = n5317 ^ x169;
  assign n5885 = n5318 ^ x168;
  assign n5145 = n5109 & n5144;
  assign n5128 = n5109 & n5127;
  assign n5169 = ~n5103 & n5128;
  assign n5185 = ~n5145 & ~n5169;
  assign n5146 = n5108 ^ n4976;
  assign n5147 = ~n5003 & ~n5146;
  assign n5148 = n5147 ^ n2995;
  assign n4978 = n4975 ^ n4782;
  assign n4979 = n4810 & n4978;
  assign n4980 = n4979 ^ n4779;
  assign n4787 = n3862 ^ n3396;
  assign n4788 = n4438 & ~n4787;
  assign n4789 = n4788 ^ n3396;
  assign n4784 = ~n4377 & n4381;
  assign n4785 = ~n4246 & ~n4784;
  assign n4786 = n4785 ^ n4234;
  assign n4809 = n4789 ^ n4786;
  assign n4981 = n4980 ^ n4809;
  assign n5002 = n4981 ^ n3007;
  assign n5149 = n5148 ^ n5002;
  assign n5186 = n5185 ^ n5149;
  assign n5886 = n5885 ^ n5186;
  assign n5997 = n5892 ^ n5886;
  assign n5825 = n4007 ^ n3420;
  assign n5826 = n4411 & n5825;
  assign n5827 = n5826 ^ n3420;
  assign n5823 = n5315 ^ x169;
  assign n5824 = n5823 ^ n5190;
  assign n5828 = n5827 ^ n5824;
  assign n4873 = ~n4377 & n4387;
  assign n4874 = ~n4266 & ~n4873;
  assign n5362 = n4271 & ~n4874;
  assign n5363 = n4278 & ~n5362;
  assign n5364 = n5363 ^ n4218;
  assign n5745 = n3990 ^ n3428;
  assign n5746 = n5364 & n5745;
  assign n5747 = n5746 ^ n3428;
  assign n5744 = n5312 ^ n5200;
  assign n5748 = n5747 ^ n5744;
  assign n4875 = n4269 ^ x135;
  assign n5063 = n4874 ^ n4269;
  assign n5064 = ~n4875 & ~n5063;
  assign n5065 = n5064 ^ x135;
  assign n5066 = n5065 ^ n4276;
  assign n5751 = n3998 ^ n3423;
  assign n5752 = n5066 & n5751;
  assign n5753 = n5752 ^ n3423;
  assign n5749 = n5309 ^ x171;
  assign n5750 = n5749 ^ n5202;
  assign n5754 = n5753 ^ n5750;
  assign n5795 = n5300 ^ n5213;
  assign n5787 = n5297 ^ n5215;
  assign n5779 = n5294 ^ n5220;
  assign n5771 = n5291 ^ n5223;
  assign n5759 = n5279 ^ x179;
  assign n5760 = n5279 ^ n5278;
  assign n5761 = ~n5759 & ~n5760;
  assign n5762 = n5761 ^ x179;
  assign n5763 = n5762 ^ n5286;
  assign n5703 = n5278 ^ x179;
  assign n5704 = n5703 ^ n5279;
  assign n5700 = n3694 ^ n3673;
  assign n5701 = n4779 & ~n5700;
  assign n5702 = n5701 ^ n3694;
  assign n5705 = n5704 ^ n5702;
  assign n5585 = n5248 & n5254;
  assign n5586 = ~n5271 & ~n5585;
  assign n5679 = n5586 ^ n5257;
  assign n5680 = n5266 & n5679;
  assign n5681 = n5680 ^ x181;
  assign n5682 = n5681 ^ n5265;
  assign n5587 = n5586 ^ n5266;
  assign n5550 = n5252 ^ x183;
  assign n5567 = n5248 & n5550;
  assign n5568 = n5567 ^ n5267;
  assign n5566 = n5250 ^ x182;
  assign n5569 = n5568 ^ n5566;
  assign n5551 = n5550 ^ n5248;
  assign n5547 = n3728 ^ n3692;
  assign n5548 = ~n4734 & ~n5547;
  assign n5549 = n5548 ^ n3728;
  assign n5552 = n5551 ^ n5549;
  assign n5534 = n5245 ^ n5226;
  assign n5531 = n3698 ^ n3667;
  assign n5532 = ~n4739 & ~n5531;
  assign n5533 = n5532 ^ n3667;
  assign n5535 = n5534 ^ n5533;
  assign n5493 = n5242 ^ x185;
  assign n5494 = n5493 ^ n5238;
  assign n5490 = n3708 ^ n3557;
  assign n5491 = ~n4750 & ~n5490;
  assign n5492 = n5491 ^ n3557;
  assign n5495 = n5494 ^ n5492;
  assign n4571 = n4570 ^ x187;
  assign n5429 = n4571 & n4587;
  assign n5430 = n5429 ^ n5234;
  assign n5431 = n5430 ^ n5233;
  assign n5426 = n3711 ^ n3546;
  assign n5427 = n4645 & n5426;
  assign n5428 = n5427 ^ n3546;
  assign n5432 = n5431 ^ n5428;
  assign n4594 = n3722 ^ n3506;
  assign n4595 = n4593 & n4594;
  assign n4596 = n4595 ^ n3506;
  assign n4588 = n4587 ^ n4571;
  assign n4597 = n4596 ^ n4588;
  assign n4600 = n3732 ^ n3472;
  assign n4601 = n4599 & ~n4600;
  assign n4602 = n4601 ^ n3472;
  assign n4598 = n4584 ^ n4573;
  assign n4603 = n4602 ^ n4598;
  assign n4608 = n4581 ^ x189;
  assign n4609 = n4608 ^ n4579;
  assign n4605 = n3737 ^ n3299;
  assign n4606 = ~n4604 & n4605;
  assign n4607 = n4606 ^ n3299;
  assign n4610 = n4609 ^ n4607;
  assign n4613 = n3742 ^ n3301;
  assign n4614 = n4612 & n4613;
  assign n4615 = n4614 ^ n3301;
  assign n4611 = n4576 ^ n4575;
  assign n4616 = n4615 ^ n4611;
  assign n4619 = n3750 ^ n3304;
  assign n4620 = n4618 & ~n4619;
  assign n4621 = n4620 ^ n3304;
  assign n4617 = n4416 ^ x191;
  assign n4622 = n4621 ^ n4617;
  assign n5060 = n3327 ^ n2724;
  assign n5061 = n3987 & ~n5060;
  assign n5062 = n5061 ^ n2724;
  assign n5067 = n5066 ^ n5062;
  assign n4876 = n4875 ^ n4874;
  assign n4870 = n3413 ^ n3028;
  assign n4871 = ~n4007 & ~n4870;
  assign n4872 = n4871 ^ n3028;
  assign n4877 = n4876 ^ n4872;
  assign n4630 = n4254 ^ x137;
  assign n4631 = ~n4377 & n4383;
  assign n4632 = ~n4252 & ~n4631;
  assign n4633 = n4229 & ~n4632;
  assign n4634 = n4227 & ~n4633;
  assign n4635 = n4634 ^ n4254;
  assign n4636 = n4630 & n4635;
  assign n4637 = n4636 ^ x137;
  assign n4638 = n4637 ^ n4220;
  assign n4627 = n3416 ^ n3012;
  assign n4628 = n3990 & ~n4627;
  assign n4629 = n4628 ^ n3012;
  assign n4639 = n4638 ^ n4629;
  assign n4783 = ~n4779 & ~n4782;
  assign n4790 = n4786 & ~n4789;
  assign n4791 = ~n4783 & ~n4790;
  assign n4792 = ~n4776 & n4791;
  assign n4793 = ~n4770 & n4792;
  assign n4794 = n4762 & n4793;
  assign n4795 = n4727 & n4794;
  assign n4808 = n4793 & n4807;
  assign n4815 = n4814 ^ n4779;
  assign n4816 = n4810 & n4815;
  assign n4817 = n4816 ^ n4782;
  assign n4818 = n4817 ^ n4786;
  assign n4819 = ~n4809 & ~n4818;
  assign n4820 = n4819 ^ n4786;
  assign n4821 = ~n4808 & n4820;
  assign n4822 = ~n4795 & n4821;
  assign n4823 = n3428 ^ n3013;
  assign n4824 = n4554 & n4823;
  assign n4825 = n4824 ^ n3013;
  assign n4826 = n4221 ^ x139;
  assign n4827 = n4632 ^ n4221;
  assign n4828 = n4826 & n4827;
  assign n4829 = n4828 ^ x139;
  assign n4830 = n4829 ^ n4224;
  assign n4831 = ~n4825 & ~n4830;
  assign n4832 = n3973 ^ n3294;
  assign n4833 = n4470 & ~n4832;
  assign n4834 = n4833 ^ n3294;
  assign n4835 = n4785 ^ n4233;
  assign n4836 = n4234 & n4835;
  assign n4837 = n4836 ^ x141;
  assign n4838 = n4837 ^ n4232;
  assign n4839 = ~n4834 & n4838;
  assign n4840 = n4826 ^ n4632;
  assign n4841 = n3423 ^ n3078;
  assign n4842 = ~n4506 & ~n4841;
  assign n4843 = n4842 ^ n3078;
  assign n4844 = n4840 & n4843;
  assign n4845 = n4634 ^ n4630;
  assign n4846 = n3420 ^ n3015;
  assign n4847 = n3998 & ~n4846;
  assign n4848 = n4847 ^ n3015;
  assign n4849 = n4845 & ~n4848;
  assign n4850 = ~n4844 & ~n4849;
  assign n4851 = ~n4839 & n4850;
  assign n4852 = ~n4831 & n4851;
  assign n4853 = ~n4822 & n4852;
  assign n4854 = n4848 ^ n4845;
  assign n4855 = n4830 ^ n4825;
  assign n4856 = n4834 & ~n4838;
  assign n4857 = n4843 ^ n4840;
  assign n4858 = ~n4856 & n4857;
  assign n4859 = n4858 ^ n4844;
  assign n4860 = n4859 ^ n4830;
  assign n4861 = n4855 & n4860;
  assign n4862 = n4861 ^ n4825;
  assign n4863 = n4862 ^ n4845;
  assign n4864 = ~n4854 & n4863;
  assign n4865 = n4864 ^ n4848;
  assign n4866 = ~n4853 & ~n4865;
  assign n4867 = n4866 ^ n4638;
  assign n4868 = ~n4639 & n4867;
  assign n4869 = n4868 ^ n4629;
  assign n5057 = n4872 ^ n4869;
  assign n5058 = n4877 & n5057;
  assign n5059 = n5058 ^ n4876;
  assign n5068 = n5067 ^ n5059;
  assign n5069 = n5068 ^ x31;
  assign n4878 = n4877 ^ n4869;
  assign n4879 = n4878 ^ n2711;
  assign n4880 = n4866 ^ n4639;
  assign n4881 = n4880 ^ n2690;
  assign n4977 = ~n2995 & n4976;
  assign n4982 = ~n3007 & n4981;
  assign n4983 = ~n4977 & ~n4982;
  assign n4984 = ~n4973 & n4983;
  assign n4985 = ~n4969 & n4984;
  assign n4986 = n4964 & n4985;
  assign n4987 = n4945 & n4986;
  assign n5001 = n4985 & n5000;
  assign n5009 = n5008 ^ n4976;
  assign n5010 = ~n5003 & ~n5009;
  assign n5011 = n5010 ^ n2995;
  assign n5012 = n5011 ^ n4981;
  assign n5013 = ~n5002 & ~n5012;
  assign n5014 = n5013 ^ n4981;
  assign n5015 = ~n5001 & n5014;
  assign n5016 = ~n4987 & n5015;
  assign n5017 = ~n4822 & ~n4839;
  assign n5018 = ~n4844 & n5017;
  assign n5019 = n4859 & ~n5018;
  assign n5020 = n5019 ^ n4855;
  assign n5021 = ~n2682 & n5020;
  assign n5022 = ~n4856 & ~n5017;
  assign n5023 = n5022 ^ n4857;
  assign n5024 = ~n2686 & n5023;
  assign n5025 = n4838 ^ n4834;
  assign n5026 = n5025 ^ n4822;
  assign n5027 = ~n3025 & ~n5026;
  assign n5028 = n5019 ^ n4830;
  assign n5029 = n4855 & n5028;
  assign n5030 = n5029 ^ n4825;
  assign n5031 = n5030 ^ n4854;
  assign n5032 = n2684 & n5031;
  assign n5033 = ~n5027 & ~n5032;
  assign n5034 = ~n5024 & n5033;
  assign n5035 = ~n5021 & n5034;
  assign n5036 = ~n5016 & n5035;
  assign n5037 = n5031 ^ n2684;
  assign n5038 = n5020 ^ n2682;
  assign n5039 = n3025 & n5026;
  assign n5040 = n5039 ^ n2686;
  assign n5041 = n5039 ^ n5023;
  assign n5042 = n5040 & n5041;
  assign n5043 = n5042 ^ n2686;
  assign n5044 = n5043 ^ n5020;
  assign n5045 = ~n5038 & n5044;
  assign n5046 = n5045 ^ n2682;
  assign n5047 = n5046 ^ n5031;
  assign n5048 = n5037 & n5047;
  assign n5049 = n5048 ^ n2684;
  assign n5050 = ~n5036 & n5049;
  assign n5051 = n5050 ^ n4880;
  assign n5052 = n4881 & n5051;
  assign n5053 = n5052 ^ n2690;
  assign n5054 = n5053 ^ n4878;
  assign n5055 = n4879 & n5054;
  assign n5056 = n5055 ^ n2711;
  assign n5070 = n5069 ^ n5056;
  assign n5129 = n5026 ^ n3025;
  assign n5130 = n5129 ^ n5016;
  assign n5131 = ~n5016 & ~n5027;
  assign n5132 = ~n5024 & n5131;
  assign n5133 = ~n5043 & ~n5132;
  assign n5134 = n5133 ^ n5038;
  assign n5135 = ~n5130 & n5134;
  assign n5136 = n5053 ^ n4879;
  assign n5137 = n5135 & n5136;
  assign n5138 = n5128 & n5137;
  assign n5139 = ~n5103 & n5138;
  assign n5150 = ~n5145 & n5149;
  assign n5151 = n5135 & ~n5150;
  assign n5152 = n5133 ^ n2682;
  assign n5153 = n5133 ^ n5020;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = n5154 ^ n2682;
  assign n5156 = n5155 ^ n5037;
  assign n5158 = ~n5039 & ~n5131;
  assign n5157 = n5023 ^ n2686;
  assign n5159 = n5158 ^ n5157;
  assign n5160 = n5134 & n5159;
  assign n5161 = ~n5156 & ~n5160;
  assign n5162 = ~n5151 & n5161;
  assign n5163 = n5050 ^ n4881;
  assign n5164 = n5162 & n5163;
  assign n5165 = n5136 & ~n5164;
  assign n5166 = ~n5139 & ~n5165;
  assign n5369 = n5070 & n5166;
  assign n5359 = n3323 ^ n3033;
  assign n5360 = n3977 & n5359;
  assign n5361 = n5360 ^ n3033;
  assign n5365 = n5364 ^ n5361;
  assign n5356 = n5066 ^ n5059;
  assign n5357 = ~n5067 & ~n5356;
  assign n5358 = n5357 ^ n5062;
  assign n5366 = n5365 ^ n5358;
  assign n5367 = n5366 ^ n2735;
  assign n5352 = n5056 ^ x31;
  assign n5353 = n5068 ^ n5056;
  assign n5354 = n5352 & ~n5353;
  assign n5355 = n5354 ^ x31;
  assign n5368 = n5367 ^ n5355;
  assign n5370 = n5369 ^ n5368;
  assign n5167 = n5166 ^ n5070;
  assign n5168 = n5167 ^ x161;
  assign n5170 = n5135 & n5169;
  assign n5171 = ~n5151 & ~n5160;
  assign n5172 = ~n5170 & n5171;
  assign n5173 = n5172 ^ n5156;
  assign n5174 = n5173 ^ x164;
  assign n5175 = n5150 & ~n5169;
  assign n5176 = ~n5130 & n5175;
  assign n5177 = n5176 ^ n5130;
  assign n5178 = ~n5159 & n5177;
  assign n5179 = n5178 ^ n5134;
  assign n5180 = n5179 ^ x165;
  assign n5181 = n5177 ^ n5159;
  assign n5182 = n5181 ^ x166;
  assign n5183 = n5175 ^ n5130;
  assign n5184 = n5183 ^ x167;
  assign n5187 = n5186 ^ x168;
  assign n5319 = n5318 ^ n5186;
  assign n5320 = ~n5187 & n5319;
  assign n5321 = n5320 ^ x168;
  assign n5322 = n5321 ^ n5183;
  assign n5323 = n5184 & ~n5322;
  assign n5324 = n5323 ^ x167;
  assign n5325 = n5324 ^ n5181;
  assign n5326 = n5182 & ~n5325;
  assign n5327 = n5326 ^ x166;
  assign n5328 = n5327 ^ n5179;
  assign n5329 = ~n5180 & n5328;
  assign n5330 = n5329 ^ x165;
  assign n5331 = n5330 ^ n5173;
  assign n5332 = n5174 & ~n5331;
  assign n5333 = n5332 ^ x164;
  assign n5334 = n5162 & ~n5170;
  assign n5335 = n5334 ^ n5163;
  assign n5336 = ~x163 & n5335;
  assign n5337 = n5163 & n5334;
  assign n5338 = n5337 ^ n5136;
  assign n5339 = ~x162 & n5338;
  assign n5340 = ~n5336 & ~n5339;
  assign n5341 = n5333 & n5340;
  assign n5342 = n5338 ^ x162;
  assign n5343 = x163 & ~n5335;
  assign n5344 = n5343 ^ n5338;
  assign n5345 = ~n5342 & n5344;
  assign n5346 = n5345 ^ x162;
  assign n5347 = ~n5341 & ~n5346;
  assign n5348 = n5347 ^ n5167;
  assign n5349 = ~n5168 & ~n5348;
  assign n5350 = n5349 ^ x161;
  assign n5351 = n5350 ^ x160;
  assign n5371 = n5370 ^ n5351;
  assign n4624 = n4041 ^ n3307;
  assign n4625 = ~n4623 & n4624;
  assign n4626 = n4625 ^ n3307;
  assign n5372 = n5371 ^ n4626;
  assign n5375 = n3758 ^ n3311;
  assign n5376 = n4694 & ~n5375;
  assign n5377 = n5376 ^ n3311;
  assign n5373 = n5347 ^ x161;
  assign n5374 = n5373 ^ n5167;
  assign n5378 = n5377 ^ n5374;
  assign n5384 = n4030 ^ n3314;
  assign n5385 = n4667 & n5384;
  assign n5386 = n5385 ^ n3314;
  assign n5379 = n5335 ^ x163;
  assign n5380 = n5335 ^ n5333;
  assign n5381 = ~n5379 & n5380;
  assign n5382 = n5381 ^ x163;
  assign n5383 = n5382 ^ n5342;
  assign n5387 = n5386 ^ n5383;
  assign n5391 = n5379 ^ n5333;
  assign n5388 = n3761 ^ n3317;
  assign n5389 = ~n4672 & n5388;
  assign n5390 = n5389 ^ n3317;
  assign n5392 = n5391 ^ n5390;
  assign n5393 = n5330 ^ x164;
  assign n5394 = n5393 ^ n5173;
  assign n5395 = n3770 ^ n3321;
  assign n5396 = n4680 & n5395;
  assign n5397 = n5396 ^ n3321;
  assign n5398 = n5394 & ~n5397;
  assign n5399 = n5398 ^ n5391;
  assign n5400 = n5392 & ~n5399;
  assign n5401 = n5400 ^ n5398;
  assign n5402 = n5401 ^ n5383;
  assign n5403 = ~n5387 & n5402;
  assign n5404 = n5403 ^ n5386;
  assign n5405 = n5404 ^ n5374;
  assign n5406 = ~n5378 & ~n5405;
  assign n5407 = n5406 ^ n5377;
  assign n5408 = n5407 ^ n5371;
  assign n5409 = n5372 & n5408;
  assign n5410 = n5409 ^ n4626;
  assign n5411 = n5410 ^ n4617;
  assign n5412 = ~n4622 & ~n5411;
  assign n5413 = n5412 ^ n4621;
  assign n5414 = n5413 ^ n4611;
  assign n5415 = ~n4616 & ~n5414;
  assign n5416 = n5415 ^ n4615;
  assign n5417 = n5416 ^ n4609;
  assign n5418 = ~n4610 & n5417;
  assign n5419 = n5418 ^ n4607;
  assign n5420 = n5419 ^ n4598;
  assign n5421 = n4603 & ~n5420;
  assign n5422 = n5421 ^ n4602;
  assign n5423 = n5422 ^ n4588;
  assign n5424 = ~n4597 & ~n5423;
  assign n5425 = n5424 ^ n4596;
  assign n5487 = n5431 ^ n5425;
  assign n5488 = n5432 & n5487;
  assign n5489 = n5488 ^ n5428;
  assign n5528 = n5494 ^ n5489;
  assign n5529 = ~n5495 & n5528;
  assign n5530 = n5529 ^ n5492;
  assign n5544 = n5534 ^ n5530;
  assign n5545 = n5535 & n5544;
  assign n5546 = n5545 ^ n5533;
  assign n5563 = n5551 ^ n5546;
  assign n5564 = ~n5552 & n5563;
  assign n5565 = n5564 ^ n5549;
  assign n5570 = n5569 ^ n5565;
  assign n5560 = n3723 ^ n3686;
  assign n5561 = n4758 & n5560;
  assign n5562 = n5561 ^ n3723;
  assign n5582 = n5569 ^ n5562;
  assign n5583 = ~n5570 & n5582;
  assign n5584 = n5583 ^ n5562;
  assign n5588 = n5587 ^ n5584;
  assign n5579 = n4083 ^ n3712;
  assign n5580 = n4766 & n5579;
  assign n5581 = n5580 ^ n3712;
  assign n5676 = n5587 ^ n5581;
  assign n5677 = ~n5588 & ~n5676;
  assign n5678 = n5677 ^ n5581;
  assign n5683 = n5682 ^ n5678;
  assign n5673 = n3700 ^ n3679;
  assign n5674 = ~n4775 & n5673;
  assign n5675 = n5674 ^ n3700;
  assign n5697 = n5682 ^ n5675;
  assign n5698 = n5683 & n5697;
  assign n5699 = n5698 ^ n5675;
  assign n5756 = n5704 ^ n5699;
  assign n5757 = n5705 & n5756;
  assign n5758 = n5757 ^ n5702;
  assign n5764 = n5763 ^ n5758;
  assign n5765 = n4100 ^ n3688;
  assign n5766 = ~n4786 & ~n5765;
  assign n5767 = n5766 ^ n3688;
  assign n5768 = n5767 ^ n5763;
  assign n5769 = ~n5764 & ~n5768;
  assign n5770 = n5769 ^ n5767;
  assign n5772 = n5771 ^ n5770;
  assign n5773 = n4115 ^ n3681;
  assign n5774 = ~n4838 & ~n5773;
  assign n5775 = n5774 ^ n3681;
  assign n5776 = n5775 ^ n5771;
  assign n5777 = n5772 & ~n5776;
  assign n5778 = n5777 ^ n5775;
  assign n5780 = n5779 ^ n5778;
  assign n5781 = n4404 ^ n3823;
  assign n5782 = ~n4840 & ~n5781;
  assign n5783 = n5782 ^ n3823;
  assign n5784 = n5783 ^ n5779;
  assign n5785 = ~n5780 & n5784;
  assign n5786 = n5785 ^ n5783;
  assign n5788 = n5787 ^ n5786;
  assign n5789 = n4438 ^ n3675;
  assign n5790 = n4830 & n5789;
  assign n5791 = n5790 ^ n3675;
  assign n5792 = n5791 ^ n5787;
  assign n5793 = ~n5788 & ~n5792;
  assign n5794 = n5793 ^ n5791;
  assign n5796 = n5795 ^ n5794;
  assign n5797 = n4470 ^ n3293;
  assign n5798 = ~n4845 & ~n5797;
  assign n5799 = n5798 ^ n3293;
  assign n5800 = n5799 ^ n5795;
  assign n5801 = ~n5796 & ~n5800;
  assign n5802 = n5801 ^ n5799;
  assign n5755 = n5303 ^ n5211;
  assign n5803 = n5802 ^ n5755;
  assign n5804 = n4506 ^ n3862;
  assign n5805 = n4638 & n5804;
  assign n5806 = n5805 ^ n3862;
  assign n5807 = n5806 ^ n5755;
  assign n5808 = ~n5803 & n5807;
  assign n5809 = n5808 ^ n5806;
  assign n5711 = n5306 ^ n5207;
  assign n5810 = n5809 ^ n5711;
  assign n5811 = n4554 ^ n3973;
  assign n5812 = n4876 & ~n5811;
  assign n5813 = n5812 ^ n3973;
  assign n5814 = n5813 ^ n5711;
  assign n5815 = ~n5810 & n5814;
  assign n5816 = n5815 ^ n5813;
  assign n5817 = n5816 ^ n5750;
  assign n5818 = n5754 & n5817;
  assign n5819 = n5818 ^ n5753;
  assign n5820 = n5819 ^ n5744;
  assign n5821 = n5748 & ~n5820;
  assign n5822 = n5821 ^ n5747;
  assign n5887 = n5824 ^ n5822;
  assign n5888 = n5828 & n5887;
  assign n5889 = n5888 ^ n5827;
  assign n5998 = n5889 ^ n5886;
  assign n5999 = ~n5997 & ~n5998;
  assign n6000 = n5999 ^ n5892;
  assign n5996 = n5321 ^ n5184;
  assign n6001 = n6000 ^ n5996;
  assign n5993 = n3977 ^ n3413;
  assign n5994 = n4480 & ~n5993;
  assign n5995 = n5994 ^ n3413;
  assign n6018 = n5996 ^ n5995;
  assign n6019 = ~n6001 & ~n6018;
  assign n6020 = n6019 ^ n5995;
  assign n6016 = n5324 ^ x166;
  assign n6017 = n6016 ^ n5181;
  assign n6021 = n6020 ^ n6017;
  assign n6013 = n3777 ^ n3327;
  assign n6014 = n4520 & ~n6013;
  assign n6015 = n6014 ^ n3327;
  assign n6022 = n6021 ^ n6015;
  assign n6002 = n6001 ^ n5995;
  assign n6009 = n6002 ^ n3028;
  assign n5893 = n5892 ^ n5889;
  assign n5894 = n5893 ^ n5886;
  assign n5895 = n5894 ^ n3012;
  assign n5829 = n5828 ^ n5822;
  assign n5830 = n5829 ^ n3015;
  assign n5831 = n5819 ^ n5747;
  assign n5832 = n5831 ^ n5744;
  assign n5833 = n5832 ^ n3013;
  assign n5834 = n5816 ^ n5753;
  assign n5835 = n5834 ^ n5750;
  assign n5836 = n5835 ^ n3078;
  assign n5837 = n5813 ^ n5810;
  assign n5838 = n5837 ^ n3294;
  assign n5839 = n5806 ^ n5803;
  assign n5840 = n5839 ^ n3396;
  assign n5841 = n5799 ^ n5796;
  assign n5842 = n5841 ^ n3383;
  assign n5843 = n5791 ^ n5788;
  assign n5844 = n5843 ^ n3355;
  assign n5845 = n5783 ^ n5780;
  assign n5846 = n5845 ^ n3338;
  assign n5847 = n5775 ^ n5772;
  assign n5848 = n5847 ^ n3330;
  assign n5849 = n5767 ^ n5764;
  assign n5850 = n5849 ^ n3331;
  assign n5706 = n5705 ^ n5699;
  assign n5851 = n5706 ^ n3287;
  assign n5684 = n5683 ^ n5675;
  assign n5692 = n5684 ^ n3276;
  assign n5589 = n5588 ^ n5581;
  assign n5668 = n5589 ^ n3263;
  assign n5571 = n5570 ^ n5562;
  assign n5572 = n5571 ^ n3150;
  assign n5553 = n5552 ^ n5546;
  assign n5556 = n5553 ^ n3144;
  assign n5536 = n5535 ^ n5530;
  assign n5537 = n5536 ^ n3139;
  assign n5496 = n5495 ^ n5489;
  assign n5524 = n5496 ^ n3130;
  assign n5433 = n5432 ^ n5425;
  assign n5434 = n5433 ^ n3124;
  assign n5435 = n5422 ^ n4597;
  assign n5436 = n5435 ^ n3116;
  assign n5437 = n5419 ^ n4603;
  assign n5438 = n5437 ^ n3111;
  assign n5439 = n5416 ^ n4610;
  assign n5440 = n5439 ^ n3105;
  assign n5441 = n5413 ^ n4616;
  assign n5442 = n5441 ^ n3095;
  assign n5443 = n5410 ^ n4622;
  assign n5444 = n5443 ^ n3047;
  assign n5445 = n5407 ^ n5372;
  assign n5446 = n5445 ^ n3045;
  assign n5447 = n5404 ^ n5378;
  assign n5448 = n5447 ^ n3042;
  assign n5449 = n5401 ^ n5387;
  assign n5450 = n5449 ^ n2719;
  assign n5451 = n5397 ^ n5394;
  assign n5452 = n2723 & ~n5451;
  assign n5453 = n5452 ^ n3036;
  assign n5454 = n5398 ^ n5390;
  assign n5455 = n5454 ^ n5391;
  assign n5456 = n5455 ^ n5452;
  assign n5457 = n5453 & n5456;
  assign n5458 = n5457 ^ n3036;
  assign n5459 = n5458 ^ n5449;
  assign n5460 = ~n5450 & n5459;
  assign n5461 = n5460 ^ n2719;
  assign n5462 = n5461 ^ n5447;
  assign n5463 = ~n5448 & n5462;
  assign n5464 = n5463 ^ n3042;
  assign n5465 = n5464 ^ n5445;
  assign n5466 = n5446 & n5465;
  assign n5467 = n5466 ^ n3045;
  assign n5468 = n5467 ^ n5443;
  assign n5469 = n5444 & ~n5468;
  assign n5470 = n5469 ^ n3047;
  assign n5471 = n5470 ^ n5441;
  assign n5472 = ~n5442 & n5471;
  assign n5473 = n5472 ^ n3095;
  assign n5474 = n5473 ^ n5439;
  assign n5475 = n5440 & ~n5474;
  assign n5476 = n5475 ^ n3105;
  assign n5477 = n5476 ^ n5437;
  assign n5478 = ~n5438 & n5477;
  assign n5479 = n5478 ^ n3111;
  assign n5480 = n5479 ^ n5435;
  assign n5481 = n5436 & ~n5480;
  assign n5482 = n5481 ^ n3116;
  assign n5483 = n5482 ^ n5433;
  assign n5484 = ~n5434 & ~n5483;
  assign n5485 = n5484 ^ n3124;
  assign n5525 = n5496 ^ n5485;
  assign n5526 = ~n5524 & n5525;
  assign n5527 = n5526 ^ n3130;
  assign n5540 = n5536 ^ n5527;
  assign n5541 = ~n5537 & ~n5540;
  assign n5542 = n5541 ^ n3139;
  assign n5557 = n5553 ^ n5542;
  assign n5558 = n5556 & n5557;
  assign n5559 = n5558 ^ n3144;
  assign n5575 = n5571 ^ n5559;
  assign n5576 = n5572 & n5575;
  assign n5577 = n5576 ^ n3150;
  assign n5669 = n5589 ^ n5577;
  assign n5670 = n5668 & n5669;
  assign n5671 = n5670 ^ n3263;
  assign n5693 = n5684 ^ n5671;
  assign n5694 = n5692 & ~n5693;
  assign n5695 = n5694 ^ n3276;
  assign n5852 = n5706 ^ n5695;
  assign n5853 = n5851 & n5852;
  assign n5854 = n5853 ^ n3287;
  assign n5855 = n5854 ^ n5849;
  assign n5856 = ~n5850 & ~n5855;
  assign n5857 = n5856 ^ n3331;
  assign n5858 = n5857 ^ n5847;
  assign n5859 = ~n5848 & ~n5858;
  assign n5860 = n5859 ^ n3330;
  assign n5861 = n5860 ^ n5845;
  assign n5862 = n5846 & ~n5861;
  assign n5863 = n5862 ^ n3338;
  assign n5864 = n5863 ^ n5843;
  assign n5865 = n5844 & n5864;
  assign n5866 = n5865 ^ n3355;
  assign n5867 = n5866 ^ n5841;
  assign n5868 = ~n5842 & n5867;
  assign n5869 = n5868 ^ n3383;
  assign n5870 = n5869 ^ n5839;
  assign n5871 = ~n5840 & n5870;
  assign n5872 = n5871 ^ n3396;
  assign n5873 = n5872 ^ n5837;
  assign n5874 = ~n5838 & n5873;
  assign n5875 = n5874 ^ n3294;
  assign n5876 = n5875 ^ n5835;
  assign n5877 = n5836 & n5876;
  assign n5878 = n5877 ^ n3078;
  assign n5879 = n5878 ^ n5832;
  assign n5880 = n5833 & n5879;
  assign n5881 = n5880 ^ n3013;
  assign n5882 = n5881 ^ n5829;
  assign n5883 = n5830 & ~n5882;
  assign n5884 = n5883 ^ n3015;
  assign n5989 = n5894 ^ n5884;
  assign n5990 = ~n5895 & ~n5989;
  assign n5991 = n5990 ^ n3012;
  assign n6010 = n6002 ^ n5991;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = n6011 ^ n3028;
  assign n6023 = n6022 ^ n6012;
  assign n6024 = n6023 ^ n2724;
  assign n5896 = n5895 ^ n5884;
  assign n5897 = n5872 ^ n3294;
  assign n5898 = n5897 ^ n5837;
  assign n5899 = n5863 ^ n3355;
  assign n5900 = n5899 ^ n5843;
  assign n5901 = n5860 ^ n3338;
  assign n5902 = n5901 ^ n5845;
  assign n5903 = n5857 ^ n3330;
  assign n5904 = n5903 ^ n5847;
  assign n5696 = n5695 ^ n3287;
  assign n5707 = n5706 ^ n5696;
  assign n5486 = n5485 ^ n3130;
  assign n5497 = n5496 ^ n5486;
  assign n5498 = n5479 ^ n3116;
  assign n5499 = n5498 ^ n5435;
  assign n5500 = n5470 ^ n5442;
  assign n5501 = n5467 ^ n3047;
  assign n5502 = n5501 ^ n5443;
  assign n5503 = n5464 ^ n5446;
  assign n5504 = n5461 ^ n3042;
  assign n5505 = n5504 ^ n5447;
  assign n5506 = n5458 ^ n5450;
  assign n5507 = n5451 ^ n2723;
  assign n5508 = n5455 ^ n5453;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~n5506 & n5509;
  assign n5511 = n5505 & ~n5510;
  assign n5512 = ~n5503 & n5511;
  assign n5513 = ~n5502 & ~n5512;
  assign n5514 = n5500 & n5513;
  assign n5515 = n5473 ^ n3105;
  assign n5516 = n5515 ^ n5439;
  assign n5517 = ~n5514 & n5516;
  assign n5518 = n5476 ^ n5438;
  assign n5519 = n5517 & ~n5518;
  assign n5520 = ~n5499 & ~n5519;
  assign n5521 = n5482 ^ n5434;
  assign n5522 = n5520 & n5521;
  assign n5523 = n5497 & ~n5522;
  assign n5538 = n5537 ^ n5527;
  assign n5539 = n5523 & n5538;
  assign n5543 = n5542 ^ n3144;
  assign n5554 = n5553 ^ n5543;
  assign n5555 = n5539 & n5554;
  assign n5573 = n5572 ^ n5559;
  assign n5574 = n5555 & ~n5573;
  assign n5578 = n5577 ^ n3263;
  assign n5590 = n5589 ^ n5578;
  assign n5667 = ~n5574 & ~n5590;
  assign n5672 = n5671 ^ n3276;
  assign n5685 = n5684 ^ n5672;
  assign n5708 = n5667 & n5685;
  assign n5905 = ~n5707 & ~n5708;
  assign n5906 = n5854 ^ n3331;
  assign n5907 = n5906 ^ n5849;
  assign n5908 = ~n5905 & n5907;
  assign n5909 = ~n5904 & n5908;
  assign n5910 = ~n5902 & n5909;
  assign n5911 = ~n5900 & n5910;
  assign n5912 = n5866 ^ n3383;
  assign n5913 = n5912 ^ n5841;
  assign n5914 = n5911 & ~n5913;
  assign n5915 = n5869 ^ n3396;
  assign n5916 = n5915 ^ n5839;
  assign n5917 = ~n5914 & n5916;
  assign n5918 = ~n5898 & ~n5917;
  assign n5919 = n5875 ^ n3078;
  assign n5920 = n5919 ^ n5835;
  assign n5921 = ~n5918 & ~n5920;
  assign n5922 = n5878 ^ n3013;
  assign n5923 = n5922 ^ n5832;
  assign n5924 = ~n5921 & ~n5923;
  assign n5925 = n5881 ^ n3015;
  assign n5926 = n5925 ^ n5829;
  assign n5927 = ~n5924 & ~n5926;
  assign n5988 = n5896 & n5927;
  assign n5992 = n5991 ^ n3028;
  assign n6003 = n6002 ^ n5992;
  assign n6025 = ~n5988 & n6003;
  assign n6044 = ~n6024 & ~n6025;
  assign n6040 = n5327 ^ n5180;
  assign n6037 = n3772 ^ n3323;
  assign n6038 = n4565 & ~n6037;
  assign n6039 = n6038 ^ n3323;
  assign n6041 = n6040 ^ n6039;
  assign n6034 = n6017 ^ n6015;
  assign n6035 = n6021 & n6034;
  assign n6036 = n6035 ^ n6015;
  assign n6042 = n6041 ^ n6036;
  assign n6043 = n6042 ^ n3033;
  assign n6045 = n6044 ^ n6043;
  assign n6031 = n6022 ^ n2724;
  assign n6032 = n6023 & n6031;
  assign n6033 = n6032 ^ n2724;
  assign n6046 = n6045 ^ n6033;
  assign n5928 = n5927 ^ n5896;
  assign n5929 = n5928 ^ x195;
  assign n5930 = n5923 ^ n5921;
  assign n5931 = n5930 ^ x197;
  assign n5932 = n5920 ^ n5918;
  assign n5933 = n5932 ^ x198;
  assign n5934 = n5917 ^ n5898;
  assign n5935 = n5934 ^ x199;
  assign n5936 = n5916 ^ n5914;
  assign n5937 = n5936 ^ x200;
  assign n5938 = n5913 ^ n5911;
  assign n5939 = n5938 ^ x201;
  assign n5940 = n5910 ^ n5900;
  assign n5941 = n5940 ^ x202;
  assign n5942 = n5909 ^ n5902;
  assign n5943 = n5942 ^ x203;
  assign n5944 = n5908 ^ n5904;
  assign n5945 = n5944 ^ x204;
  assign n5946 = n5907 ^ n5905;
  assign n5947 = n5946 ^ x205;
  assign n5709 = n5708 ^ n5707;
  assign n5948 = n5709 ^ x206;
  assign n5686 = n5685 ^ n5667;
  assign n5591 = n5590 ^ n5574;
  assign n5592 = n5591 ^ x208;
  assign n5593 = n5573 ^ n5555;
  assign n5594 = n5593 ^ x209;
  assign n5595 = n5554 ^ n5539;
  assign n5596 = n5595 ^ x210;
  assign n5597 = n5538 ^ n5523;
  assign n5598 = n5597 ^ x211;
  assign n5599 = n5522 ^ n5497;
  assign n5600 = n5599 ^ x212;
  assign n5601 = n5521 ^ n5520;
  assign n5602 = n5601 ^ x213;
  assign n5603 = n5519 ^ n5499;
  assign n5604 = n5603 ^ x214;
  assign n5605 = n5518 ^ n5517;
  assign n5606 = n5605 ^ x215;
  assign n5607 = n5516 ^ n5514;
  assign n5608 = n5607 ^ x216;
  assign n5609 = n5513 ^ n5500;
  assign n5610 = n5609 ^ x217;
  assign n5611 = n5512 ^ n5502;
  assign n5612 = n5611 ^ x218;
  assign n5613 = n5511 ^ n5503;
  assign n5614 = n5613 ^ x219;
  assign n5615 = n5510 ^ n5505;
  assign n5616 = n5615 ^ x220;
  assign n5617 = n5509 ^ n5506;
  assign n5618 = n5617 ^ x221;
  assign n5619 = x223 & n5507;
  assign n5620 = n5619 ^ x222;
  assign n5621 = n5508 ^ n5507;
  assign n5622 = n5621 ^ n5619;
  assign n5623 = n5620 & ~n5622;
  assign n5624 = n5623 ^ x222;
  assign n5625 = n5624 ^ n5617;
  assign n5626 = ~n5618 & n5625;
  assign n5627 = n5626 ^ x221;
  assign n5628 = n5627 ^ n5615;
  assign n5629 = n5616 & ~n5628;
  assign n5630 = n5629 ^ x220;
  assign n5631 = n5630 ^ n5613;
  assign n5632 = n5614 & ~n5631;
  assign n5633 = n5632 ^ x219;
  assign n5634 = n5633 ^ n5611;
  assign n5635 = n5612 & ~n5634;
  assign n5636 = n5635 ^ x218;
  assign n5637 = n5636 ^ n5609;
  assign n5638 = n5610 & ~n5637;
  assign n5639 = n5638 ^ x217;
  assign n5640 = n5639 ^ n5607;
  assign n5641 = n5608 & ~n5640;
  assign n5642 = n5641 ^ x216;
  assign n5643 = n5642 ^ n5605;
  assign n5644 = n5606 & ~n5643;
  assign n5645 = n5644 ^ x215;
  assign n5646 = n5645 ^ n5603;
  assign n5647 = n5604 & ~n5646;
  assign n5648 = n5647 ^ x214;
  assign n5649 = n5648 ^ n5601;
  assign n5650 = n5602 & ~n5649;
  assign n5651 = n5650 ^ x213;
  assign n5652 = n5651 ^ n5599;
  assign n5653 = n5600 & ~n5652;
  assign n5654 = n5653 ^ x212;
  assign n5655 = n5654 ^ n5597;
  assign n5656 = ~n5598 & n5655;
  assign n5657 = n5656 ^ x211;
  assign n5658 = n5657 ^ n5595;
  assign n5659 = ~n5596 & n5658;
  assign n5660 = n5659 ^ x210;
  assign n5661 = n5660 ^ n5593;
  assign n5662 = n5594 & ~n5661;
  assign n5663 = n5662 ^ x209;
  assign n5664 = n5663 ^ n5591;
  assign n5665 = n5592 & ~n5664;
  assign n5666 = n5665 ^ x208;
  assign n5687 = n5686 ^ n5666;
  assign n5688 = n5686 ^ x207;
  assign n5689 = ~n5687 & n5688;
  assign n5690 = n5689 ^ x207;
  assign n5949 = n5709 ^ n5690;
  assign n5950 = ~n5948 & n5949;
  assign n5951 = n5950 ^ x206;
  assign n5952 = n5951 ^ n5946;
  assign n5953 = ~n5947 & n5952;
  assign n5954 = n5953 ^ x205;
  assign n5955 = n5954 ^ n5944;
  assign n5956 = ~n5945 & n5955;
  assign n5957 = n5956 ^ x204;
  assign n5958 = n5957 ^ n5942;
  assign n5959 = ~n5943 & n5958;
  assign n5960 = n5959 ^ x203;
  assign n5961 = n5960 ^ n5940;
  assign n5962 = ~n5941 & n5961;
  assign n5963 = n5962 ^ x202;
  assign n5964 = n5963 ^ n5938;
  assign n5965 = ~n5939 & n5964;
  assign n5966 = n5965 ^ x201;
  assign n5967 = n5966 ^ n5936;
  assign n5968 = n5937 & ~n5967;
  assign n5969 = n5968 ^ x200;
  assign n5970 = n5969 ^ n5934;
  assign n5971 = n5935 & ~n5970;
  assign n5972 = n5971 ^ x199;
  assign n5973 = n5972 ^ n5932;
  assign n5974 = ~n5933 & n5973;
  assign n5975 = n5974 ^ x198;
  assign n5976 = n5975 ^ n5930;
  assign n5977 = n5931 & ~n5976;
  assign n5978 = n5977 ^ x197;
  assign n5979 = n5978 ^ x196;
  assign n5980 = n5926 ^ n5924;
  assign n5981 = n5980 ^ n5978;
  assign n5982 = n5979 & n5981;
  assign n5983 = n5982 ^ x196;
  assign n5984 = n5983 ^ n5928;
  assign n5985 = ~n5929 & n5984;
  assign n5986 = n5985 ^ x195;
  assign n5987 = n5986 ^ x194;
  assign n6004 = n6003 ^ n5988;
  assign n6005 = n6004 ^ n5986;
  assign n6006 = n5987 & n6005;
  assign n6007 = n6006 ^ x194;
  assign n6008 = n6007 ^ x193;
  assign n6026 = n6025 ^ n6024;
  assign n6027 = n6026 ^ n6007;
  assign n6028 = n6008 & n6027;
  assign n6029 = n6028 ^ x193;
  assign n6030 = n6029 ^ x192;
  assign n6047 = n6046 ^ n6030;
  assign n5741 = n4612 ^ n4041;
  assign n5742 = n4588 & n5741;
  assign n5743 = n5742 ^ n4041;
  assign n6048 = n6047 ^ n5743;
  assign n6052 = n6026 ^ n6008;
  assign n6049 = n4618 ^ n3758;
  assign n6050 = n4598 & n6049;
  assign n6051 = n6050 ^ n3758;
  assign n6053 = n6052 ^ n6051;
  assign n6057 = n6004 ^ n5987;
  assign n6054 = n4623 ^ n4030;
  assign n6055 = ~n4609 & ~n6054;
  assign n6056 = n6055 ^ n4030;
  assign n6058 = n6057 ^ n6056;
  assign n6060 = n4694 ^ n3761;
  assign n6061 = ~n4611 & n6060;
  assign n6062 = n6061 ^ n3761;
  assign n6059 = n5983 ^ n5929;
  assign n6063 = n6062 ^ n6059;
  assign n6064 = n5980 ^ n5979;
  assign n6065 = n4667 ^ n3770;
  assign n6066 = n4617 & ~n6065;
  assign n6067 = n6066 ^ n3770;
  assign n6068 = ~n6064 & ~n6067;
  assign n6069 = n6068 ^ n6059;
  assign n6070 = n6063 & ~n6069;
  assign n6071 = n6070 ^ n6068;
  assign n6072 = n6071 ^ n6057;
  assign n6073 = ~n6058 & n6072;
  assign n6074 = n6073 ^ n6056;
  assign n6075 = n6074 ^ n6052;
  assign n6076 = ~n6053 & n6075;
  assign n6077 = n6076 ^ n6051;
  assign n6078 = n6077 ^ n6047;
  assign n6079 = ~n6048 & n6078;
  assign n6080 = n6079 ^ n5743;
  assign n5739 = n5507 ^ x223;
  assign n5736 = n4604 ^ n3750;
  assign n5737 = n5431 & ~n5736;
  assign n5738 = n5737 ^ n3750;
  assign n5740 = n5739 ^ n5738;
  assign n6112 = n6080 ^ n5740;
  assign n6113 = n6112 ^ n3304;
  assign n6114 = n6077 ^ n6048;
  assign n6115 = n6114 ^ n3307;
  assign n6116 = n6074 ^ n6053;
  assign n6117 = n6116 ^ n3311;
  assign n6118 = n6071 ^ n6058;
  assign n6119 = n6118 ^ n3314;
  assign n6120 = n6067 ^ n6064;
  assign n6121 = ~n3321 & n6120;
  assign n6122 = n6121 ^ n3317;
  assign n6123 = n6068 ^ n6062;
  assign n6124 = n6123 ^ n6059;
  assign n6125 = n6124 ^ n6121;
  assign n6126 = n6122 & n6125;
  assign n6127 = n6126 ^ n3317;
  assign n6128 = n6127 ^ n6118;
  assign n6129 = ~n6119 & n6128;
  assign n6130 = n6129 ^ n3314;
  assign n6131 = n6130 ^ n6116;
  assign n6132 = n6117 & n6131;
  assign n6133 = n6132 ^ n3311;
  assign n6134 = n6133 ^ n6114;
  assign n6135 = ~n6115 & ~n6134;
  assign n6136 = n6135 ^ n3307;
  assign n6137 = n6136 ^ n6112;
  assign n6138 = ~n6113 & ~n6137;
  assign n6139 = n6138 ^ n3304;
  assign n6181 = n6139 ^ n3301;
  assign n6081 = n6080 ^ n5739;
  assign n6082 = n5740 & ~n6081;
  assign n6083 = n6082 ^ n5738;
  assign n5732 = n4599 ^ n3742;
  assign n5733 = ~n5494 & n5732;
  assign n5734 = n5733 ^ n3742;
  assign n5731 = n5621 ^ n5620;
  assign n5735 = n5734 ^ n5731;
  assign n6110 = n6083 ^ n5735;
  assign n6182 = n6181 ^ n6110;
  assign n6168 = n6133 ^ n3307;
  assign n6169 = n6168 ^ n6114;
  assign n6170 = n6130 ^ n6117;
  assign n6171 = n6127 ^ n3314;
  assign n6172 = n6171 ^ n6118;
  assign n6173 = n6120 ^ n3321;
  assign n6174 = n6124 ^ n6122;
  assign n6175 = ~n6173 & ~n6174;
  assign n6176 = ~n6172 & n6175;
  assign n6177 = ~n6170 & ~n6176;
  assign n6178 = ~n6169 & n6177;
  assign n6179 = n6136 ^ n6113;
  assign n6180 = ~n6178 & ~n6179;
  assign n6202 = n6182 ^ n6180;
  assign n6203 = n6202 ^ x249;
  assign n6204 = n6179 ^ n6178;
  assign n6205 = n6204 ^ x250;
  assign n6206 = n6177 ^ n6169;
  assign n6207 = n6206 ^ x251;
  assign n6208 = n6176 ^ n6170;
  assign n6209 = n6208 ^ x252;
  assign n6210 = n6175 ^ n6172;
  assign n6211 = n6210 ^ x253;
  assign n6212 = x255 & n6173;
  assign n6213 = n6212 ^ x254;
  assign n6214 = n6174 ^ n6173;
  assign n6215 = n6214 ^ n6212;
  assign n6216 = n6213 & ~n6215;
  assign n6217 = n6216 ^ x254;
  assign n6218 = n6217 ^ n6210;
  assign n6219 = ~n6211 & n6218;
  assign n6220 = n6219 ^ x253;
  assign n6221 = n6220 ^ n6208;
  assign n6222 = ~n6209 & n6221;
  assign n6223 = n6222 ^ x252;
  assign n6224 = n6223 ^ n6206;
  assign n6225 = n6207 & ~n6224;
  assign n6226 = n6225 ^ x251;
  assign n6227 = n6226 ^ n6204;
  assign n6228 = n6205 & ~n6227;
  assign n6229 = n6228 ^ x250;
  assign n6230 = n6229 ^ n6202;
  assign n6231 = ~n6203 & n6230;
  assign n6232 = n6231 ^ x249;
  assign n6301 = n6232 ^ x248;
  assign n6111 = n6110 ^ n3301;
  assign n6140 = n6139 ^ n6110;
  assign n6141 = n6111 & n6140;
  assign n6142 = n6141 ^ n3301;
  assign n6084 = n6083 ^ n5731;
  assign n6085 = n5735 & ~n6084;
  assign n6086 = n6085 ^ n5734;
  assign n5727 = n4593 ^ n3737;
  assign n5728 = ~n5534 & n5727;
  assign n5729 = n5728 ^ n3737;
  assign n5726 = n5624 ^ n5618;
  assign n5730 = n5729 ^ n5726;
  assign n6108 = n6086 ^ n5730;
  assign n6109 = n6108 ^ n3299;
  assign n6184 = n6142 ^ n6109;
  assign n6183 = n6180 & ~n6182;
  assign n6200 = n6184 ^ n6183;
  assign n6302 = n6301 ^ n6200;
  assign n6297 = n5654 ^ n5598;
  assign n6298 = n5771 ^ n4758;
  assign n6299 = ~n6297 & n6298;
  assign n6300 = n6299 ^ n4758;
  assign n6303 = n6302 ^ n6300;
  assign n6305 = n5651 ^ x212;
  assign n6306 = n6305 ^ n5599;
  assign n6307 = n5763 ^ n4734;
  assign n6308 = n6306 & ~n6307;
  assign n6309 = n6308 ^ n4734;
  assign n6304 = n6229 ^ n6203;
  assign n6310 = n6309 ^ n6304;
  assign n6315 = n6226 ^ x250;
  assign n6316 = n6315 ^ n6204;
  assign n6311 = n5648 ^ n5602;
  assign n6312 = n5704 ^ n4739;
  assign n6313 = n6311 & ~n6312;
  assign n6314 = n6313 ^ n4739;
  assign n6317 = n6316 ^ n6314;
  assign n6319 = n5645 ^ n5604;
  assign n6320 = n5682 ^ n4750;
  assign n6321 = n6319 & n6320;
  assign n6322 = n6321 ^ n4750;
  assign n6318 = n6223 ^ n6207;
  assign n6323 = n6322 ^ n6318;
  assign n6329 = n6220 ^ x252;
  assign n6330 = n6329 ^ n6208;
  assign n6324 = n5642 ^ x215;
  assign n6325 = n6324 ^ n5605;
  assign n6326 = n5587 ^ n4645;
  assign n6327 = n6325 & ~n6326;
  assign n6328 = n6327 ^ n4645;
  assign n6331 = n6330 ^ n6328;
  assign n6335 = n6217 ^ n6211;
  assign n6261 = n5639 ^ x216;
  assign n6262 = n6261 ^ n5607;
  assign n6332 = n5569 ^ n4593;
  assign n6333 = n6262 & ~n6332;
  assign n6334 = n6333 ^ n4593;
  assign n6336 = n6335 ^ n6334;
  assign n6340 = n6214 ^ n6213;
  assign n6162 = n5636 ^ n5610;
  assign n6337 = n5551 ^ n4599;
  assign n6338 = n6162 & n6337;
  assign n6339 = n6338 ^ n4599;
  assign n6341 = n6340 ^ n6339;
  assign n6099 = n5633 ^ x218;
  assign n6100 = n6099 ^ n5611;
  assign n6343 = n5534 ^ n4604;
  assign n6344 = n6100 & n6343;
  assign n6345 = n6344 ^ n4604;
  assign n6342 = n6173 ^ x255;
  assign n6346 = n6345 ^ n6342;
  assign n5718 = n5630 ^ n5614;
  assign n6751 = n5494 ^ n4612;
  assign n6752 = n5718 & ~n6751;
  assign n6753 = n6752 ^ n4612;
  assign n5723 = n5627 ^ x220;
  assign n5724 = n5723 ^ n5615;
  assign n6721 = n5431 ^ n4618;
  assign n6722 = n5724 & n6721;
  assign n6723 = n6722 ^ n4618;
  assign n6538 = n5963 ^ n5939;
  assign n6534 = n4480 ^ n4007;
  assign n6535 = n5394 & ~n6534;
  assign n6536 = n6535 ^ n4007;
  assign n6450 = n5960 ^ x202;
  assign n6451 = n6450 ^ n5940;
  assign n6446 = n4445 ^ n3990;
  assign n6447 = ~n6040 & n6446;
  assign n6448 = n6447 ^ n3990;
  assign n6530 = n6451 ^ n6448;
  assign n6348 = n4411 ^ n3998;
  assign n6349 = n6017 & n6348;
  assign n6350 = n6349 ^ n3998;
  assign n6347 = n5957 ^ n5943;
  assign n6351 = n6350 ^ n6347;
  assign n6354 = n5364 ^ n4554;
  assign n6355 = n5996 & n6354;
  assign n6356 = n6355 ^ n4554;
  assign n6352 = n5954 ^ x204;
  assign n6353 = n6352 ^ n5944;
  assign n6357 = n6356 ^ n6353;
  assign n6359 = n5066 ^ n4506;
  assign n6360 = ~n5886 & ~n6359;
  assign n6361 = n6360 ^ n4506;
  assign n6358 = n5951 ^ n5947;
  assign n6362 = n6361 ^ n6358;
  assign n6363 = n4876 ^ n4470;
  assign n6364 = ~n5824 & n6363;
  assign n6365 = n6364 ^ n4470;
  assign n5691 = n5690 ^ x206;
  assign n5710 = n5709 ^ n5691;
  assign n6366 = n6365 ^ n5710;
  assign n6367 = n4638 ^ n4438;
  assign n6368 = n5744 & n6367;
  assign n6369 = n6368 ^ n4438;
  assign n6269 = n5687 ^ x207;
  assign n6370 = n6369 ^ n6269;
  assign n6371 = n4845 ^ n4404;
  assign n6372 = n5750 & ~n6371;
  assign n6373 = n6372 ^ n4404;
  assign n6276 = n5663 ^ x208;
  assign n6277 = n6276 ^ n5591;
  assign n6374 = n6373 ^ n6277;
  assign n6375 = n4830 ^ n4115;
  assign n6376 = ~n5711 & n6375;
  assign n6377 = n6376 ^ n4115;
  assign n6283 = n5660 ^ n5594;
  assign n6378 = n6377 ^ n6283;
  assign n6379 = n4840 ^ n4100;
  assign n6380 = ~n5755 & ~n6379;
  assign n6381 = n6380 ^ n4100;
  assign n6291 = n5657 ^ x210;
  assign n6292 = n6291 ^ n5595;
  assign n6382 = n6381 ^ n6292;
  assign n6383 = n4838 ^ n3673;
  assign n6384 = n5795 & n6383;
  assign n6385 = n6384 ^ n3673;
  assign n6386 = n6385 ^ n6297;
  assign n6387 = n4786 ^ n3679;
  assign n6388 = ~n5787 & n6387;
  assign n6389 = n6388 ^ n3679;
  assign n6390 = n6389 ^ n6306;
  assign n6391 = n4779 ^ n4083;
  assign n6392 = ~n5779 & n6391;
  assign n6393 = n6392 ^ n4083;
  assign n6394 = n6393 ^ n6311;
  assign n6395 = n4775 ^ n3686;
  assign n6396 = n5771 & n6395;
  assign n6397 = n6396 ^ n3686;
  assign n6398 = n6397 ^ n6319;
  assign n6399 = n4766 ^ n3692;
  assign n6400 = n5763 & n6399;
  assign n6401 = n6400 ^ n3692;
  assign n6402 = n6401 ^ n6325;
  assign n6257 = n4758 ^ n3698;
  assign n6258 = n5704 & n6257;
  assign n6259 = n6258 ^ n3698;
  assign n6403 = n6262 ^ n6259;
  assign n6158 = n4734 ^ n3708;
  assign n6159 = ~n5682 & n6158;
  assign n6160 = n6159 ^ n3708;
  assign n6253 = n6162 ^ n6160;
  assign n6096 = n4739 ^ n3711;
  assign n6097 = ~n5587 & ~n6096;
  assign n6098 = n6097 ^ n3711;
  assign n6101 = n6100 ^ n6098;
  assign n5715 = n4750 ^ n3722;
  assign n5716 = ~n5569 & n5715;
  assign n5717 = n5716 ^ n3722;
  assign n5719 = n5718 ^ n5717;
  assign n5720 = n4645 ^ n3732;
  assign n5721 = n5551 & ~n5720;
  assign n5722 = n5721 ^ n3732;
  assign n5725 = n5724 ^ n5722;
  assign n6087 = n6086 ^ n5726;
  assign n6088 = ~n5730 & n6087;
  assign n6089 = n6088 ^ n5729;
  assign n6090 = n6089 ^ n5724;
  assign n6091 = ~n5725 & ~n6090;
  assign n6092 = n6091 ^ n5722;
  assign n6093 = n6092 ^ n5718;
  assign n6094 = ~n5719 & n6093;
  assign n6095 = n6094 ^ n5717;
  assign n6155 = n6100 ^ n6095;
  assign n6156 = n6101 & n6155;
  assign n6157 = n6156 ^ n6098;
  assign n6254 = n6162 ^ n6157;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = n6255 ^ n6160;
  assign n6404 = n6262 ^ n6256;
  assign n6405 = n6403 & n6404;
  assign n6406 = n6405 ^ n6259;
  assign n6407 = n6406 ^ n6325;
  assign n6408 = n6402 & ~n6407;
  assign n6409 = n6408 ^ n6401;
  assign n6410 = n6409 ^ n6319;
  assign n6411 = ~n6398 & ~n6410;
  assign n6412 = n6411 ^ n6397;
  assign n6413 = n6412 ^ n6311;
  assign n6414 = n6394 & n6413;
  assign n6415 = n6414 ^ n6393;
  assign n6416 = n6415 ^ n6306;
  assign n6417 = ~n6390 & ~n6416;
  assign n6418 = n6417 ^ n6389;
  assign n6419 = n6418 ^ n6297;
  assign n6420 = n6386 & ~n6419;
  assign n6421 = n6420 ^ n6385;
  assign n6422 = n6421 ^ n6292;
  assign n6423 = ~n6382 & ~n6422;
  assign n6424 = n6423 ^ n6381;
  assign n6425 = n6424 ^ n6283;
  assign n6426 = n6378 & ~n6425;
  assign n6427 = n6426 ^ n6377;
  assign n6428 = n6427 ^ n6277;
  assign n6429 = n6374 & ~n6428;
  assign n6430 = n6429 ^ n6373;
  assign n6431 = n6430 ^ n6269;
  assign n6432 = n6370 & ~n6431;
  assign n6433 = n6432 ^ n6369;
  assign n6434 = n6433 ^ n5710;
  assign n6435 = ~n6366 & n6434;
  assign n6436 = n6435 ^ n6365;
  assign n6437 = n6436 ^ n6358;
  assign n6438 = n6362 & n6437;
  assign n6439 = n6438 ^ n6361;
  assign n6440 = n6439 ^ n6353;
  assign n6441 = ~n6357 & ~n6440;
  assign n6442 = n6441 ^ n6356;
  assign n6443 = n6442 ^ n6347;
  assign n6444 = ~n6351 & n6443;
  assign n6445 = n6444 ^ n6350;
  assign n6531 = n6451 ^ n6445;
  assign n6532 = ~n6530 & n6531;
  assign n6533 = n6532 ^ n6448;
  assign n6537 = n6536 ^ n6533;
  assign n6539 = n6538 ^ n6537;
  assign n6449 = n6448 ^ n6445;
  assign n6452 = n6451 ^ n6449;
  assign n6453 = n6452 ^ n3428;
  assign n6454 = n6442 ^ n6351;
  assign n6455 = n6454 ^ n3423;
  assign n6456 = n6439 ^ n6357;
  assign n6457 = n6456 ^ n3973;
  assign n6458 = n6436 ^ n6362;
  assign n6459 = n6458 ^ n3862;
  assign n6460 = n6433 ^ n6366;
  assign n6461 = n6460 ^ n3293;
  assign n6462 = n6430 ^ n6370;
  assign n6463 = n6462 ^ n3675;
  assign n6464 = n6427 ^ n6374;
  assign n6465 = n6464 ^ n3823;
  assign n6466 = n6424 ^ n6378;
  assign n6467 = n6466 ^ n3681;
  assign n6468 = n6421 ^ n6382;
  assign n6469 = n6468 ^ n3688;
  assign n6470 = n6418 ^ n6386;
  assign n6471 = n6470 ^ n3694;
  assign n6472 = n6415 ^ n6390;
  assign n6473 = n6472 ^ n3700;
  assign n6474 = n6412 ^ n6393;
  assign n6475 = n6474 ^ n6311;
  assign n6476 = n6475 ^ n3712;
  assign n6477 = n6409 ^ n6397;
  assign n6478 = n6477 ^ n6319;
  assign n6479 = n6478 ^ n3723;
  assign n6480 = n6406 ^ n6401;
  assign n6481 = n6480 ^ n6325;
  assign n6482 = n6481 ^ n3728;
  assign n6260 = n6259 ^ n6256;
  assign n6263 = n6262 ^ n6260;
  assign n6483 = n6263 ^ n3667;
  assign n6161 = n6160 ^ n6157;
  assign n6163 = n6162 ^ n6161;
  assign n6164 = n6163 ^ n3557;
  assign n6102 = n6101 ^ n6095;
  assign n6103 = n6102 ^ n3546;
  assign n6104 = n6092 ^ n5719;
  assign n6105 = n6104 ^ n3506;
  assign n6106 = n6089 ^ n5725;
  assign n6107 = n6106 ^ n3472;
  assign n6143 = n6142 ^ n6108;
  assign n6144 = ~n6109 & n6143;
  assign n6145 = n6144 ^ n3299;
  assign n6146 = n6145 ^ n6106;
  assign n6147 = ~n6107 & n6146;
  assign n6148 = n6147 ^ n3472;
  assign n6149 = n6148 ^ n6104;
  assign n6150 = ~n6105 & ~n6149;
  assign n6151 = n6150 ^ n3506;
  assign n6152 = n6151 ^ n6102;
  assign n6153 = ~n6103 & ~n6152;
  assign n6154 = n6153 ^ n3546;
  assign n6249 = n6163 ^ n6154;
  assign n6250 = ~n6164 & n6249;
  assign n6251 = n6250 ^ n3557;
  assign n6484 = n6263 ^ n6251;
  assign n6485 = n6483 & n6484;
  assign n6486 = n6485 ^ n3667;
  assign n6487 = n6486 ^ n6481;
  assign n6488 = ~n6482 & n6487;
  assign n6489 = n6488 ^ n3728;
  assign n6490 = n6489 ^ n6478;
  assign n6491 = n6479 & ~n6490;
  assign n6492 = n6491 ^ n3723;
  assign n6493 = n6492 ^ n6475;
  assign n6494 = ~n6476 & ~n6493;
  assign n6495 = n6494 ^ n3712;
  assign n6496 = n6495 ^ n6472;
  assign n6497 = n6473 & n6496;
  assign n6498 = n6497 ^ n3700;
  assign n6499 = n6498 ^ n6470;
  assign n6500 = ~n6471 & ~n6499;
  assign n6501 = n6500 ^ n3694;
  assign n6502 = n6501 ^ n6468;
  assign n6503 = ~n6469 & ~n6502;
  assign n6504 = n6503 ^ n3688;
  assign n6505 = n6504 ^ n6466;
  assign n6506 = ~n6467 & n6505;
  assign n6507 = n6506 ^ n3681;
  assign n6508 = n6507 ^ n6464;
  assign n6509 = ~n6465 & n6508;
  assign n6510 = n6509 ^ n3823;
  assign n6511 = n6510 ^ n6462;
  assign n6512 = n6463 & n6511;
  assign n6513 = n6512 ^ n3675;
  assign n6514 = n6513 ^ n6460;
  assign n6515 = n6461 & n6514;
  assign n6516 = n6515 ^ n3293;
  assign n6517 = n6516 ^ n6458;
  assign n6518 = ~n6459 & n6517;
  assign n6519 = n6518 ^ n3862;
  assign n6520 = n6519 ^ n6456;
  assign n6521 = ~n6457 & n6520;
  assign n6522 = n6521 ^ n3973;
  assign n6523 = n6522 ^ n6454;
  assign n6524 = ~n6455 & ~n6523;
  assign n6525 = n6524 ^ n3423;
  assign n6526 = n6525 ^ n6452;
  assign n6527 = ~n6453 & n6526;
  assign n6528 = n6527 ^ n3428;
  assign n6529 = n6528 ^ n3420;
  assign n6540 = n6539 ^ n6529;
  assign n6541 = n6501 ^ n3688;
  assign n6542 = n6541 ^ n6468;
  assign n6543 = n6498 ^ n6471;
  assign n6544 = n6489 ^ n3723;
  assign n6545 = n6544 ^ n6478;
  assign n6546 = n6486 ^ n3728;
  assign n6547 = n6546 ^ n6481;
  assign n6165 = n6164 ^ n6154;
  assign n6166 = n6151 ^ n3546;
  assign n6167 = n6166 ^ n6102;
  assign n6185 = ~n6183 & n6184;
  assign n6186 = n6145 ^ n3472;
  assign n6187 = n6186 ^ n6106;
  assign n6188 = n6185 & n6187;
  assign n6189 = n6148 ^ n6105;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = n6167 & n6190;
  assign n6248 = n6165 & ~n6191;
  assign n6252 = n6251 ^ n3667;
  assign n6264 = n6263 ^ n6252;
  assign n6548 = n6248 & ~n6264;
  assign n6549 = ~n6547 & n6548;
  assign n6550 = n6545 & n6549;
  assign n6551 = n6492 ^ n3712;
  assign n6552 = n6551 ^ n6475;
  assign n6553 = ~n6550 & n6552;
  assign n6554 = n6495 ^ n6473;
  assign n6555 = n6553 & n6554;
  assign n6556 = ~n6543 & ~n6555;
  assign n6557 = ~n6542 & ~n6556;
  assign n6558 = n6504 ^ n6467;
  assign n6559 = n6557 & n6558;
  assign n6560 = n6507 ^ n3823;
  assign n6561 = n6560 ^ n6464;
  assign n6562 = n6559 & n6561;
  assign n6563 = n6510 ^ n6463;
  assign n6564 = n6562 & ~n6563;
  assign n6565 = n6513 ^ n3293;
  assign n6566 = n6565 ^ n6460;
  assign n6567 = n6564 & n6566;
  assign n6568 = n6516 ^ n6459;
  assign n6569 = ~n6567 & ~n6568;
  assign n6570 = n6519 ^ n6457;
  assign n6571 = ~n6569 & n6570;
  assign n6572 = n6522 ^ n6455;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = n6525 ^ n3428;
  assign n6575 = n6574 ^ n6452;
  assign n6576 = ~n6573 & ~n6575;
  assign n6577 = n6540 & ~n6576;
  assign n6591 = n5966 ^ x200;
  assign n6592 = n6591 ^ n5936;
  assign n6587 = n4520 ^ n3987;
  assign n6588 = ~n5391 & n6587;
  assign n6589 = n6588 ^ n3987;
  assign n6583 = n6538 ^ n6536;
  assign n6584 = n6538 ^ n6533;
  assign n6585 = n6583 & n6584;
  assign n6586 = n6585 ^ n6536;
  assign n6590 = n6589 ^ n6586;
  assign n6593 = n6592 ^ n6590;
  assign n6578 = n6539 ^ n3420;
  assign n6579 = n6539 ^ n6528;
  assign n6580 = ~n6578 & ~n6579;
  assign n6581 = n6580 ^ n3420;
  assign n6582 = n6581 ^ n3416;
  assign n6594 = n6593 ^ n6582;
  assign n6595 = n6577 & ~n6594;
  assign n6608 = n5969 ^ x199;
  assign n6609 = n6608 ^ n5934;
  assign n6604 = n6592 ^ n6589;
  assign n6605 = n6592 ^ n6586;
  assign n6606 = n6604 & n6605;
  assign n6607 = n6606 ^ n6589;
  assign n6610 = n6609 ^ n6607;
  assign n6601 = n4565 ^ n3977;
  assign n6602 = ~n5383 & n6601;
  assign n6603 = n6602 ^ n3977;
  assign n6611 = n6610 ^ n6603;
  assign n6596 = n6593 ^ n3416;
  assign n6597 = n6593 ^ n6581;
  assign n6598 = ~n6596 & ~n6597;
  assign n6599 = n6598 ^ n3416;
  assign n6600 = n6599 ^ n3413;
  assign n6612 = n6611 ^ n6600;
  assign n6718 = ~n6595 & ~n6612;
  assign n6713 = n5972 ^ x198;
  assign n6714 = n6713 ^ n5932;
  assign n6710 = n6609 ^ n6603;
  assign n6711 = ~n6610 & n6710;
  assign n6712 = n6711 ^ n6603;
  assign n6715 = n6714 ^ n6712;
  assign n6707 = n4680 ^ n3777;
  assign n6708 = n5374 & ~n6707;
  assign n6709 = n6708 ^ n3777;
  assign n6716 = n6715 ^ n6709;
  assign n6702 = n6611 ^ n3413;
  assign n6703 = n6611 ^ n6599;
  assign n6704 = ~n6702 & ~n6703;
  assign n6705 = n6704 ^ n3413;
  assign n6706 = n6705 ^ n3327;
  assign n6717 = n6716 ^ n6706;
  assign n6719 = n6718 ^ n6717;
  assign n6613 = n6612 ^ n6595;
  assign n6614 = n6613 ^ x226;
  assign n6615 = n6594 ^ n6577;
  assign n6616 = n6615 ^ x227;
  assign n6617 = n6576 ^ n6540;
  assign n6618 = n6617 ^ x228;
  assign n6619 = n6575 ^ n6573;
  assign n6620 = n6619 ^ x229;
  assign n6621 = n6572 ^ n6571;
  assign n6622 = n6621 ^ x230;
  assign n6623 = n6570 ^ n6569;
  assign n6624 = n6623 ^ x231;
  assign n6625 = n6568 ^ n6567;
  assign n6626 = n6625 ^ x232;
  assign n6627 = n6566 ^ n6564;
  assign n6628 = n6627 ^ x233;
  assign n6629 = n6563 ^ n6562;
  assign n6630 = n6629 ^ x234;
  assign n6631 = n6561 ^ n6559;
  assign n6632 = n6631 ^ x235;
  assign n6633 = n6558 ^ n6557;
  assign n6634 = n6633 ^ x236;
  assign n6635 = n6556 ^ n6542;
  assign n6636 = n6635 ^ x237;
  assign n6637 = n6555 ^ n6543;
  assign n6638 = n6637 ^ x238;
  assign n6657 = n6554 ^ n6553;
  assign n6639 = n6552 ^ n6550;
  assign n6640 = n6639 ^ x240;
  assign n6641 = n6549 ^ n6545;
  assign n6642 = n6641 ^ x241;
  assign n6643 = n6548 ^ n6547;
  assign n6644 = n6643 ^ x242;
  assign n6265 = n6264 ^ n6248;
  assign n6266 = n6265 ^ x243;
  assign n6192 = n6191 ^ n6165;
  assign n6193 = n6192 ^ x244;
  assign n6194 = n6190 ^ n6167;
  assign n6195 = n6194 ^ x245;
  assign n6196 = n6189 ^ n6188;
  assign n6197 = n6196 ^ x246;
  assign n6198 = n6187 ^ n6185;
  assign n6199 = n6198 ^ x247;
  assign n6201 = n6200 ^ x248;
  assign n6233 = n6232 ^ n6200;
  assign n6234 = n6201 & ~n6233;
  assign n6235 = n6234 ^ x248;
  assign n6236 = n6235 ^ n6198;
  assign n6237 = ~n6199 & n6236;
  assign n6238 = n6237 ^ x247;
  assign n6239 = n6238 ^ n6196;
  assign n6240 = n6197 & ~n6239;
  assign n6241 = n6240 ^ x246;
  assign n6242 = n6241 ^ n6194;
  assign n6243 = n6195 & ~n6242;
  assign n6244 = n6243 ^ x245;
  assign n6245 = n6244 ^ n6192;
  assign n6246 = n6193 & ~n6245;
  assign n6247 = n6246 ^ x244;
  assign n6645 = n6265 ^ n6247;
  assign n6646 = n6266 & ~n6645;
  assign n6647 = n6646 ^ x243;
  assign n6648 = n6647 ^ n6643;
  assign n6649 = n6644 & ~n6648;
  assign n6650 = n6649 ^ x242;
  assign n6651 = n6650 ^ n6641;
  assign n6652 = ~n6642 & n6651;
  assign n6653 = n6652 ^ x241;
  assign n6654 = n6653 ^ n6639;
  assign n6655 = ~n6640 & n6654;
  assign n6656 = n6655 ^ x240;
  assign n6658 = n6657 ^ n6656;
  assign n6659 = n6657 ^ x239;
  assign n6660 = ~n6658 & n6659;
  assign n6661 = n6660 ^ x239;
  assign n6662 = n6661 ^ n6637;
  assign n6663 = ~n6638 & n6662;
  assign n6664 = n6663 ^ x238;
  assign n6665 = n6664 ^ n6635;
  assign n6666 = n6636 & ~n6665;
  assign n6667 = n6666 ^ x237;
  assign n6668 = n6667 ^ n6633;
  assign n6669 = n6634 & ~n6668;
  assign n6670 = n6669 ^ x236;
  assign n6671 = n6670 ^ n6631;
  assign n6672 = n6632 & ~n6671;
  assign n6673 = n6672 ^ x235;
  assign n6674 = n6673 ^ n6629;
  assign n6675 = ~n6630 & n6674;
  assign n6676 = n6675 ^ x234;
  assign n6677 = n6676 ^ n6627;
  assign n6678 = n6628 & ~n6677;
  assign n6679 = n6678 ^ x233;
  assign n6680 = n6679 ^ n6625;
  assign n6681 = ~n6626 & n6680;
  assign n6682 = n6681 ^ x232;
  assign n6683 = n6682 ^ n6623;
  assign n6684 = ~n6624 & n6683;
  assign n6685 = n6684 ^ x231;
  assign n6686 = n6685 ^ n6621;
  assign n6687 = ~n6622 & n6686;
  assign n6688 = n6687 ^ x230;
  assign n6689 = n6688 ^ n6619;
  assign n6690 = n6620 & ~n6689;
  assign n6691 = n6690 ^ x229;
  assign n6692 = n6691 ^ n6617;
  assign n6693 = n6618 & ~n6692;
  assign n6694 = n6693 ^ x228;
  assign n6695 = n6694 ^ n6615;
  assign n6696 = n6616 & ~n6695;
  assign n6697 = n6696 ^ x227;
  assign n6698 = n6697 ^ n6613;
  assign n6699 = n6614 & ~n6698;
  assign n6700 = n6699 ^ x226;
  assign n6701 = n6700 ^ x225;
  assign n6720 = n6719 ^ n6701;
  assign n6724 = n6723 ^ n6720;
  assign n6728 = n6697 ^ x226;
  assign n6729 = n6728 ^ n6613;
  assign n6725 = n4623 ^ n4588;
  assign n6726 = ~n5726 & ~n6725;
  assign n6727 = n6726 ^ n4623;
  assign n6730 = n6729 ^ n6727;
  assign n6732 = n4694 ^ n4598;
  assign n6733 = n5731 & n6732;
  assign n6734 = n6733 ^ n4694;
  assign n6731 = n6694 ^ n6616;
  assign n6735 = n6734 ^ n6731;
  assign n6736 = n4667 ^ n4609;
  assign n6737 = n5739 & ~n6736;
  assign n6738 = n6737 ^ n4667;
  assign n6739 = n6691 ^ x228;
  assign n6740 = n6739 ^ n6617;
  assign n6741 = n6738 & n6740;
  assign n6742 = n6741 ^ n6731;
  assign n6743 = ~n6735 & n6742;
  assign n6744 = n6743 ^ n6741;
  assign n6745 = n6744 ^ n6729;
  assign n6746 = ~n6730 & ~n6745;
  assign n6747 = n6746 ^ n6727;
  assign n6748 = n6747 ^ n6720;
  assign n6749 = n6724 & n6748;
  assign n6750 = n6749 ^ n6723;
  assign n6754 = n6753 ^ n6750;
  assign n6771 = n5975 ^ n5931;
  assign n6768 = n4672 ^ n3772;
  assign n6769 = n5371 & n6768;
  assign n6770 = n6769 ^ n3772;
  assign n6772 = n6771 ^ n6770;
  assign n6773 = n6772 ^ n3323;
  assign n6765 = n6714 ^ n6709;
  assign n6766 = n6715 & n6765;
  assign n6767 = n6766 ^ n6709;
  assign n6774 = n6773 ^ n6767;
  assign n6764 = n6717 & ~n6718;
  assign n6775 = n6774 ^ n6764;
  assign n6760 = n6716 ^ n3327;
  assign n6761 = n6716 ^ n6705;
  assign n6762 = n6760 & n6761;
  assign n6763 = n6762 ^ n3327;
  assign n6776 = n6775 ^ n6763;
  assign n6755 = n6719 ^ x225;
  assign n6756 = n6719 ^ n6700;
  assign n6757 = n6755 & ~n6756;
  assign n6758 = n6757 ^ x225;
  assign n6759 = n6758 ^ x224;
  assign n6777 = n6776 ^ n6759;
  assign n6778 = n6777 ^ n6750;
  assign n6779 = n6754 & n6778;
  assign n6780 = n6779 ^ n6753;
  assign n6781 = n6780 ^ n6342;
  assign n6782 = ~n6346 & ~n6781;
  assign n6783 = n6782 ^ n6345;
  assign n6784 = n6783 ^ n6340;
  assign n6785 = n6341 & n6784;
  assign n6786 = n6785 ^ n6339;
  assign n6787 = n6786 ^ n6335;
  assign n6788 = ~n6336 & n6787;
  assign n6789 = n6788 ^ n6334;
  assign n6790 = n6789 ^ n6330;
  assign n6791 = ~n6331 & n6790;
  assign n6792 = n6791 ^ n6328;
  assign n6793 = n6792 ^ n6318;
  assign n6794 = ~n6323 & ~n6793;
  assign n6795 = n6794 ^ n6322;
  assign n6796 = n6795 ^ n6316;
  assign n6797 = ~n6317 & n6796;
  assign n6798 = n6797 ^ n6314;
  assign n6799 = n6798 ^ n6304;
  assign n6800 = n6310 & ~n6799;
  assign n6801 = n6800 ^ n6309;
  assign n6802 = n6801 ^ n6302;
  assign n6803 = n6303 & n6802;
  assign n6804 = n6803 ^ n6300;
  assign n6293 = n5779 ^ n4766;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = n6294 ^ n4766;
  assign n6838 = n6804 ^ n6295;
  assign n6289 = n6235 ^ x247;
  assign n6290 = n6289 ^ n6198;
  assign n6839 = n6838 ^ n6290;
  assign n6840 = n6839 ^ n3692;
  assign n6841 = n6801 ^ n6303;
  assign n6842 = n6841 ^ n3698;
  assign n6843 = n6798 ^ n6309;
  assign n6844 = n6843 ^ n6304;
  assign n6845 = n6844 ^ n3708;
  assign n6846 = n6795 ^ n6317;
  assign n6847 = n6846 ^ n3711;
  assign n6848 = n6792 ^ n6322;
  assign n6849 = n6848 ^ n6318;
  assign n6850 = n6849 ^ n3722;
  assign n6851 = n6789 ^ n6331;
  assign n6852 = n6851 ^ n3732;
  assign n6853 = n6786 ^ n6334;
  assign n6854 = n6853 ^ n6335;
  assign n6855 = n6854 ^ n3737;
  assign n6856 = n6783 ^ n6341;
  assign n6857 = n6856 ^ n3742;
  assign n6858 = n6780 ^ n6346;
  assign n6859 = n6858 ^ n3750;
  assign n6860 = n6777 ^ n6753;
  assign n6861 = n6860 ^ n6750;
  assign n6862 = n6861 ^ n4041;
  assign n6863 = n6747 ^ n6723;
  assign n6864 = n6863 ^ n6720;
  assign n6865 = n6864 ^ n3758;
  assign n6866 = n6744 ^ n6730;
  assign n6867 = n6866 ^ n4030;
  assign n6868 = n6740 ^ n6738;
  assign n6869 = ~n3770 & n6868;
  assign n6870 = n6869 ^ n3761;
  assign n6871 = n6741 ^ n6734;
  assign n6872 = n6871 ^ n6731;
  assign n6873 = n6872 ^ n6869;
  assign n6874 = n6870 & ~n6873;
  assign n6875 = n6874 ^ n3761;
  assign n6876 = n6875 ^ n6866;
  assign n6877 = ~n6867 & n6876;
  assign n6878 = n6877 ^ n4030;
  assign n6879 = n6878 ^ n6864;
  assign n6880 = ~n6865 & n6879;
  assign n6881 = n6880 ^ n3758;
  assign n6882 = n6881 ^ n6861;
  assign n6883 = ~n6862 & n6882;
  assign n6884 = n6883 ^ n4041;
  assign n6885 = n6884 ^ n6858;
  assign n6886 = ~n6859 & n6885;
  assign n6887 = n6886 ^ n3750;
  assign n6888 = n6887 ^ n6856;
  assign n6889 = ~n6857 & n6888;
  assign n6890 = n6889 ^ n3742;
  assign n6891 = n6890 ^ n6854;
  assign n6892 = ~n6855 & n6891;
  assign n6893 = n6892 ^ n3737;
  assign n6894 = n6893 ^ n6851;
  assign n6895 = n6852 & n6894;
  assign n6896 = n6895 ^ n3732;
  assign n6897 = n6896 ^ n6849;
  assign n6898 = n6850 & ~n6897;
  assign n6899 = n6898 ^ n3722;
  assign n6900 = n6899 ^ n6846;
  assign n6901 = n6847 & n6900;
  assign n6902 = n6901 ^ n3711;
  assign n6903 = n6902 ^ n6844;
  assign n6904 = n6845 & n6903;
  assign n6905 = n6904 ^ n3708;
  assign n6906 = n6905 ^ n6841;
  assign n6907 = ~n6842 & ~n6906;
  assign n6908 = n6907 ^ n3698;
  assign n6909 = n6908 ^ n6839;
  assign n6910 = ~n6840 & n6909;
  assign n6911 = n6910 ^ n3692;
  assign n6973 = n6911 ^ n3686;
  assign n6296 = n6295 ^ n6290;
  assign n6805 = n6804 ^ n6290;
  assign n6806 = ~n6296 & n6805;
  assign n6807 = n6806 ^ n6295;
  assign n6287 = n6238 ^ n6197;
  assign n6284 = n5787 ^ n4775;
  assign n6285 = n6283 & n6284;
  assign n6286 = n6285 ^ n4775;
  assign n6288 = n6287 ^ n6286;
  assign n6836 = n6807 ^ n6288;
  assign n6974 = n6973 ^ n6836;
  assign n6940 = n6893 ^ n3732;
  assign n6941 = n6940 ^ n6851;
  assign n6942 = n6887 ^ n3742;
  assign n6943 = n6942 ^ n6856;
  assign n6944 = n6875 ^ n4030;
  assign n6945 = n6944 ^ n6866;
  assign n6946 = n6872 ^ n6870;
  assign n6947 = n6868 ^ n3770;
  assign n6948 = n6946 & ~n6947;
  assign n6949 = ~n6945 & n6948;
  assign n6950 = n6878 ^ n6865;
  assign n6951 = ~n6949 & n6950;
  assign n6952 = n6881 ^ n4041;
  assign n6953 = n6952 ^ n6861;
  assign n6954 = n6951 & n6953;
  assign n6955 = n6884 ^ n6859;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~n6943 & n6956;
  assign n6958 = n6890 ^ n6855;
  assign n6959 = ~n6957 & n6958;
  assign n6960 = ~n6941 & n6959;
  assign n6961 = n6896 ^ n6850;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = n6899 ^ n3711;
  assign n6964 = n6963 ^ n6846;
  assign n6965 = n6962 & ~n6964;
  assign n6966 = n6902 ^ n6845;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = n6905 ^ n3698;
  assign n6969 = n6968 ^ n6841;
  assign n6970 = n6967 & ~n6969;
  assign n6971 = n6908 ^ n6840;
  assign n6972 = n6970 & n6971;
  assign n7121 = n6974 ^ n6972;
  assign n7122 = n7121 ^ x273;
  assign n7123 = n6971 ^ n6970;
  assign n7124 = n7123 ^ x274;
  assign n7125 = n6969 ^ n6967;
  assign n7126 = n7125 ^ x275;
  assign n7127 = n6966 ^ n6965;
  assign n7128 = n7127 ^ x276;
  assign n7129 = n6964 ^ n6962;
  assign n7130 = n7129 ^ x277;
  assign n7131 = n6961 ^ n6960;
  assign n7132 = n7131 ^ x278;
  assign n7133 = n6959 ^ n6941;
  assign n7134 = n7133 ^ x279;
  assign n7135 = n6958 ^ n6957;
  assign n7136 = n7135 ^ x280;
  assign n7137 = n6956 ^ n6943;
  assign n7138 = n7137 ^ x281;
  assign n7139 = n6955 ^ n6954;
  assign n7140 = n7139 ^ x282;
  assign n7141 = n6953 ^ n6951;
  assign n7142 = n7141 ^ x283;
  assign n7143 = n6950 ^ n6949;
  assign n7144 = n7143 ^ x284;
  assign n7145 = n6948 ^ n6945;
  assign n7146 = n7145 ^ x285;
  assign n7147 = x287 & n6947;
  assign n7148 = n7147 ^ x286;
  assign n7149 = n6947 ^ n6946;
  assign n7150 = n7149 ^ n7147;
  assign n7151 = n7148 & n7150;
  assign n7152 = n7151 ^ x286;
  assign n7153 = n7152 ^ n7145;
  assign n7154 = ~n7146 & n7153;
  assign n7155 = n7154 ^ x285;
  assign n7156 = n7155 ^ n7143;
  assign n7157 = n7144 & ~n7156;
  assign n7158 = n7157 ^ x284;
  assign n7159 = n7158 ^ n7141;
  assign n7160 = ~n7142 & n7159;
  assign n7161 = n7160 ^ x283;
  assign n7162 = n7161 ^ n7139;
  assign n7163 = n7140 & ~n7162;
  assign n7164 = n7163 ^ x282;
  assign n7165 = n7164 ^ n7137;
  assign n7166 = ~n7138 & n7165;
  assign n7167 = n7166 ^ x281;
  assign n7168 = n7167 ^ n7135;
  assign n7169 = n7136 & ~n7168;
  assign n7170 = n7169 ^ x280;
  assign n7171 = n7170 ^ n7133;
  assign n7172 = n7134 & ~n7171;
  assign n7173 = n7172 ^ x279;
  assign n7174 = n7173 ^ n7131;
  assign n7175 = n7132 & ~n7174;
  assign n7176 = n7175 ^ x278;
  assign n7177 = n7176 ^ n7129;
  assign n7178 = ~n7130 & n7177;
  assign n7179 = n7178 ^ x277;
  assign n7180 = n7179 ^ n7127;
  assign n7181 = ~n7128 & n7180;
  assign n7182 = n7181 ^ x276;
  assign n7183 = n7182 ^ n7125;
  assign n7184 = n7126 & ~n7183;
  assign n7185 = n7184 ^ x275;
  assign n7186 = n7185 ^ n7123;
  assign n7187 = ~n7124 & n7186;
  assign n7188 = n7187 ^ x274;
  assign n7189 = n7188 ^ n7121;
  assign n7190 = n7122 & ~n7189;
  assign n7191 = n7190 ^ x273;
  assign n7755 = n7191 ^ x272;
  assign n6837 = n6836 ^ n3686;
  assign n6912 = n6911 ^ n6836;
  assign n6913 = n6837 & n6912;
  assign n6914 = n6913 ^ n3686;
  assign n6808 = n6807 ^ n6287;
  assign n6809 = ~n6288 & ~n6808;
  assign n6810 = n6809 ^ n6286;
  assign n6278 = n5795 ^ n4779;
  assign n6279 = n6277 & n6278;
  assign n6280 = n6279 ^ n4779;
  assign n6833 = n6810 ^ n6280;
  assign n6281 = n6241 ^ n6195;
  assign n6834 = n6833 ^ n6281;
  assign n6835 = n6834 ^ n4083;
  assign n6976 = n6914 ^ n6835;
  assign n6975 = n6972 & ~n6974;
  assign n7119 = n6976 ^ n6975;
  assign n7756 = n7755 ^ n7119;
  assign n7027 = n6661 ^ x238;
  assign n7028 = n7027 ^ n6637;
  assign n7839 = n7028 ^ n5710;
  assign n7840 = ~n7756 & n7839;
  assign n7841 = n7840 ^ n5710;
  assign n7347 = n6319 ^ n5569;
  assign n7348 = n6302 & ~n7347;
  assign n7349 = n7348 ^ n5569;
  assign n7346 = n7152 ^ n7146;
  assign n7350 = n7349 ^ n7346;
  assign n7454 = n7149 ^ n7148;
  assign n7352 = n6262 ^ n5534;
  assign n7353 = n6316 & ~n7352;
  assign n7354 = n7353 ^ n5534;
  assign n7351 = n6947 ^ x287;
  assign n7355 = n7354 ^ n7351;
  assign n7421 = n6162 ^ n5494;
  assign n7422 = n6318 & ~n7421;
  assign n7423 = n7422 ^ n5494;
  assign n7371 = n6682 ^ n6624;
  assign n7277 = n6679 ^ x232;
  assign n7278 = n7277 ^ n6625;
  assign n7273 = n5374 ^ n4520;
  assign n7274 = ~n6059 & n7273;
  assign n7275 = n7274 ^ n4520;
  assign n7367 = n7278 ^ n7275;
  assign n7245 = n6676 ^ n6628;
  assign n7241 = n5383 ^ n4480;
  assign n7242 = ~n6064 & ~n7241;
  assign n7243 = n7242 ^ n4480;
  assign n7269 = n7245 ^ n7243;
  assign n7095 = n6673 ^ x234;
  assign n7096 = n7095 ^ n6629;
  assign n7091 = n5391 ^ n4445;
  assign n7092 = n6771 & ~n7091;
  assign n7093 = n7092 ^ n4445;
  assign n7237 = n7096 ^ n7093;
  assign n7078 = n6670 ^ n6632;
  assign n7074 = n5394 ^ n4411;
  assign n7075 = ~n6714 & n7074;
  assign n7076 = n7075 ^ n4411;
  assign n7087 = n7078 ^ n7076;
  assign n7060 = n6667 ^ x236;
  assign n7061 = n7060 ^ n6633;
  assign n7057 = n6040 ^ n5364;
  assign n7058 = n6609 & ~n7057;
  assign n7059 = n7058 ^ n5364;
  assign n7062 = n7061 ^ n7059;
  assign n7045 = n6664 ^ n6636;
  assign n7041 = n6017 ^ n5066;
  assign n7042 = n6592 & n7041;
  assign n7043 = n7042 ^ n5066;
  assign n7053 = n7045 ^ n7043;
  assign n7011 = n6658 ^ x239;
  assign n6995 = n6653 ^ x240;
  assign n6996 = n6995 ^ n6639;
  assign n6992 = n5824 ^ n4845;
  assign n6993 = ~n6347 & n6992;
  assign n6994 = n6993 ^ n4845;
  assign n6997 = n6996 ^ n6994;
  assign n6933 = n6650 ^ n6642;
  assign n6930 = n5744 ^ n4830;
  assign n6931 = ~n6353 & n6930;
  assign n6932 = n6931 ^ n4830;
  assign n6934 = n6933 ^ n6932;
  assign n6823 = n6647 ^ x242;
  assign n6824 = n6823 ^ n6643;
  assign n6820 = n5750 ^ n4840;
  assign n6821 = ~n6358 & ~n6820;
  assign n6822 = n6821 ^ n4840;
  assign n6825 = n6824 ^ n6822;
  assign n6267 = n6266 ^ n6247;
  assign n5712 = n5711 ^ n4838;
  assign n5713 = ~n5710 & n5712;
  assign n5714 = n5713 ^ n4838;
  assign n6268 = n6267 ^ n5714;
  assign n6273 = n6244 ^ x244;
  assign n6274 = n6273 ^ n6192;
  assign n6270 = n5755 ^ n4786;
  assign n6271 = n6269 & n6270;
  assign n6272 = n6271 ^ n4786;
  assign n6275 = n6274 ^ n6272;
  assign n6282 = n6281 ^ n6280;
  assign n6811 = n6810 ^ n6281;
  assign n6812 = n6282 & n6811;
  assign n6813 = n6812 ^ n6280;
  assign n6814 = n6813 ^ n6274;
  assign n6815 = ~n6275 & ~n6814;
  assign n6816 = n6815 ^ n6272;
  assign n6817 = n6816 ^ n6267;
  assign n6818 = ~n6268 & n6817;
  assign n6819 = n6818 ^ n5714;
  assign n6927 = n6824 ^ n6819;
  assign n6928 = ~n6825 & n6927;
  assign n6929 = n6928 ^ n6822;
  assign n6989 = n6933 ^ n6929;
  assign n6990 = ~n6934 & ~n6989;
  assign n6991 = n6990 ^ n6932;
  assign n7008 = n6996 ^ n6991;
  assign n7009 = n6997 & n7008;
  assign n7010 = n7009 ^ n6994;
  assign n7012 = n7011 ^ n7010;
  assign n7005 = n5886 ^ n4638;
  assign n7006 = ~n6451 & ~n7005;
  assign n7007 = n7006 ^ n4638;
  assign n7024 = n7011 ^ n7007;
  assign n7025 = n7012 & n7024;
  assign n7026 = n7025 ^ n7007;
  assign n7029 = n7028 ^ n7026;
  assign n7021 = n5996 ^ n4876;
  assign n7022 = ~n6538 & n7021;
  assign n7023 = n7022 ^ n4876;
  assign n7038 = n7028 ^ n7023;
  assign n7039 = n7029 & ~n7038;
  assign n7040 = n7039 ^ n7023;
  assign n7054 = n7045 ^ n7040;
  assign n7055 = n7053 & ~n7054;
  assign n7056 = n7055 ^ n7043;
  assign n7071 = n7061 ^ n7056;
  assign n7072 = n7062 & ~n7071;
  assign n7073 = n7072 ^ n7059;
  assign n7088 = n7078 ^ n7073;
  assign n7089 = n7087 & ~n7088;
  assign n7090 = n7089 ^ n7076;
  assign n7238 = n7096 ^ n7090;
  assign n7239 = ~n7237 & n7238;
  assign n7240 = n7239 ^ n7093;
  assign n7270 = n7245 ^ n7240;
  assign n7271 = n7269 & ~n7270;
  assign n7272 = n7271 ^ n7243;
  assign n7368 = n7278 ^ n7272;
  assign n7369 = ~n7367 & n7368;
  assign n7370 = n7369 ^ n7275;
  assign n7372 = n7371 ^ n7370;
  assign n7364 = n5371 ^ n4565;
  assign n7365 = ~n6057 & n7364;
  assign n7366 = n7365 ^ n4565;
  assign n7373 = n7372 ^ n7366;
  assign n7276 = n7275 ^ n7272;
  assign n7279 = n7278 ^ n7276;
  assign n7359 = n7279 ^ n3987;
  assign n7244 = n7243 ^ n7240;
  assign n7246 = n7245 ^ n7244;
  assign n7264 = n7246 ^ n4007;
  assign n7094 = n7093 ^ n7090;
  assign n7097 = n7096 ^ n7094;
  assign n7232 = n7097 ^ n3990;
  assign n7077 = n7076 ^ n7073;
  assign n7079 = n7078 ^ n7077;
  assign n7082 = n7079 ^ n3998;
  assign n7063 = n7062 ^ n7056;
  assign n7064 = n7063 ^ n4554;
  assign n7044 = n7043 ^ n7040;
  assign n7046 = n7045 ^ n7044;
  assign n7049 = n7046 ^ n4506;
  assign n7030 = n7029 ^ n7023;
  assign n7033 = n7030 ^ n4470;
  assign n7013 = n7012 ^ n7007;
  assign n7014 = n7013 ^ n4438;
  assign n6998 = n6997 ^ n6991;
  assign n7001 = n6998 ^ n4404;
  assign n6935 = n6934 ^ n6929;
  assign n6936 = n6935 ^ n4115;
  assign n6826 = n6825 ^ n6819;
  assign n6827 = n6826 ^ n4100;
  assign n6828 = n6816 ^ n5714;
  assign n6829 = n6828 ^ n6267;
  assign n6830 = n6829 ^ n3673;
  assign n6831 = n6813 ^ n6275;
  assign n6832 = n6831 ^ n3679;
  assign n6915 = n6914 ^ n6834;
  assign n6916 = ~n6835 & ~n6915;
  assign n6917 = n6916 ^ n4083;
  assign n6918 = n6917 ^ n6831;
  assign n6919 = n6832 & n6918;
  assign n6920 = n6919 ^ n3679;
  assign n6921 = n6920 ^ n6829;
  assign n6922 = ~n6830 & n6921;
  assign n6923 = n6922 ^ n3673;
  assign n6924 = n6923 ^ n6826;
  assign n6925 = n6827 & n6924;
  assign n6926 = n6925 ^ n4100;
  assign n6985 = n6935 ^ n6926;
  assign n6986 = n6936 & ~n6985;
  assign n6987 = n6986 ^ n4115;
  assign n7002 = n6998 ^ n6987;
  assign n7003 = n7001 & ~n7002;
  assign n7004 = n7003 ^ n4404;
  assign n7017 = n7013 ^ n7004;
  assign n7018 = ~n7014 & n7017;
  assign n7019 = n7018 ^ n4438;
  assign n7034 = n7030 ^ n7019;
  assign n7035 = ~n7033 & n7034;
  assign n7036 = n7035 ^ n4470;
  assign n7050 = n7046 ^ n7036;
  assign n7051 = ~n7049 & ~n7050;
  assign n7052 = n7051 ^ n4506;
  assign n7067 = n7063 ^ n7052;
  assign n7068 = n7064 & n7067;
  assign n7069 = n7068 ^ n4554;
  assign n7083 = n7079 ^ n7069;
  assign n7084 = n7082 & ~n7083;
  assign n7085 = n7084 ^ n3998;
  assign n7233 = n7097 ^ n7085;
  assign n7234 = ~n7232 & n7233;
  assign n7235 = n7234 ^ n3990;
  assign n7265 = n7246 ^ n7235;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = n7266 ^ n4007;
  assign n7360 = n7279 ^ n7267;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = n7361 ^ n3987;
  assign n7363 = n7362 ^ n3977;
  assign n7374 = n7373 ^ n7363;
  assign n6937 = n6936 ^ n6926;
  assign n6938 = n6923 ^ n4100;
  assign n6939 = n6938 ^ n6826;
  assign n6977 = ~n6975 & n6976;
  assign n6978 = n6917 ^ n6832;
  assign n6979 = n6977 & n6978;
  assign n6980 = n6920 ^ n3673;
  assign n6981 = n6980 ^ n6829;
  assign n6982 = ~n6979 & ~n6981;
  assign n6983 = ~n6939 & ~n6982;
  assign n6984 = n6937 & n6983;
  assign n6988 = n6987 ^ n4404;
  assign n6999 = n6998 ^ n6988;
  assign n7000 = n6984 & n6999;
  assign n7015 = n7014 ^ n7004;
  assign n7016 = n7000 & ~n7015;
  assign n7020 = n7019 ^ n4470;
  assign n7031 = n7030 ^ n7020;
  assign n7032 = n7016 & ~n7031;
  assign n7037 = n7036 ^ n4506;
  assign n7047 = n7046 ^ n7037;
  assign n7048 = ~n7032 & n7047;
  assign n7065 = n7064 ^ n7052;
  assign n7066 = ~n7048 & ~n7065;
  assign n7070 = n7069 ^ n3998;
  assign n7080 = n7079 ^ n7070;
  assign n7081 = ~n7066 & ~n7080;
  assign n7086 = n7085 ^ n3990;
  assign n7098 = n7097 ^ n7086;
  assign n7231 = ~n7081 & ~n7098;
  assign n7236 = n7235 ^ n4007;
  assign n7247 = n7246 ^ n7236;
  assign n7263 = ~n7231 & n7247;
  assign n7268 = n7267 ^ n3987;
  assign n7280 = n7279 ^ n7268;
  assign n7375 = n7263 & ~n7280;
  assign n7402 = ~n7374 & ~n7375;
  assign n7397 = n6685 ^ x230;
  assign n7398 = n7397 ^ n6621;
  assign n7394 = n7371 ^ n7366;
  assign n7395 = n7372 & ~n7394;
  assign n7396 = n7395 ^ n7366;
  assign n7399 = n7398 ^ n7396;
  assign n7391 = n4680 ^ n4617;
  assign n7392 = ~n6052 & n7391;
  assign n7393 = n7392 ^ n4680;
  assign n7400 = n7399 ^ n7393;
  assign n7386 = n7373 ^ n3977;
  assign n7387 = n7373 ^ n7362;
  assign n7388 = ~n7386 & n7387;
  assign n7389 = n7388 ^ n3977;
  assign n7390 = n7389 ^ n3777;
  assign n7401 = n7400 ^ n7390;
  assign n7403 = n7402 ^ n7401;
  assign n7376 = n7375 ^ n7374;
  assign n7377 = n7376 ^ x258;
  assign n7281 = n7280 ^ n7263;
  assign n7378 = n7281 ^ x259;
  assign n7248 = n7247 ^ n7231;
  assign n7258 = n7248 ^ x260;
  assign n7099 = n7098 ^ n7081;
  assign n7100 = n7099 ^ x261;
  assign n7101 = n7080 ^ n7066;
  assign n7102 = n7101 ^ x262;
  assign n7103 = n7065 ^ n7048;
  assign n7104 = n7103 ^ x263;
  assign n7105 = n7047 ^ n7032;
  assign n7106 = n7105 ^ x264;
  assign n7107 = n7031 ^ n7016;
  assign n7108 = n7107 ^ x265;
  assign n7109 = n7015 ^ n7000;
  assign n7110 = n7109 ^ x266;
  assign n7111 = n6999 ^ n6984;
  assign n7112 = n7111 ^ x267;
  assign n7113 = n6983 ^ n6937;
  assign n7114 = n7113 ^ x268;
  assign n7115 = n6982 ^ n6939;
  assign n7116 = n7115 ^ x269;
  assign n7117 = n6981 ^ n6979;
  assign n7118 = n7117 ^ x270;
  assign n7195 = n6978 ^ n6977;
  assign n7120 = n7119 ^ x272;
  assign n7192 = n7191 ^ n7119;
  assign n7193 = ~n7120 & n7192;
  assign n7194 = n7193 ^ x272;
  assign n7196 = n7195 ^ n7194;
  assign n7197 = n7195 ^ x271;
  assign n7198 = ~n7196 & n7197;
  assign n7199 = n7198 ^ x271;
  assign n7200 = n7199 ^ n7117;
  assign n7201 = ~n7118 & n7200;
  assign n7202 = n7201 ^ x270;
  assign n7203 = n7202 ^ n7115;
  assign n7204 = n7116 & ~n7203;
  assign n7205 = n7204 ^ x269;
  assign n7206 = n7205 ^ n7113;
  assign n7207 = n7114 & ~n7206;
  assign n7208 = n7207 ^ x268;
  assign n7209 = n7208 ^ n7111;
  assign n7210 = n7112 & ~n7209;
  assign n7211 = n7210 ^ x267;
  assign n7212 = n7211 ^ n7109;
  assign n7213 = ~n7110 & n7212;
  assign n7214 = n7213 ^ x266;
  assign n7215 = n7214 ^ n7107;
  assign n7216 = ~n7108 & n7215;
  assign n7217 = n7216 ^ x265;
  assign n7218 = n7217 ^ n7105;
  assign n7219 = n7106 & ~n7218;
  assign n7220 = n7219 ^ x264;
  assign n7221 = n7220 ^ n7103;
  assign n7222 = n7104 & ~n7221;
  assign n7223 = n7222 ^ x263;
  assign n7224 = n7223 ^ n7101;
  assign n7225 = ~n7102 & n7224;
  assign n7226 = n7225 ^ x262;
  assign n7227 = n7226 ^ n7099;
  assign n7228 = n7100 & ~n7227;
  assign n7229 = n7228 ^ x261;
  assign n7259 = n7248 ^ n7229;
  assign n7260 = n7258 & ~n7259;
  assign n7261 = n7260 ^ x260;
  assign n7379 = n7281 ^ n7261;
  assign n7380 = n7378 & ~n7379;
  assign n7381 = n7380 ^ x259;
  assign n7382 = n7381 ^ n7376;
  assign n7383 = n7377 & ~n7382;
  assign n7384 = n7383 ^ x258;
  assign n7385 = n7384 ^ x257;
  assign n7404 = n7403 ^ n7385;
  assign n7356 = n6100 ^ n5431;
  assign n7357 = ~n6330 & n7356;
  assign n7358 = n7357 ^ n5431;
  assign n7405 = n7404 ^ n7358;
  assign n7410 = n5718 ^ n4588;
  assign n7411 = ~n6335 & n7410;
  assign n7412 = n7411 ^ n4588;
  assign n7262 = n7261 ^ x259;
  assign n7282 = n7281 ^ n7262;
  assign n7254 = n5724 ^ n4598;
  assign n7255 = n6340 & n7254;
  assign n7256 = n7255 ^ n4598;
  assign n7406 = n7282 ^ n7256;
  assign n7230 = n7229 ^ x260;
  assign n7249 = n7248 ^ n7230;
  assign n7250 = n5726 ^ n4609;
  assign n7251 = n6342 & n7250;
  assign n7252 = n7251 ^ n4609;
  assign n7253 = n7249 & ~n7252;
  assign n7407 = n7282 ^ n7253;
  assign n7408 = ~n7406 & n7407;
  assign n7409 = n7408 ^ n7253;
  assign n7413 = n7412 ^ n7409;
  assign n7414 = n7381 ^ n7377;
  assign n7415 = n7414 ^ n7409;
  assign n7416 = n7413 & ~n7415;
  assign n7417 = n7416 ^ n7412;
  assign n7418 = n7417 ^ n7404;
  assign n7419 = ~n7405 & n7418;
  assign n7420 = n7419 ^ n7358;
  assign n7424 = n7423 ^ n7420;
  assign n7441 = n6688 ^ n6620;
  assign n7438 = n4672 ^ n4611;
  assign n7439 = ~n6047 & n7438;
  assign n7440 = n7439 ^ n4672;
  assign n7442 = n7441 ^ n7440;
  assign n7443 = n7442 ^ n3772;
  assign n7435 = n7398 ^ n7393;
  assign n7436 = n7399 & ~n7435;
  assign n7437 = n7436 ^ n7393;
  assign n7444 = n7443 ^ n7437;
  assign n7434 = ~n7401 & ~n7402;
  assign n7445 = n7444 ^ n7434;
  assign n7430 = n7400 ^ n3777;
  assign n7431 = n7400 ^ n7389;
  assign n7432 = n7430 & n7431;
  assign n7433 = n7432 ^ n3777;
  assign n7446 = n7445 ^ n7433;
  assign n7425 = n7403 ^ x257;
  assign n7426 = n7403 ^ n7384;
  assign n7427 = ~n7425 & n7426;
  assign n7428 = n7427 ^ x257;
  assign n7429 = n7428 ^ x256;
  assign n7447 = n7446 ^ n7429;
  assign n7448 = n7447 ^ n7420;
  assign n7449 = ~n7424 & ~n7448;
  assign n7450 = n7449 ^ n7423;
  assign n7451 = n7450 ^ n7351;
  assign n7452 = ~n7355 & n7451;
  assign n7453 = n7452 ^ n7354;
  assign n7455 = n7454 ^ n7453;
  assign n7456 = n6325 ^ n5551;
  assign n7457 = ~n6304 & n7456;
  assign n7458 = n7457 ^ n5551;
  assign n7459 = n7458 ^ n7454;
  assign n7460 = ~n7455 & ~n7459;
  assign n7461 = n7460 ^ n7458;
  assign n7462 = n7461 ^ n7346;
  assign n7463 = n7350 & n7462;
  assign n7464 = n7463 ^ n7349;
  assign n7342 = n6311 ^ n5587;
  assign n7343 = ~n6290 & ~n7342;
  assign n7344 = n7343 ^ n5587;
  assign n7517 = n7464 ^ n7344;
  assign n7293 = n7155 ^ x284;
  assign n7294 = n7293 ^ n7143;
  assign n7518 = n7517 ^ n7294;
  assign n7519 = n7518 ^ n4645;
  assign n7520 = n7461 ^ n7349;
  assign n7521 = n7520 ^ n7346;
  assign n7522 = n7521 ^ n4593;
  assign n7523 = n7458 ^ n7455;
  assign n7524 = n7523 ^ n4599;
  assign n7525 = n7450 ^ n7354;
  assign n7526 = n7525 ^ n7351;
  assign n7527 = n7526 ^ n4604;
  assign n7528 = n7447 ^ n7424;
  assign n7529 = n7528 ^ n4612;
  assign n7530 = n7417 ^ n7358;
  assign n7531 = n7530 ^ n7404;
  assign n7532 = n7531 ^ n4618;
  assign n7533 = n7414 ^ n7413;
  assign n7534 = n7533 ^ n4623;
  assign n7284 = n7252 ^ n7249;
  assign n7285 = n4667 & ~n7284;
  assign n7286 = n7285 ^ n4694;
  assign n7257 = n7256 ^ n7253;
  assign n7283 = n7282 ^ n7257;
  assign n7535 = n7285 ^ n7283;
  assign n7536 = n7286 & ~n7535;
  assign n7537 = n7536 ^ n4694;
  assign n7538 = n7537 ^ n7533;
  assign n7539 = ~n7534 & ~n7538;
  assign n7540 = n7539 ^ n4623;
  assign n7541 = n7540 ^ n7531;
  assign n7542 = ~n7532 & ~n7541;
  assign n7543 = n7542 ^ n4618;
  assign n7544 = n7543 ^ n7528;
  assign n7545 = ~n7529 & n7544;
  assign n7546 = n7545 ^ n4612;
  assign n7547 = n7546 ^ n7526;
  assign n7548 = ~n7527 & ~n7547;
  assign n7549 = n7548 ^ n4604;
  assign n7550 = n7549 ^ n7523;
  assign n7551 = n7524 & n7550;
  assign n7552 = n7551 ^ n4599;
  assign n7553 = n7552 ^ n7521;
  assign n7554 = n7522 & ~n7553;
  assign n7555 = n7554 ^ n4593;
  assign n7556 = n7555 ^ n7518;
  assign n7557 = n7519 & ~n7556;
  assign n7558 = n7557 ^ n4645;
  assign n7619 = n7558 ^ n4750;
  assign n7345 = n7344 ^ n7294;
  assign n7465 = n7464 ^ n7294;
  assign n7466 = ~n7345 & n7465;
  assign n7467 = n7466 ^ n7344;
  assign n7338 = n6306 ^ n5682;
  assign n7339 = n6287 & ~n7338;
  assign n7340 = n7339 ^ n5682;
  assign n7514 = n7467 ^ n7340;
  assign n7337 = n7158 ^ n7142;
  assign n7515 = n7514 ^ n7337;
  assign n7620 = n7619 ^ n7515;
  assign n7598 = n7555 ^ n4645;
  assign n7599 = n7598 ^ n7518;
  assign n7600 = n7552 ^ n4593;
  assign n7601 = n7600 ^ n7521;
  assign n7602 = n7540 ^ n7532;
  assign n7287 = n7286 ^ n7283;
  assign n7288 = n7284 ^ n4667;
  assign n7603 = n7287 & ~n7288;
  assign n7604 = n7537 ^ n4623;
  assign n7605 = n7604 ^ n7533;
  assign n7606 = n7603 & ~n7605;
  assign n7607 = ~n7602 & ~n7606;
  assign n7608 = n7543 ^ n4612;
  assign n7609 = n7608 ^ n7528;
  assign n7610 = n7607 & n7609;
  assign n7611 = n7546 ^ n4604;
  assign n7612 = n7611 ^ n7526;
  assign n7613 = ~n7610 & ~n7612;
  assign n7614 = n7549 ^ n4599;
  assign n7615 = n7614 ^ n7523;
  assign n7616 = n7613 & ~n7615;
  assign n7617 = ~n7601 & ~n7616;
  assign n7618 = ~n7599 & n7617;
  assign n7674 = n7620 ^ n7618;
  assign n7675 = n7674 ^ x310;
  assign n7676 = n7617 ^ n7599;
  assign n7677 = n7676 ^ x311;
  assign n7678 = n7616 ^ n7601;
  assign n7679 = n7678 ^ x312;
  assign n7680 = n7615 ^ n7613;
  assign n7681 = n7680 ^ x313;
  assign n7682 = n7612 ^ n7610;
  assign n7683 = n7682 ^ x314;
  assign n7684 = n7609 ^ n7607;
  assign n7685 = n7684 ^ x315;
  assign n7686 = n7606 ^ n7602;
  assign n7687 = n7686 ^ x316;
  assign n7688 = n7605 ^ n7603;
  assign n7689 = n7688 ^ x317;
  assign n7290 = x319 & n7288;
  assign n7291 = n7290 ^ x318;
  assign n7289 = n7288 ^ n7287;
  assign n7690 = n7290 ^ n7289;
  assign n7691 = n7291 & n7690;
  assign n7692 = n7691 ^ x318;
  assign n7693 = n7692 ^ n7688;
  assign n7694 = ~n7689 & n7693;
  assign n7695 = n7694 ^ x317;
  assign n7696 = n7695 ^ n7686;
  assign n7697 = ~n7687 & n7696;
  assign n7698 = n7697 ^ x316;
  assign n7699 = n7698 ^ n7684;
  assign n7700 = ~n7685 & n7699;
  assign n7701 = n7700 ^ x315;
  assign n7702 = n7701 ^ n7682;
  assign n7703 = n7683 & ~n7702;
  assign n7704 = n7703 ^ x314;
  assign n7705 = n7704 ^ n7680;
  assign n7706 = ~n7681 & n7705;
  assign n7707 = n7706 ^ x313;
  assign n7708 = n7707 ^ n7678;
  assign n7709 = ~n7679 & n7708;
  assign n7710 = n7709 ^ x312;
  assign n7711 = n7710 ^ n7676;
  assign n7712 = n7677 & ~n7711;
  assign n7713 = n7712 ^ x311;
  assign n7714 = n7713 ^ n7674;
  assign n7715 = ~n7675 & n7714;
  assign n7716 = n7715 ^ x310;
  assign n7516 = n7515 ^ n4750;
  assign n7559 = n7558 ^ n7515;
  assign n7560 = n7516 & n7559;
  assign n7561 = n7560 ^ n4750;
  assign n7622 = n7561 ^ n4739;
  assign n7341 = n7340 ^ n7337;
  assign n7468 = n7467 ^ n7337;
  assign n7469 = n7341 & ~n7468;
  assign n7470 = n7469 ^ n7340;
  assign n7333 = n6297 ^ n5704;
  assign n7334 = n6281 & ~n7333;
  assign n7335 = n7334 ^ n5704;
  assign n7331 = n7161 ^ x282;
  assign n7332 = n7331 ^ n7139;
  assign n7336 = n7335 ^ n7332;
  assign n7512 = n7470 ^ n7336;
  assign n7623 = n7622 ^ n7512;
  assign n7621 = ~n7618 & n7620;
  assign n7672 = n7623 ^ n7621;
  assign n7673 = n7672 ^ x309;
  assign n7838 = n7716 ^ n7673;
  assign n7842 = n7841 ^ n7838;
  assign n7846 = n7713 ^ x310;
  assign n7847 = n7846 ^ n7674;
  assign n7650 = n7188 ^ n7122;
  assign n7843 = n7011 ^ n6269;
  assign n7844 = n7650 & n7843;
  assign n7845 = n7844 ^ n6269;
  assign n7848 = n7847 ^ n7845;
  assign n7852 = n7710 ^ x311;
  assign n7853 = n7852 ^ n7676;
  assign n7593 = n7185 ^ x274;
  assign n7594 = n7593 ^ n7123;
  assign n7849 = n6996 ^ n6277;
  assign n7850 = ~n7594 & ~n7849;
  assign n7851 = n7850 ^ n6277;
  assign n7854 = n7853 ^ n7851;
  assign n7858 = n7707 ^ x312;
  assign n7859 = n7858 ^ n7678;
  assign n7495 = n7182 ^ n7126;
  assign n7855 = n6933 ^ n6283;
  assign n7856 = n7495 & ~n7855;
  assign n7857 = n7856 ^ n6283;
  assign n7860 = n7859 ^ n7857;
  assign n7864 = n7704 ^ n7681;
  assign n7301 = n7179 ^ x276;
  assign n7302 = n7301 ^ n7127;
  assign n7861 = n6824 ^ n6292;
  assign n7862 = ~n7302 & ~n7861;
  assign n7863 = n7862 ^ n6292;
  assign n7865 = n7864 ^ n7863;
  assign n7869 = n7701 ^ x314;
  assign n7870 = n7869 ^ n7682;
  assign n7307 = n7176 ^ n7130;
  assign n7866 = n6297 ^ n6267;
  assign n7867 = ~n7307 & ~n7866;
  assign n7868 = n7867 ^ n6297;
  assign n7871 = n7870 ^ n7868;
  assign n7875 = n7698 ^ n7685;
  assign n7312 = n7173 ^ n7132;
  assign n7872 = n6306 ^ n6274;
  assign n7873 = n7312 & n7872;
  assign n7874 = n7873 ^ n6306;
  assign n7876 = n7875 ^ n7874;
  assign n7880 = n7695 ^ x316;
  assign n7881 = n7880 ^ n7686;
  assign n7314 = n7170 ^ x279;
  assign n7315 = n7314 ^ n7133;
  assign n7877 = n6311 ^ n6281;
  assign n7878 = n7315 & n7877;
  assign n7879 = n7878 ^ n6311;
  assign n7882 = n7881 ^ n7879;
  assign n7320 = n7167 ^ x280;
  assign n7321 = n7320 ^ n7135;
  assign n7884 = n6319 ^ n6287;
  assign n7885 = n7321 & n7884;
  assign n7886 = n7885 ^ n6319;
  assign n7883 = n7692 ^ n7689;
  assign n7887 = n7886 ^ n7883;
  assign n7326 = n7164 ^ n7138;
  assign n7888 = n6325 ^ n6290;
  assign n7889 = ~n7326 & ~n7888;
  assign n7890 = n7889 ^ n6325;
  assign n7292 = n7291 ^ n7289;
  assign n7891 = n7890 ^ n7292;
  assign n7893 = n6302 ^ n6262;
  assign n7894 = n7332 & n7893;
  assign n7895 = n7894 ^ n6262;
  assign n7892 = n7288 ^ x319;
  assign n7896 = n7895 ^ n7892;
  assign n8113 = n5731 ^ n4611;
  assign n8114 = ~n6777 & ~n8113;
  assign n8115 = n8114 ^ n4611;
  assign n8112 = n7226 ^ n7100;
  assign n8116 = n8115 ^ n8112;
  assign n8117 = n8116 ^ n4672;
  assign n7903 = n6052 ^ n5374;
  assign n7904 = n6731 & ~n7903;
  assign n7905 = n7904 ^ n5374;
  assign n7784 = n7217 ^ x264;
  assign n7785 = n7784 ^ n7105;
  assign n7906 = n7905 ^ n7785;
  assign n7907 = n6057 ^ n5383;
  assign n7908 = n6740 & n7907;
  assign n7909 = n7908 ^ n5383;
  assign n7792 = n7214 ^ n7108;
  assign n7910 = n7909 ^ n7792;
  assign n7911 = n6059 ^ n5391;
  assign n7912 = n7441 & n7911;
  assign n7913 = n7912 ^ n5391;
  assign n7798 = n7211 ^ x266;
  assign n7799 = n7798 ^ n7109;
  assign n7914 = n7913 ^ n7799;
  assign n7915 = n6064 ^ n5394;
  assign n7916 = ~n7398 & ~n7915;
  assign n7917 = n7916 ^ n5394;
  assign n7806 = n7208 ^ n7112;
  assign n7918 = n7917 ^ n7806;
  assign n7919 = n6771 ^ n6040;
  assign n7920 = ~n7371 & ~n7919;
  assign n7921 = n7920 ^ n6040;
  assign n7812 = n7205 ^ x268;
  assign n7813 = n7812 ^ n7113;
  assign n7922 = n7921 ^ n7813;
  assign n7923 = n6714 ^ n6017;
  assign n7924 = ~n7278 & ~n7923;
  assign n7925 = n7924 ^ n6017;
  assign n7820 = n7202 ^ n7116;
  assign n7926 = n7925 ^ n7820;
  assign n7927 = n6609 ^ n5996;
  assign n7928 = n7245 & n7927;
  assign n7929 = n7928 ^ n5996;
  assign n7826 = n7199 ^ x270;
  assign n7827 = n7826 ^ n7117;
  assign n7930 = n7929 ^ n7827;
  assign n7931 = n6592 ^ n5886;
  assign n7932 = ~n7096 & ~n7931;
  assign n7933 = n7932 ^ n5886;
  assign n7833 = n7196 ^ x271;
  assign n7934 = n7933 ^ n7833;
  assign n7752 = n6538 ^ n5824;
  assign n7753 = n7078 & n7752;
  assign n7754 = n7753 ^ n5824;
  assign n7757 = n7756 ^ n7754;
  assign n7647 = n6451 ^ n5744;
  assign n7648 = n7061 & ~n7647;
  assign n7649 = n7648 ^ n5744;
  assign n7651 = n7650 ^ n7649;
  assign n7590 = n6347 ^ n5750;
  assign n7591 = n7045 & ~n7590;
  assign n7592 = n7591 ^ n5750;
  assign n7595 = n7594 ^ n7592;
  assign n7492 = n6353 ^ n5711;
  assign n7493 = ~n7028 & n7492;
  assign n7494 = n7493 ^ n5711;
  assign n7496 = n7495 ^ n7494;
  assign n7298 = n6358 ^ n5755;
  assign n7299 = n7011 & n7298;
  assign n7300 = n7299 ^ n5755;
  assign n7303 = n7302 ^ n7300;
  assign n7304 = n5795 ^ n5710;
  assign n7305 = ~n6996 & ~n7304;
  assign n7306 = n7305 ^ n5795;
  assign n7308 = n7307 ^ n7306;
  assign n7309 = n6269 ^ n5787;
  assign n7310 = ~n6933 & ~n7309;
  assign n7311 = n7310 ^ n5787;
  assign n7313 = n7312 ^ n7311;
  assign n7316 = n6277 ^ n5779;
  assign n7317 = n6824 & ~n7316;
  assign n7318 = n7317 ^ n5779;
  assign n7319 = n7318 ^ n7315;
  assign n7322 = n6283 ^ n5771;
  assign n7323 = n6267 & n7322;
  assign n7324 = n7323 ^ n5771;
  assign n7325 = n7324 ^ n7321;
  assign n7327 = n6292 ^ n5763;
  assign n7328 = n6274 & ~n7327;
  assign n7329 = n7328 ^ n5763;
  assign n7330 = n7329 ^ n7326;
  assign n7471 = n7470 ^ n7332;
  assign n7472 = n7336 & n7471;
  assign n7473 = n7472 ^ n7335;
  assign n7474 = n7473 ^ n7326;
  assign n7475 = ~n7330 & n7474;
  assign n7476 = n7475 ^ n7329;
  assign n7477 = n7476 ^ n7321;
  assign n7478 = n7325 & ~n7477;
  assign n7479 = n7478 ^ n7324;
  assign n7480 = n7479 ^ n7315;
  assign n7481 = ~n7319 & ~n7480;
  assign n7482 = n7481 ^ n7318;
  assign n7483 = n7482 ^ n7312;
  assign n7484 = ~n7313 & n7483;
  assign n7485 = n7484 ^ n7311;
  assign n7486 = n7485 ^ n7307;
  assign n7487 = ~n7308 & ~n7486;
  assign n7488 = n7487 ^ n7306;
  assign n7489 = n7488 ^ n7302;
  assign n7490 = n7303 & n7489;
  assign n7491 = n7490 ^ n7300;
  assign n7587 = n7495 ^ n7491;
  assign n7588 = ~n7496 & n7587;
  assign n7589 = n7588 ^ n7494;
  assign n7652 = n7594 ^ n7589;
  assign n7653 = ~n7595 & ~n7652;
  assign n7654 = n7653 ^ n7592;
  assign n7758 = n7654 ^ n7650;
  assign n7759 = n7651 & ~n7758;
  assign n7760 = n7759 ^ n7649;
  assign n7935 = n7760 ^ n7756;
  assign n7936 = n7757 & n7935;
  assign n7937 = n7936 ^ n7754;
  assign n7938 = n7937 ^ n7833;
  assign n7939 = ~n7934 & n7938;
  assign n7940 = n7939 ^ n7933;
  assign n7941 = n7940 ^ n7827;
  assign n7942 = ~n7930 & ~n7941;
  assign n7943 = n7942 ^ n7929;
  assign n7944 = n7943 ^ n7820;
  assign n7945 = n7926 & ~n7944;
  assign n7946 = n7945 ^ n7925;
  assign n7947 = n7946 ^ n7813;
  assign n7948 = ~n7922 & ~n7947;
  assign n7949 = n7948 ^ n7921;
  assign n7950 = n7949 ^ n7806;
  assign n7951 = n7918 & n7950;
  assign n7952 = n7951 ^ n7917;
  assign n7953 = n7952 ^ n7799;
  assign n7954 = n7914 & n7953;
  assign n7955 = n7954 ^ n7913;
  assign n7956 = n7955 ^ n7792;
  assign n7957 = n7910 & ~n7956;
  assign n7958 = n7957 ^ n7909;
  assign n7959 = n7958 ^ n7785;
  assign n7960 = n7906 & n7959;
  assign n7961 = n7960 ^ n7905;
  assign n7778 = n7220 ^ n7104;
  assign n7962 = n7961 ^ n7778;
  assign n7900 = n6047 ^ n5371;
  assign n7901 = n6729 & ~n7900;
  assign n7902 = n7901 ^ n5371;
  assign n8020 = n7902 ^ n7778;
  assign n8021 = ~n7962 & n8020;
  assign n8022 = n8021 ^ n7902;
  assign n7770 = n7223 ^ x262;
  assign n7771 = n7770 ^ n7101;
  assign n8023 = n8022 ^ n7771;
  assign n8017 = n5739 ^ n4617;
  assign n8018 = n6720 & n8017;
  assign n8019 = n8018 ^ n4617;
  assign n8109 = n8019 ^ n7771;
  assign n8110 = n8023 & ~n8109;
  assign n8111 = n8110 ^ n8019;
  assign n8118 = n8117 ^ n8111;
  assign n8024 = n8023 ^ n8019;
  assign n7963 = n7962 ^ n7902;
  assign n7964 = n7963 ^ n4565;
  assign n7965 = n7958 ^ n7905;
  assign n7966 = n7965 ^ n7785;
  assign n7967 = n7966 ^ n4520;
  assign n7968 = n7955 ^ n7909;
  assign n7969 = n7968 ^ n7792;
  assign n7970 = n7969 ^ n4480;
  assign n7971 = n7952 ^ n7913;
  assign n7972 = n7971 ^ n7799;
  assign n7973 = n7972 ^ n4445;
  assign n7974 = n7949 ^ n7917;
  assign n7975 = n7974 ^ n7806;
  assign n7976 = n7975 ^ n4411;
  assign n7977 = n7946 ^ n7922;
  assign n7978 = n7977 ^ n5364;
  assign n7979 = n7943 ^ n7926;
  assign n7980 = n7979 ^ n5066;
  assign n7981 = n7940 ^ n7930;
  assign n7982 = n7981 ^ n4876;
  assign n7983 = n7937 ^ n7934;
  assign n7984 = n7983 ^ n4638;
  assign n7761 = n7760 ^ n7757;
  assign n7985 = n7761 ^ n4845;
  assign n7655 = n7654 ^ n7651;
  assign n7656 = n7655 ^ n4830;
  assign n7596 = n7595 ^ n7589;
  assign n7643 = n7596 ^ n4840;
  assign n7497 = n7496 ^ n7491;
  assign n7498 = n7497 ^ n4838;
  assign n7499 = n7488 ^ n7300;
  assign n7500 = n7499 ^ n7302;
  assign n7501 = n7500 ^ n4786;
  assign n7502 = n7485 ^ n7308;
  assign n7503 = n7502 ^ n4779;
  assign n7504 = n7482 ^ n7313;
  assign n7505 = n7504 ^ n4775;
  assign n7506 = n7479 ^ n7319;
  assign n7507 = n7506 ^ n4766;
  assign n7508 = n7476 ^ n7325;
  assign n7509 = n7508 ^ n4758;
  assign n7510 = n7473 ^ n7330;
  assign n7511 = n7510 ^ n4734;
  assign n7513 = n7512 ^ n4739;
  assign n7562 = n7561 ^ n7512;
  assign n7563 = n7513 & ~n7562;
  assign n7564 = n7563 ^ n4739;
  assign n7565 = n7564 ^ n7510;
  assign n7566 = n7511 & ~n7565;
  assign n7567 = n7566 ^ n4734;
  assign n7568 = n7567 ^ n7508;
  assign n7569 = n7509 & n7568;
  assign n7570 = n7569 ^ n4758;
  assign n7571 = n7570 ^ n7506;
  assign n7572 = ~n7507 & n7571;
  assign n7573 = n7572 ^ n4766;
  assign n7574 = n7573 ^ n7504;
  assign n7575 = ~n7505 & ~n7574;
  assign n7576 = n7575 ^ n4775;
  assign n7577 = n7576 ^ n7502;
  assign n7578 = n7503 & n7577;
  assign n7579 = n7578 ^ n4779;
  assign n7580 = n7579 ^ n7500;
  assign n7581 = ~n7501 & ~n7580;
  assign n7582 = n7581 ^ n4786;
  assign n7583 = n7582 ^ n7497;
  assign n7584 = ~n7498 & n7583;
  assign n7585 = n7584 ^ n4838;
  assign n7644 = n7596 ^ n7585;
  assign n7645 = ~n7643 & n7644;
  assign n7646 = n7645 ^ n4840;
  assign n7762 = n7655 ^ n7646;
  assign n7763 = n7656 & n7762;
  assign n7764 = n7763 ^ n4830;
  assign n7986 = n7764 ^ n7761;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = n7987 ^ n4845;
  assign n7989 = n7988 ^ n7983;
  assign n7990 = n7984 & n7989;
  assign n7991 = n7990 ^ n4638;
  assign n7992 = n7991 ^ n7981;
  assign n7993 = n7982 & ~n7992;
  assign n7994 = n7993 ^ n4876;
  assign n7995 = n7994 ^ n7979;
  assign n7996 = n7980 & ~n7995;
  assign n7997 = n7996 ^ n5066;
  assign n7998 = n7997 ^ n7977;
  assign n7999 = ~n7978 & n7998;
  assign n8000 = n7999 ^ n5364;
  assign n8001 = n8000 ^ n7975;
  assign n8002 = ~n7976 & n8001;
  assign n8003 = n8002 ^ n4411;
  assign n8004 = n8003 ^ n7972;
  assign n8005 = n7973 & ~n8004;
  assign n8006 = n8005 ^ n4445;
  assign n8007 = n8006 ^ n7969;
  assign n8008 = ~n7970 & n8007;
  assign n8009 = n8008 ^ n4480;
  assign n8010 = n8009 ^ n7966;
  assign n8011 = ~n7967 & n8010;
  assign n8012 = n8011 ^ n4520;
  assign n8013 = n8012 ^ n7963;
  assign n8014 = n7964 & ~n8013;
  assign n8015 = n8014 ^ n4565;
  assign n8016 = n8015 ^ n4680;
  assign n8025 = n8024 ^ n8016;
  assign n8026 = n8012 ^ n4565;
  assign n8027 = n8026 ^ n7963;
  assign n8028 = n8009 ^ n4520;
  assign n8029 = n8028 ^ n7966;
  assign n7586 = n7585 ^ n4840;
  assign n7597 = n7596 ^ n7586;
  assign n7624 = n7621 & ~n7623;
  assign n7625 = n7564 ^ n7511;
  assign n7626 = ~n7624 & n7625;
  assign n7627 = n7567 ^ n4758;
  assign n7628 = n7627 ^ n7508;
  assign n7629 = n7626 & n7628;
  assign n7630 = n7570 ^ n7507;
  assign n7631 = n7629 & n7630;
  assign n7632 = n7573 ^ n4775;
  assign n7633 = n7632 ^ n7504;
  assign n7634 = n7631 & n7633;
  assign n7635 = n7576 ^ n4779;
  assign n7636 = n7635 ^ n7502;
  assign n7637 = ~n7634 & ~n7636;
  assign n7638 = n7579 ^ n7501;
  assign n7639 = n7637 & ~n7638;
  assign n7640 = n7582 ^ n7498;
  assign n7641 = ~n7639 & ~n7640;
  assign n7642 = n7597 & ~n7641;
  assign n7657 = n7656 ^ n7646;
  assign n7751 = n7642 & ~n7657;
  assign n7765 = n7764 ^ n4845;
  assign n7766 = n7765 ^ n7761;
  assign n8030 = n7751 & ~n7766;
  assign n8031 = n7988 ^ n7984;
  assign n8032 = n8030 & ~n8031;
  assign n8033 = n7991 ^ n4876;
  assign n8034 = n8033 ^ n7981;
  assign n8035 = n8032 & n8034;
  assign n8036 = n7994 ^ n7980;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = n7997 ^ n7978;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = n8000 ^ n7976;
  assign n8041 = ~n8039 & n8040;
  assign n8042 = n8003 ^ n4445;
  assign n8043 = n8042 ^ n7972;
  assign n8044 = ~n8041 & n8043;
  assign n8045 = n8006 ^ n4480;
  assign n8046 = n8045 ^ n7969;
  assign n8047 = ~n8044 & n8046;
  assign n8048 = n8029 & n8047;
  assign n8049 = n8027 & ~n8048;
  assign n8108 = n8025 & ~n8049;
  assign n8119 = n8118 ^ n8108;
  assign n8104 = n8024 ^ n4680;
  assign n8105 = n8024 ^ n8015;
  assign n8106 = ~n8104 & n8105;
  assign n8107 = n8106 ^ n4680;
  assign n8120 = n8119 ^ n8107;
  assign n8050 = n8049 ^ n8025;
  assign n8051 = n8050 ^ x289;
  assign n8095 = n8048 ^ n8027;
  assign n8052 = n8047 ^ n8029;
  assign n8053 = n8052 ^ x291;
  assign n8054 = n8046 ^ n8044;
  assign n8055 = n8054 ^ x292;
  assign n8056 = n8043 ^ n8041;
  assign n8057 = n8056 ^ x293;
  assign n8058 = n8040 ^ n8039;
  assign n8059 = n8058 ^ x294;
  assign n8060 = n8038 ^ n8037;
  assign n8061 = n8060 ^ x295;
  assign n8062 = n8036 ^ n8035;
  assign n8063 = n8062 ^ x296;
  assign n8064 = n8034 ^ n8032;
  assign n8065 = n8064 ^ x297;
  assign n8066 = n8031 ^ n8030;
  assign n8067 = n8066 ^ x298;
  assign n7767 = n7766 ^ n7751;
  assign n7768 = n7767 ^ x299;
  assign n7658 = n7657 ^ n7642;
  assign n7659 = n7658 ^ x300;
  assign n7660 = n7641 ^ n7597;
  assign n7661 = n7660 ^ x301;
  assign n7662 = n7640 ^ n7639;
  assign n7663 = n7662 ^ x302;
  assign n7737 = n7638 ^ n7637;
  assign n7664 = n7636 ^ n7634;
  assign n7665 = n7664 ^ x304;
  assign n7666 = n7633 ^ n7631;
  assign n7667 = n7666 ^ x305;
  assign n7668 = n7630 ^ n7629;
  assign n7669 = n7668 ^ x306;
  assign n7670 = n7628 ^ n7626;
  assign n7671 = n7670 ^ x307;
  assign n7720 = n7625 ^ n7624;
  assign n7717 = n7716 ^ n7672;
  assign n7718 = ~n7673 & n7717;
  assign n7719 = n7718 ^ x309;
  assign n7721 = n7720 ^ n7719;
  assign n7722 = n7720 ^ x308;
  assign n7723 = ~n7721 & n7722;
  assign n7724 = n7723 ^ x308;
  assign n7725 = n7724 ^ n7670;
  assign n7726 = ~n7671 & n7725;
  assign n7727 = n7726 ^ x307;
  assign n7728 = n7727 ^ n7668;
  assign n7729 = ~n7669 & n7728;
  assign n7730 = n7729 ^ x306;
  assign n7731 = n7730 ^ n7666;
  assign n7732 = ~n7667 & n7731;
  assign n7733 = n7732 ^ x305;
  assign n7734 = n7733 ^ n7664;
  assign n7735 = n7665 & ~n7734;
  assign n7736 = n7735 ^ x304;
  assign n7738 = n7737 ^ n7736;
  assign n7739 = n7737 ^ x303;
  assign n7740 = n7738 & ~n7739;
  assign n7741 = n7740 ^ x303;
  assign n7742 = n7741 ^ n7662;
  assign n7743 = ~n7663 & n7742;
  assign n7744 = n7743 ^ x302;
  assign n7745 = n7744 ^ n7660;
  assign n7746 = ~n7661 & n7745;
  assign n7747 = n7746 ^ x301;
  assign n7748 = n7747 ^ n7658;
  assign n7749 = ~n7659 & n7748;
  assign n7750 = n7749 ^ x300;
  assign n8068 = n7767 ^ n7750;
  assign n8069 = ~n7768 & n8068;
  assign n8070 = n8069 ^ x299;
  assign n8071 = n8070 ^ n8066;
  assign n8072 = ~n8067 & n8071;
  assign n8073 = n8072 ^ x298;
  assign n8074 = n8073 ^ n8064;
  assign n8075 = n8065 & ~n8074;
  assign n8076 = n8075 ^ x297;
  assign n8077 = n8076 ^ n8062;
  assign n8078 = ~n8063 & n8077;
  assign n8079 = n8078 ^ x296;
  assign n8080 = n8079 ^ n8060;
  assign n8081 = n8061 & ~n8080;
  assign n8082 = n8081 ^ x295;
  assign n8083 = n8082 ^ n8058;
  assign n8084 = n8059 & ~n8083;
  assign n8085 = n8084 ^ x294;
  assign n8086 = n8085 ^ n8056;
  assign n8087 = ~n8057 & n8086;
  assign n8088 = n8087 ^ x293;
  assign n8089 = n8088 ^ n8054;
  assign n8090 = n8055 & ~n8089;
  assign n8091 = n8090 ^ x292;
  assign n8092 = n8091 ^ n8052;
  assign n8093 = ~n8053 & n8092;
  assign n8094 = n8093 ^ x291;
  assign n8096 = n8095 ^ n8094;
  assign n8097 = n8095 ^ x290;
  assign n8098 = n8096 & ~n8097;
  assign n8099 = n8098 ^ x290;
  assign n8100 = n8099 ^ n8050;
  assign n8101 = n8051 & ~n8100;
  assign n8102 = n8101 ^ x289;
  assign n8103 = n8102 ^ x288;
  assign n8121 = n8120 ^ n8103;
  assign n7897 = n6304 ^ n6162;
  assign n7898 = ~n7337 & ~n7897;
  assign n7899 = n7898 ^ n6162;
  assign n8122 = n8121 ^ n7899;
  assign n8126 = n8099 ^ x289;
  assign n8127 = n8126 ^ n8050;
  assign n8123 = n6316 ^ n6100;
  assign n8124 = n7294 & n8123;
  assign n8125 = n8124 ^ n6100;
  assign n8128 = n8127 ^ n8125;
  assign n8132 = n8096 ^ x290;
  assign n8129 = n6318 ^ n5718;
  assign n8130 = ~n7346 & n8129;
  assign n8131 = n8130 ^ n5718;
  assign n8133 = n8132 ^ n8131;
  assign n8135 = n6330 ^ n5724;
  assign n8136 = ~n7454 & ~n8135;
  assign n8137 = n8136 ^ n5724;
  assign n8134 = n8091 ^ n8053;
  assign n8138 = n8137 ^ n8134;
  assign n8139 = n8088 ^ x292;
  assign n8140 = n8139 ^ n8054;
  assign n8141 = n6335 ^ n5726;
  assign n8142 = n7351 & n8141;
  assign n8143 = n8142 ^ n5726;
  assign n8144 = n8140 & ~n8143;
  assign n8145 = n8144 ^ n8134;
  assign n8146 = n8138 & ~n8145;
  assign n8147 = n8146 ^ n8144;
  assign n8148 = n8147 ^ n8132;
  assign n8149 = ~n8133 & n8148;
  assign n8150 = n8149 ^ n8131;
  assign n8151 = n8150 ^ n8127;
  assign n8152 = n8128 & ~n8151;
  assign n8153 = n8152 ^ n8125;
  assign n8154 = n8153 ^ n8121;
  assign n8155 = ~n8122 & n8154;
  assign n8156 = n8155 ^ n7899;
  assign n8157 = n8156 ^ n7892;
  assign n8158 = n7896 & ~n8157;
  assign n8159 = n8158 ^ n7895;
  assign n8160 = n8159 ^ n7292;
  assign n8161 = ~n7891 & n8160;
  assign n8162 = n8161 ^ n7890;
  assign n8163 = n8162 ^ n7883;
  assign n8164 = ~n7887 & n8163;
  assign n8165 = n8164 ^ n7886;
  assign n8166 = n8165 ^ n7881;
  assign n8167 = ~n7882 & n8166;
  assign n8168 = n8167 ^ n7879;
  assign n8169 = n8168 ^ n7875;
  assign n8170 = ~n7876 & n8169;
  assign n8171 = n8170 ^ n7874;
  assign n8172 = n8171 ^ n7870;
  assign n8173 = ~n7871 & ~n8172;
  assign n8174 = n8173 ^ n7868;
  assign n8175 = n8174 ^ n7864;
  assign n8176 = n7865 & ~n8175;
  assign n8177 = n8176 ^ n7863;
  assign n8178 = n8177 ^ n7859;
  assign n8179 = ~n7860 & ~n8178;
  assign n8180 = n8179 ^ n7857;
  assign n8181 = n8180 ^ n7853;
  assign n8182 = n7854 & ~n8181;
  assign n8183 = n8182 ^ n7851;
  assign n8184 = n8183 ^ n7847;
  assign n8185 = ~n7848 & n8184;
  assign n8186 = n8185 ^ n7845;
  assign n8187 = n8186 ^ n7838;
  assign n8188 = n7842 & n8187;
  assign n8189 = n8188 ^ n7841;
  assign n7834 = n7045 ^ n6358;
  assign n7835 = n7833 & ~n7834;
  assign n7836 = n7835 ^ n6358;
  assign n8257 = n8189 ^ n7836;
  assign n7832 = n7721 ^ x308;
  assign n8258 = n8257 ^ n7832;
  assign n8259 = n8258 ^ n5755;
  assign n8260 = n8186 ^ n7841;
  assign n8261 = n8260 ^ n7838;
  assign n8262 = n8261 ^ n5795;
  assign n8263 = n8183 ^ n7848;
  assign n8264 = n8263 ^ n5787;
  assign n8265 = n8180 ^ n7854;
  assign n8266 = n8265 ^ n5779;
  assign n8267 = n8177 ^ n7860;
  assign n8268 = n8267 ^ n5771;
  assign n8269 = n8174 ^ n7865;
  assign n8270 = n8269 ^ n5763;
  assign n8271 = n8171 ^ n7871;
  assign n8272 = n8271 ^ n5704;
  assign n8273 = n8168 ^ n7876;
  assign n8274 = n8273 ^ n5682;
  assign n8275 = n8165 ^ n7882;
  assign n8276 = n8275 ^ n5587;
  assign n8277 = n8162 ^ n7887;
  assign n8278 = n8277 ^ n5569;
  assign n8279 = n8159 ^ n7891;
  assign n8280 = n8279 ^ n5551;
  assign n8281 = n8156 ^ n7896;
  assign n8282 = n8281 ^ n5534;
  assign n8283 = n8153 ^ n8122;
  assign n8284 = n8283 ^ n5494;
  assign n8285 = n8150 ^ n8128;
  assign n8286 = n8285 ^ n5431;
  assign n8287 = n8147 ^ n8133;
  assign n8288 = n8287 ^ n4588;
  assign n8289 = n8143 ^ n8140;
  assign n8290 = ~n4609 & ~n8289;
  assign n8291 = n8290 ^ n4598;
  assign n8292 = n8144 ^ n8137;
  assign n8293 = n8292 ^ n8134;
  assign n8294 = n8293 ^ n8290;
  assign n8295 = n8291 & n8294;
  assign n8296 = n8295 ^ n4598;
  assign n8297 = n8296 ^ n8287;
  assign n8298 = ~n8288 & n8297;
  assign n8299 = n8298 ^ n4588;
  assign n8300 = n8299 ^ n8285;
  assign n8301 = n8286 & ~n8300;
  assign n8302 = n8301 ^ n5431;
  assign n8303 = n8302 ^ n8283;
  assign n8304 = n8284 & n8303;
  assign n8305 = n8304 ^ n5494;
  assign n8306 = n8305 ^ n8281;
  assign n8307 = ~n8282 & n8306;
  assign n8308 = n8307 ^ n5534;
  assign n8309 = n8308 ^ n8279;
  assign n8310 = ~n8280 & ~n8309;
  assign n8311 = n8310 ^ n5551;
  assign n8312 = n8311 ^ n8277;
  assign n8313 = n8278 & n8312;
  assign n8314 = n8313 ^ n5569;
  assign n8315 = n8314 ^ n8275;
  assign n8316 = n8276 & ~n8315;
  assign n8317 = n8316 ^ n5587;
  assign n8318 = n8317 ^ n8273;
  assign n8319 = n8274 & ~n8318;
  assign n8320 = n8319 ^ n5682;
  assign n8321 = n8320 ^ n8271;
  assign n8322 = ~n8272 & ~n8321;
  assign n8323 = n8322 ^ n5704;
  assign n8324 = n8323 ^ n8269;
  assign n8325 = ~n8270 & n8324;
  assign n8326 = n8325 ^ n5763;
  assign n8327 = n8326 ^ n8267;
  assign n8328 = n8268 & ~n8327;
  assign n8329 = n8328 ^ n5771;
  assign n8330 = n8329 ^ n8265;
  assign n8331 = ~n8266 & ~n8330;
  assign n8332 = n8331 ^ n5779;
  assign n8333 = n8332 ^ n8263;
  assign n8334 = n8264 & ~n8333;
  assign n8335 = n8334 ^ n5787;
  assign n8336 = n8335 ^ n8261;
  assign n8337 = n8262 & n8336;
  assign n8338 = n8337 ^ n5795;
  assign n8339 = n8338 ^ n8258;
  assign n8340 = ~n8259 & ~n8339;
  assign n8341 = n8340 ^ n5755;
  assign n7837 = n7836 ^ n7832;
  assign n8190 = n8189 ^ n7832;
  assign n8191 = ~n7837 & n8190;
  assign n8192 = n8191 ^ n7836;
  assign n7828 = n7061 ^ n6353;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = n7829 ^ n6353;
  assign n7825 = n7724 ^ n7671;
  assign n7831 = n7830 ^ n7825;
  assign n8255 = n8192 ^ n7831;
  assign n8256 = n8255 ^ n5711;
  assign n8377 = n8341 ^ n8256;
  assign n8378 = n8332 ^ n8264;
  assign n8379 = n8320 ^ n8272;
  assign n8380 = n8317 ^ n8274;
  assign n8381 = n8314 ^ n8276;
  assign n8382 = n8299 ^ n8286;
  assign n8383 = n8296 ^ n4588;
  assign n8384 = n8383 ^ n8287;
  assign n8385 = n8289 ^ n4609;
  assign n8386 = n8293 ^ n8291;
  assign n8387 = n8385 & ~n8386;
  assign n8388 = ~n8384 & n8387;
  assign n8389 = ~n8382 & ~n8388;
  assign n8390 = n8302 ^ n8284;
  assign n8391 = n8389 & ~n8390;
  assign n8392 = n8305 ^ n8282;
  assign n8393 = ~n8391 & n8392;
  assign n8394 = n8308 ^ n8280;
  assign n8395 = n8393 & n8394;
  assign n8396 = n8311 ^ n8278;
  assign n8397 = ~n8395 & ~n8396;
  assign n8398 = n8381 & n8397;
  assign n8399 = ~n8380 & ~n8398;
  assign n8400 = n8379 & n8399;
  assign n8401 = n8323 ^ n8270;
  assign n8402 = ~n8400 & n8401;
  assign n8403 = n8326 ^ n8268;
  assign n8404 = n8402 & ~n8403;
  assign n8405 = n8329 ^ n8266;
  assign n8406 = n8404 & n8405;
  assign n8407 = n8378 & n8406;
  assign n8408 = n8335 ^ n8262;
  assign n8409 = ~n8407 & ~n8408;
  assign n8410 = n8338 ^ n8259;
  assign n8411 = n8409 & ~n8410;
  assign n8412 = n8377 & ~n8411;
  assign n8342 = n8341 ^ n8255;
  assign n8343 = n8256 & ~n8342;
  assign n8344 = n8343 ^ n5711;
  assign n8193 = n8192 ^ n7825;
  assign n8194 = n7831 & ~n8193;
  assign n8195 = n8194 ^ n7830;
  assign n7821 = n7078 ^ n6347;
  assign n7822 = n7820 & ~n7821;
  assign n7823 = n7822 ^ n6347;
  assign n7818 = n7727 ^ x306;
  assign n7819 = n7818 ^ n7668;
  assign n7824 = n7823 ^ n7819;
  assign n8253 = n8195 ^ n7824;
  assign n8254 = n8253 ^ n5750;
  assign n8413 = n8344 ^ n8254;
  assign n8414 = ~n8412 & n8413;
  assign n8345 = n8344 ^ n8253;
  assign n8346 = ~n8254 & ~n8345;
  assign n8347 = n8346 ^ n5750;
  assign n8375 = n8347 ^ n5744;
  assign n8196 = n8195 ^ n7819;
  assign n8197 = n7824 & ~n8196;
  assign n8198 = n8197 ^ n7823;
  assign n7814 = n7096 ^ n6451;
  assign n7815 = n7813 & n7814;
  assign n7816 = n7815 ^ n6451;
  assign n7811 = n7730 ^ n7667;
  assign n7817 = n7816 ^ n7811;
  assign n8251 = n8198 ^ n7817;
  assign n8376 = n8375 ^ n8251;
  assign n8446 = n8414 ^ n8376;
  assign n8447 = n8446 ^ x332;
  assign n8448 = n8413 ^ n8412;
  assign n8449 = n8448 ^ x333;
  assign n8450 = n8411 ^ n8377;
  assign n8451 = n8450 ^ x334;
  assign n8528 = n8410 ^ n8409;
  assign n8452 = n8408 ^ n8407;
  assign n8453 = n8452 ^ x336;
  assign n8454 = n8406 ^ n8378;
  assign n8455 = n8454 ^ x337;
  assign n8456 = n8405 ^ n8404;
  assign n8457 = n8456 ^ x338;
  assign n8458 = n8403 ^ n8402;
  assign n8459 = n8458 ^ x339;
  assign n8460 = n8401 ^ n8400;
  assign n8461 = n8460 ^ x340;
  assign n8462 = n8399 ^ n8379;
  assign n8463 = n8462 ^ x341;
  assign n8464 = n8398 ^ n8380;
  assign n8465 = n8464 ^ x342;
  assign n8466 = n8397 ^ n8381;
  assign n8467 = n8466 ^ x343;
  assign n8468 = n8396 ^ n8395;
  assign n8469 = n8468 ^ x344;
  assign n8470 = n8394 ^ n8393;
  assign n8471 = n8470 ^ x345;
  assign n8472 = n8392 ^ n8391;
  assign n8473 = n8472 ^ x346;
  assign n8474 = n8390 ^ n8389;
  assign n8475 = n8474 ^ x347;
  assign n8476 = n8388 ^ n8382;
  assign n8477 = n8476 ^ x348;
  assign n8478 = n8387 ^ n8384;
  assign n8479 = n8478 ^ x349;
  assign n8480 = x351 & ~n8385;
  assign n8481 = n8480 ^ x350;
  assign n8482 = n8386 ^ n8385;
  assign n8483 = n8482 ^ n8480;
  assign n8484 = n8481 & n8483;
  assign n8485 = n8484 ^ x350;
  assign n8486 = n8485 ^ n8478;
  assign n8487 = ~n8479 & n8486;
  assign n8488 = n8487 ^ x349;
  assign n8489 = n8488 ^ n8476;
  assign n8490 = ~n8477 & n8489;
  assign n8491 = n8490 ^ x348;
  assign n8492 = n8491 ^ n8474;
  assign n8493 = n8475 & ~n8492;
  assign n8494 = n8493 ^ x347;
  assign n8495 = n8494 ^ n8472;
  assign n8496 = ~n8473 & n8495;
  assign n8497 = n8496 ^ x346;
  assign n8498 = n8497 ^ n8470;
  assign n8499 = n8471 & ~n8498;
  assign n8500 = n8499 ^ x345;
  assign n8501 = n8500 ^ n8468;
  assign n8502 = ~n8469 & n8501;
  assign n8503 = n8502 ^ x344;
  assign n8504 = n8503 ^ n8466;
  assign n8505 = ~n8467 & n8504;
  assign n8506 = n8505 ^ x343;
  assign n8507 = n8506 ^ n8464;
  assign n8508 = n8465 & ~n8507;
  assign n8509 = n8508 ^ x342;
  assign n8510 = n8509 ^ n8462;
  assign n8511 = n8463 & ~n8510;
  assign n8512 = n8511 ^ x341;
  assign n8513 = n8512 ^ n8460;
  assign n8514 = n8461 & ~n8513;
  assign n8515 = n8514 ^ x340;
  assign n8516 = n8515 ^ n8458;
  assign n8517 = n8459 & ~n8516;
  assign n8518 = n8517 ^ x339;
  assign n8519 = n8518 ^ n8456;
  assign n8520 = ~n8457 & n8519;
  assign n8521 = n8520 ^ x338;
  assign n8522 = n8521 ^ n8454;
  assign n8523 = ~n8455 & n8522;
  assign n8524 = n8523 ^ x337;
  assign n8525 = n8524 ^ n8452;
  assign n8526 = n8453 & ~n8525;
  assign n8527 = n8526 ^ x336;
  assign n8529 = n8528 ^ n8527;
  assign n8530 = n8528 ^ x335;
  assign n8531 = n8529 & ~n8530;
  assign n8532 = n8531 ^ x335;
  assign n8533 = n8532 ^ n8450;
  assign n8534 = n8451 & ~n8533;
  assign n8535 = n8534 ^ x334;
  assign n8536 = n8535 ^ n8448;
  assign n8537 = ~n8449 & n8536;
  assign n8538 = n8537 ^ x333;
  assign n8539 = n8538 ^ n8446;
  assign n8540 = ~n8447 & n8539;
  assign n8541 = n8540 ^ x332;
  assign n8415 = ~n8376 & n8414;
  assign n8252 = n8251 ^ n5744;
  assign n8348 = n8347 ^ n8251;
  assign n8349 = ~n8252 & n8348;
  assign n8350 = n8349 ^ n5744;
  assign n8199 = n8198 ^ n7811;
  assign n8200 = n7817 & ~n8199;
  assign n8201 = n8200 ^ n7816;
  assign n7807 = n7245 ^ n6538;
  assign n7808 = n7806 & ~n7807;
  assign n7809 = n7808 ^ n6538;
  assign n7804 = n7733 ^ x304;
  assign n7805 = n7804 ^ n7664;
  assign n7810 = n7809 ^ n7805;
  assign n8249 = n8201 ^ n7810;
  assign n8250 = n8249 ^ n5824;
  assign n8374 = n8350 ^ n8250;
  assign n8444 = n8415 ^ n8374;
  assign n8445 = n8444 ^ x331;
  assign n9126 = n8541 ^ n8445;
  assign n8233 = n8073 ^ n8065;
  assign n9127 = n8233 ^ n7792;
  assign n9128 = ~n9126 & ~n9127;
  assign n9129 = n9128 ^ n7792;
  assign n8759 = n7594 ^ n6824;
  assign n8760 = n7832 & ~n8759;
  assign n8761 = n8760 ^ n6824;
  assign n8734 = n8497 ^ n8471;
  assign n8762 = n8761 ^ n8734;
  assign n8765 = n7495 ^ n6267;
  assign n8766 = ~n7838 & n8765;
  assign n8767 = n8766 ^ n6267;
  assign n8763 = n8494 ^ x346;
  assign n8764 = n8763 ^ n8472;
  assign n8768 = n8767 ^ n8764;
  assign n8770 = n7302 ^ n6274;
  assign n8771 = ~n7847 & ~n8770;
  assign n8772 = n8771 ^ n6274;
  assign n8769 = n8491 ^ n8475;
  assign n8773 = n8772 ^ n8769;
  assign n8776 = n7307 ^ n6281;
  assign n8777 = n7853 & ~n8776;
  assign n8778 = n8777 ^ n6281;
  assign n8774 = n8488 ^ x348;
  assign n8775 = n8774 ^ n8476;
  assign n8779 = n8778 ^ n8775;
  assign n8783 = n8485 ^ x349;
  assign n8784 = n8783 ^ n8478;
  assign n8780 = n7312 ^ n6287;
  assign n8781 = ~n7859 & n8780;
  assign n8782 = n8781 ^ n6287;
  assign n8785 = n8784 ^ n8782;
  assign n8787 = n7315 ^ n6290;
  assign n8788 = ~n7864 & ~n8787;
  assign n8789 = n8788 ^ n6290;
  assign n8786 = n8482 ^ n8481;
  assign n8790 = n8789 ^ n8786;
  assign n8792 = n7321 ^ n6302;
  assign n8793 = n7870 & n8792;
  assign n8794 = n8793 ^ n6302;
  assign n8791 = n8385 ^ x351;
  assign n8795 = n8794 ^ n8791;
  assign n8719 = n8085 ^ n8057;
  assign n8716 = n6340 ^ n5731;
  assign n8717 = n7447 & n8716;
  assign n8718 = n8717 ^ n5731;
  assign n8720 = n8719 ^ n8718;
  assign n8721 = n8720 ^ n4611;
  assign n8660 = n8082 ^ x294;
  assign n8661 = n8660 ^ n8058;
  assign n8616 = n8079 ^ n8061;
  assign n8579 = n8076 ^ x296;
  assign n8580 = n8579 ^ n8062;
  assign n8575 = n6720 ^ n6052;
  assign n8576 = n7282 & ~n8575;
  assign n8577 = n8576 ^ n6052;
  assign n8612 = n8580 ^ n8577;
  assign n8229 = n6729 ^ n6057;
  assign n8230 = n7249 & ~n8229;
  assign n8231 = n8230 ^ n6057;
  assign n8571 = n8233 ^ n8231;
  assign n8220 = n8070 ^ x298;
  assign n8221 = n8220 ^ n8066;
  assign n7772 = n6740 ^ n6064;
  assign n7773 = ~n7771 & ~n7772;
  assign n7774 = n7773 ^ n6064;
  assign n7769 = n7768 ^ n7750;
  assign n7775 = n7774 ^ n7769;
  assign n7779 = n7441 ^ n6771;
  assign n7780 = n7778 & n7779;
  assign n7781 = n7780 ^ n6771;
  assign n7776 = n7747 ^ x300;
  assign n7777 = n7776 ^ n7658;
  assign n7782 = n7781 ^ n7777;
  assign n7786 = n7398 ^ n6714;
  assign n7787 = n7785 & n7786;
  assign n7788 = n7787 ^ n6714;
  assign n7783 = n7744 ^ n7661;
  assign n7789 = n7788 ^ n7783;
  assign n7793 = n7371 ^ n6609;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = n7794 ^ n6609;
  assign n7790 = n7741 ^ x302;
  assign n7791 = n7790 ^ n7662;
  assign n7796 = n7795 ^ n7791;
  assign n7800 = n7278 ^ n6592;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = n7801 ^ n6592;
  assign n7797 = n7738 ^ x303;
  assign n7803 = n7802 ^ n7797;
  assign n8202 = n8201 ^ n7805;
  assign n8203 = ~n7810 & n8202;
  assign n8204 = n8203 ^ n7809;
  assign n8205 = n8204 ^ n7797;
  assign n8206 = ~n7803 & ~n8205;
  assign n8207 = n8206 ^ n7802;
  assign n8208 = n8207 ^ n7791;
  assign n8209 = ~n7796 & n8208;
  assign n8210 = n8209 ^ n7795;
  assign n8211 = n8210 ^ n7783;
  assign n8212 = n7789 & n8211;
  assign n8213 = n8212 ^ n7788;
  assign n8214 = n8213 ^ n7777;
  assign n8215 = ~n7782 & ~n8214;
  assign n8216 = n8215 ^ n7781;
  assign n8217 = n8216 ^ n7769;
  assign n8218 = n7775 & n8217;
  assign n8219 = n8218 ^ n7774;
  assign n8222 = n8221 ^ n8219;
  assign n8223 = n6731 ^ n6059;
  assign n8224 = n8112 & ~n8223;
  assign n8225 = n8224 ^ n6059;
  assign n8226 = n8225 ^ n8219;
  assign n8227 = n8222 & ~n8226;
  assign n8228 = n8227 ^ n8221;
  assign n8572 = n8233 ^ n8228;
  assign n8573 = ~n8571 & n8572;
  assign n8574 = n8573 ^ n8231;
  assign n8613 = n8580 ^ n8574;
  assign n8614 = n8612 & ~n8613;
  assign n8615 = n8614 ^ n8577;
  assign n8617 = n8616 ^ n8615;
  assign n8609 = n6777 ^ n6047;
  assign n8610 = n7414 & n8609;
  assign n8611 = n8610 ^ n6047;
  assign n8657 = n8616 ^ n8611;
  assign n8658 = n8617 & ~n8657;
  assign n8659 = n8658 ^ n8611;
  assign n8662 = n8661 ^ n8659;
  assign n8654 = n6342 ^ n5739;
  assign n8655 = ~n7404 & n8654;
  assign n8656 = n8655 ^ n5739;
  assign n8713 = n8661 ^ n8656;
  assign n8714 = n8662 & n8713;
  assign n8715 = n8714 ^ n8656;
  assign n8722 = n8721 ^ n8715;
  assign n8663 = n8662 ^ n8656;
  assign n8618 = n8617 ^ n8611;
  assign n8649 = n8618 ^ n5371;
  assign n8578 = n8577 ^ n8574;
  assign n8581 = n8580 ^ n8578;
  assign n8604 = n8581 ^ n5374;
  assign n8232 = n8231 ^ n8228;
  assign n8234 = n8233 ^ n8232;
  assign n8566 = n8234 ^ n5383;
  assign n8235 = n8225 ^ n8221;
  assign n8236 = n8235 ^ n8219;
  assign n8237 = n8236 ^ n5391;
  assign n8238 = n8216 ^ n7774;
  assign n8239 = n8238 ^ n7769;
  assign n8240 = n8239 ^ n5394;
  assign n8241 = n8213 ^ n7782;
  assign n8242 = n8241 ^ n6040;
  assign n8243 = n8210 ^ n7789;
  assign n8244 = n8243 ^ n6017;
  assign n8245 = n8207 ^ n7796;
  assign n8246 = n8245 ^ n5996;
  assign n8247 = n8204 ^ n7803;
  assign n8248 = n8247 ^ n5886;
  assign n8351 = n8350 ^ n8249;
  assign n8352 = ~n8250 & ~n8351;
  assign n8353 = n8352 ^ n5824;
  assign n8354 = n8353 ^ n8247;
  assign n8355 = ~n8248 & n8354;
  assign n8356 = n8355 ^ n5886;
  assign n8357 = n8356 ^ n8245;
  assign n8358 = ~n8246 & ~n8357;
  assign n8359 = n8358 ^ n5996;
  assign n8360 = n8359 ^ n8243;
  assign n8361 = n8244 & ~n8360;
  assign n8362 = n8361 ^ n6017;
  assign n8363 = n8362 ^ n8241;
  assign n8364 = ~n8242 & ~n8363;
  assign n8365 = n8364 ^ n6040;
  assign n8366 = n8365 ^ n8239;
  assign n8367 = n8240 & n8366;
  assign n8368 = n8367 ^ n5394;
  assign n8369 = n8368 ^ n8236;
  assign n8370 = n8237 & n8369;
  assign n8371 = n8370 ^ n5391;
  assign n8567 = n8371 ^ n8234;
  assign n8568 = ~n8566 & n8567;
  assign n8569 = n8568 ^ n5383;
  assign n8605 = n8581 ^ n8569;
  assign n8606 = ~n8604 & ~n8605;
  assign n8607 = n8606 ^ n5374;
  assign n8650 = n8618 ^ n8607;
  assign n8651 = n8649 & ~n8650;
  assign n8652 = n8651 ^ n5371;
  assign n8653 = n8652 ^ n4617;
  assign n8664 = n8663 ^ n8653;
  assign n8608 = n8607 ^ n5371;
  assign n8619 = n8618 ^ n8608;
  assign n8570 = n8569 ^ n5374;
  assign n8582 = n8581 ^ n8570;
  assign n8372 = n8371 ^ n5383;
  assign n8373 = n8372 ^ n8234;
  assign n8416 = ~n8374 & n8415;
  assign n8417 = n8353 ^ n8248;
  assign n8418 = n8416 & n8417;
  assign n8419 = n8356 ^ n8246;
  assign n8420 = n8418 & n8419;
  assign n8421 = n8359 ^ n8244;
  assign n8422 = ~n8420 & ~n8421;
  assign n8423 = n8362 ^ n8242;
  assign n8424 = ~n8422 & ~n8423;
  assign n8425 = n8365 ^ n8240;
  assign n8426 = ~n8424 & n8425;
  assign n8427 = n8368 ^ n5391;
  assign n8428 = n8427 ^ n8236;
  assign n8429 = ~n8426 & n8428;
  assign n8583 = ~n8373 & ~n8429;
  assign n8620 = ~n8582 & n8583;
  assign n8665 = n8619 & ~n8620;
  assign n8712 = n8664 & ~n8665;
  assign n8723 = n8722 ^ n8712;
  assign n8708 = n8663 ^ n4617;
  assign n8709 = n8663 ^ n8652;
  assign n8710 = ~n8708 & n8709;
  assign n8711 = n8710 ^ n4617;
  assign n8724 = n8723 ^ n8711;
  assign n8666 = n8665 ^ n8664;
  assign n8703 = n8666 ^ x321;
  assign n8621 = n8620 ^ n8619;
  assign n8644 = n8621 ^ x322;
  assign n8584 = n8583 ^ n8582;
  assign n8585 = n8584 ^ x323;
  assign n8430 = n8429 ^ n8373;
  assign n8431 = n8430 ^ x324;
  assign n8432 = n8428 ^ n8426;
  assign n8433 = n8432 ^ x325;
  assign n8434 = n8425 ^ n8424;
  assign n8435 = n8434 ^ x326;
  assign n8436 = n8423 ^ n8422;
  assign n8437 = n8436 ^ x327;
  assign n8438 = n8421 ^ n8420;
  assign n8439 = n8438 ^ x328;
  assign n8440 = n8419 ^ n8418;
  assign n8441 = n8440 ^ x329;
  assign n8442 = n8417 ^ n8416;
  assign n8443 = n8442 ^ x330;
  assign n8542 = n8541 ^ n8444;
  assign n8543 = ~n8445 & n8542;
  assign n8544 = n8543 ^ x331;
  assign n8545 = n8544 ^ n8442;
  assign n8546 = n8443 & ~n8545;
  assign n8547 = n8546 ^ x330;
  assign n8548 = n8547 ^ n8440;
  assign n8549 = n8441 & ~n8548;
  assign n8550 = n8549 ^ x329;
  assign n8551 = n8550 ^ n8438;
  assign n8552 = ~n8439 & n8551;
  assign n8553 = n8552 ^ x328;
  assign n8554 = n8553 ^ n8436;
  assign n8555 = n8437 & ~n8554;
  assign n8556 = n8555 ^ x327;
  assign n8557 = n8556 ^ n8434;
  assign n8558 = n8435 & ~n8557;
  assign n8559 = n8558 ^ x326;
  assign n8560 = n8559 ^ n8432;
  assign n8561 = ~n8433 & n8560;
  assign n8562 = n8561 ^ x325;
  assign n8563 = n8562 ^ n8430;
  assign n8564 = ~n8431 & n8563;
  assign n8565 = n8564 ^ x324;
  assign n8600 = n8584 ^ n8565;
  assign n8601 = n8585 & ~n8600;
  assign n8602 = n8601 ^ x323;
  assign n8645 = n8621 ^ n8602;
  assign n8646 = ~n8644 & n8645;
  assign n8647 = n8646 ^ x322;
  assign n8704 = n8666 ^ n8647;
  assign n8705 = n8703 & ~n8704;
  assign n8706 = n8705 ^ x321;
  assign n8707 = n8706 ^ x320;
  assign n8725 = n8724 ^ n8707;
  assign n8700 = n7326 ^ n6304;
  assign n8701 = ~n7875 & n8700;
  assign n8702 = n8701 ^ n6304;
  assign n8726 = n8725 ^ n8702;
  assign n8648 = n8647 ^ x321;
  assign n8667 = n8666 ^ n8648;
  assign n8640 = n7332 ^ n6316;
  assign n8641 = ~n7881 & n8640;
  assign n8642 = n8641 ^ n6316;
  assign n8696 = n8667 ^ n8642;
  assign n8603 = n8602 ^ x322;
  assign n8622 = n8621 ^ n8603;
  assign n8597 = n7337 ^ n6318;
  assign n8598 = ~n7883 & ~n8597;
  assign n8599 = n8598 ^ n6318;
  assign n8623 = n8622 ^ n8599;
  assign n8586 = n8585 ^ n8565;
  assign n7295 = n7294 ^ n6330;
  assign n7296 = ~n7292 & ~n7295;
  assign n7297 = n7296 ^ n6330;
  assign n8587 = n8586 ^ n7297;
  assign n8588 = n8562 ^ x324;
  assign n8589 = n8588 ^ n8430;
  assign n8590 = n7346 ^ n6335;
  assign n8591 = n7892 & n8590;
  assign n8592 = n8591 ^ n6335;
  assign n8593 = ~n8589 & ~n8592;
  assign n8594 = n8593 ^ n8586;
  assign n8595 = n8587 & n8594;
  assign n8596 = n8595 ^ n8593;
  assign n8637 = n8622 ^ n8596;
  assign n8638 = ~n8623 & n8637;
  assign n8639 = n8638 ^ n8599;
  assign n8697 = n8667 ^ n8639;
  assign n8698 = n8696 & ~n8697;
  assign n8699 = n8698 ^ n8642;
  assign n8796 = n8725 ^ n8699;
  assign n8797 = n8726 & n8796;
  assign n8798 = n8797 ^ n8702;
  assign n8799 = n8798 ^ n8791;
  assign n8800 = ~n8795 & ~n8799;
  assign n8801 = n8800 ^ n8794;
  assign n8802 = n8801 ^ n8786;
  assign n8803 = n8790 & n8802;
  assign n8804 = n8803 ^ n8789;
  assign n8805 = n8804 ^ n8784;
  assign n8806 = ~n8785 & ~n8805;
  assign n8807 = n8806 ^ n8782;
  assign n8808 = n8807 ^ n8775;
  assign n8809 = ~n8779 & n8808;
  assign n8810 = n8809 ^ n8778;
  assign n8811 = n8810 ^ n8769;
  assign n8812 = n8773 & ~n8811;
  assign n8813 = n8812 ^ n8772;
  assign n8814 = n8813 ^ n8764;
  assign n8815 = ~n8768 & n8814;
  assign n8816 = n8815 ^ n8767;
  assign n8817 = n8816 ^ n8734;
  assign n8818 = n8762 & ~n8817;
  assign n8819 = n8818 ^ n8761;
  assign n8755 = n7650 ^ n6933;
  assign n8756 = ~n7825 & ~n8755;
  assign n8757 = n8756 ^ n6933;
  assign n8753 = n8500 ^ x344;
  assign n8754 = n8753 ^ n8468;
  assign n8758 = n8757 ^ n8754;
  assign n8837 = n8819 ^ n8758;
  assign n8838 = n8837 ^ n6283;
  assign n8839 = n8816 ^ n8761;
  assign n8840 = n8839 ^ n8734;
  assign n8841 = n8840 ^ n6292;
  assign n8842 = n8813 ^ n8768;
  assign n8843 = n8842 ^ n6297;
  assign n8844 = n8810 ^ n8772;
  assign n8845 = n8844 ^ n8769;
  assign n8846 = n8845 ^ n6306;
  assign n8847 = n8807 ^ n8778;
  assign n8848 = n8847 ^ n8775;
  assign n8849 = n8848 ^ n6311;
  assign n8850 = n8804 ^ n8782;
  assign n8851 = n8850 ^ n8784;
  assign n8852 = n8851 ^ n6319;
  assign n8853 = n8801 ^ n8790;
  assign n8854 = n8853 ^ n6325;
  assign n8855 = n8798 ^ n8795;
  assign n8856 = n8855 ^ n6262;
  assign n8727 = n8726 ^ n8699;
  assign n8728 = n8727 ^ n6162;
  assign n8643 = n8642 ^ n8639;
  assign n8668 = n8667 ^ n8643;
  assign n8669 = n8668 ^ n6100;
  assign n8624 = n8623 ^ n8596;
  assign n8625 = n8624 ^ n5718;
  assign n8626 = n8592 ^ n8589;
  assign n8627 = ~n5726 & n8626;
  assign n8628 = n8627 ^ n5724;
  assign n8629 = n8593 ^ n7297;
  assign n8630 = n8629 ^ n8586;
  assign n8631 = n8630 ^ n8627;
  assign n8632 = n8628 & n8631;
  assign n8633 = n8632 ^ n5724;
  assign n8634 = n8633 ^ n8624;
  assign n8635 = ~n8625 & n8634;
  assign n8636 = n8635 ^ n5718;
  assign n8693 = n8668 ^ n8636;
  assign n8694 = n8669 & ~n8693;
  assign n8695 = n8694 ^ n6100;
  assign n8857 = n8727 ^ n8695;
  assign n8858 = n8728 & ~n8857;
  assign n8859 = n8858 ^ n6162;
  assign n8860 = n8859 ^ n8855;
  assign n8861 = n8856 & ~n8860;
  assign n8862 = n8861 ^ n6262;
  assign n8863 = n8862 ^ n8853;
  assign n8864 = n8854 & ~n8863;
  assign n8865 = n8864 ^ n6325;
  assign n8866 = n8865 ^ n8851;
  assign n8867 = n8852 & ~n8866;
  assign n8868 = n8867 ^ n6319;
  assign n8869 = n8868 ^ n8848;
  assign n8870 = ~n8849 & n8869;
  assign n8871 = n8870 ^ n6311;
  assign n8872 = n8871 ^ n8845;
  assign n8873 = n8846 & ~n8872;
  assign n8874 = n8873 ^ n6306;
  assign n8875 = n8874 ^ n8842;
  assign n8876 = n8843 & n8875;
  assign n8877 = n8876 ^ n6297;
  assign n8878 = n8877 ^ n8840;
  assign n8879 = ~n8841 & n8878;
  assign n8880 = n8879 ^ n6292;
  assign n8881 = n8880 ^ n8837;
  assign n8882 = n8838 & n8881;
  assign n8883 = n8882 ^ n6283;
  assign n8907 = n8883 ^ n6277;
  assign n8820 = n8819 ^ n8754;
  assign n8821 = n8758 & n8820;
  assign n8822 = n8821 ^ n8757;
  assign n8749 = n7756 ^ n6996;
  assign n8750 = ~n7819 & n8749;
  assign n8751 = n8750 ^ n6996;
  assign n8834 = n8822 ^ n8751;
  assign n8747 = n8503 ^ x343;
  assign n8748 = n8747 ^ n8466;
  assign n8835 = n8834 ^ n8748;
  assign n8908 = n8907 ^ n8835;
  assign n8909 = n8880 ^ n8838;
  assign n8910 = n8877 ^ n8841;
  assign n8729 = n8728 ^ n8695;
  assign n8670 = n8669 ^ n8636;
  assign n8671 = n8633 ^ n5718;
  assign n8672 = n8671 ^ n8624;
  assign n8673 = n8626 ^ n5726;
  assign n8674 = n8630 ^ n8628;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = ~n8672 & n8675;
  assign n8730 = ~n8670 & ~n8676;
  assign n8911 = ~n8729 & n8730;
  assign n8912 = n8859 ^ n8856;
  assign n8913 = ~n8911 & n8912;
  assign n8914 = n8862 ^ n8854;
  assign n8915 = n8913 & n8914;
  assign n8916 = n8865 ^ n8852;
  assign n8917 = ~n8915 & ~n8916;
  assign n8918 = n8868 ^ n8849;
  assign n8919 = n8917 & n8918;
  assign n8920 = n8871 ^ n8846;
  assign n8921 = ~n8919 & n8920;
  assign n8922 = n8874 ^ n6297;
  assign n8923 = n8922 ^ n8842;
  assign n8924 = n8921 & n8923;
  assign n8925 = ~n8910 & ~n8924;
  assign n8926 = n8909 & n8925;
  assign n8927 = n8908 & n8926;
  assign n8836 = n8835 ^ n6277;
  assign n8884 = n8883 ^ n8835;
  assign n8885 = ~n8836 & n8884;
  assign n8886 = n8885 ^ n6277;
  assign n8752 = n8751 ^ n8748;
  assign n8823 = n8822 ^ n8748;
  assign n8824 = n8752 & ~n8823;
  assign n8825 = n8824 ^ n8751;
  assign n8743 = n7833 ^ n7011;
  assign n8744 = ~n7811 & n8743;
  assign n8745 = n8744 ^ n7011;
  assign n8742 = n8506 ^ n8465;
  assign n8746 = n8745 ^ n8742;
  assign n8832 = n8825 ^ n8746;
  assign n8833 = n8832 ^ n6269;
  assign n8906 = n8886 ^ n8833;
  assign n9003 = n8927 ^ n8906;
  assign n9004 = n9003 ^ x369;
  assign n9005 = n8926 ^ n8908;
  assign n9006 = n9005 ^ x370;
  assign n9007 = n8925 ^ n8909;
  assign n9008 = n9007 ^ x371;
  assign n9009 = n8924 ^ n8910;
  assign n9010 = n9009 ^ x372;
  assign n9011 = n8923 ^ n8921;
  assign n9012 = n9011 ^ x373;
  assign n9013 = n8920 ^ n8919;
  assign n9014 = n9013 ^ x374;
  assign n9015 = n8918 ^ n8917;
  assign n9016 = n9015 ^ x375;
  assign n9017 = n8916 ^ n8915;
  assign n9018 = n9017 ^ x376;
  assign n9019 = n8914 ^ n8913;
  assign n9020 = n9019 ^ x377;
  assign n9021 = n8912 ^ n8911;
  assign n9022 = n9021 ^ x378;
  assign n8731 = n8730 ^ n8729;
  assign n8732 = n8731 ^ x379;
  assign n8677 = n8676 ^ n8670;
  assign n8678 = n8677 ^ x380;
  assign n8679 = n8675 ^ n8672;
  assign n8680 = n8679 ^ x381;
  assign n8681 = x383 & n8673;
  assign n8682 = n8681 ^ x382;
  assign n8683 = n8674 ^ n8673;
  assign n8684 = n8683 ^ n8681;
  assign n8685 = n8682 & ~n8684;
  assign n8686 = n8685 ^ x382;
  assign n8687 = n8686 ^ n8679;
  assign n8688 = ~n8680 & n8687;
  assign n8689 = n8688 ^ x381;
  assign n8690 = n8689 ^ n8677;
  assign n8691 = ~n8678 & n8690;
  assign n8692 = n8691 ^ x380;
  assign n9023 = n8731 ^ n8692;
  assign n9024 = n8732 & ~n9023;
  assign n9025 = n9024 ^ x379;
  assign n9026 = n9025 ^ n9021;
  assign n9027 = ~n9022 & n9026;
  assign n9028 = n9027 ^ x378;
  assign n9029 = n9028 ^ n9019;
  assign n9030 = n9020 & ~n9029;
  assign n9031 = n9030 ^ x377;
  assign n9032 = n9031 ^ n9017;
  assign n9033 = ~n9018 & n9032;
  assign n9034 = n9033 ^ x376;
  assign n9035 = n9034 ^ n9015;
  assign n9036 = ~n9016 & n9035;
  assign n9037 = n9036 ^ x375;
  assign n9038 = n9037 ^ n9013;
  assign n9039 = ~n9014 & n9038;
  assign n9040 = n9039 ^ x374;
  assign n9041 = n9040 ^ n9011;
  assign n9042 = n9012 & ~n9041;
  assign n9043 = n9042 ^ x373;
  assign n9044 = n9043 ^ n9009;
  assign n9045 = ~n9010 & n9044;
  assign n9046 = n9045 ^ x372;
  assign n9047 = n9046 ^ n9007;
  assign n9048 = ~n9008 & n9047;
  assign n9049 = n9048 ^ x371;
  assign n9050 = n9049 ^ n9005;
  assign n9051 = ~n9006 & n9050;
  assign n9052 = n9051 ^ x370;
  assign n9053 = n9052 ^ n9003;
  assign n9054 = ~n9004 & n9053;
  assign n9055 = n9054 ^ x369;
  assign n9124 = n9055 ^ x368;
  assign n8887 = n8886 ^ n8832;
  assign n8888 = ~n8833 & n8887;
  assign n8889 = n8888 ^ n6269;
  assign n8826 = n8825 ^ n8742;
  assign n8827 = n8746 & n8826;
  assign n8828 = n8827 ^ n8745;
  assign n8739 = n7827 ^ n7028;
  assign n8740 = n7805 & n8739;
  assign n8741 = n8740 ^ n7028;
  assign n8829 = n8828 ^ n8741;
  assign n8738 = n8509 ^ n8463;
  assign n8830 = n8829 ^ n8738;
  assign n8831 = n8830 ^ n5710;
  assign n8929 = n8889 ^ n8831;
  assign n8928 = n8906 & n8927;
  assign n9001 = n8929 ^ n8928;
  assign n9125 = n9124 ^ n9001;
  assign n9130 = n9129 ^ n9125;
  assign n9132 = n8538 ^ x332;
  assign n9133 = n9132 ^ n8446;
  assign n9134 = n8221 ^ n7799;
  assign n9135 = ~n9133 & n9134;
  assign n9136 = n9135 ^ n7799;
  assign n9131 = n9052 ^ n9004;
  assign n9137 = n9136 ^ n9131;
  assign n9142 = n9049 ^ x370;
  assign n9143 = n9142 ^ n9005;
  assign n9138 = n8535 ^ n8449;
  assign n9139 = n7806 ^ n7769;
  assign n9140 = ~n9138 & ~n9139;
  assign n9141 = n9140 ^ n7806;
  assign n9144 = n9143 ^ n9141;
  assign n9150 = n9046 ^ n9008;
  assign n9145 = n8532 ^ x334;
  assign n9146 = n9145 ^ n8450;
  assign n9147 = n7813 ^ n7777;
  assign n9148 = n9146 & ~n9147;
  assign n9149 = n9148 ^ n7813;
  assign n9151 = n9150 ^ n9149;
  assign n9155 = n9043 ^ x372;
  assign n9156 = n9155 ^ n9009;
  assign n9087 = n8529 ^ x335;
  assign n9152 = n7820 ^ n7783;
  assign n9153 = ~n9087 & ~n9152;
  assign n9154 = n9153 ^ n7820;
  assign n9157 = n9156 ^ n9154;
  assign n9161 = n9040 ^ n9012;
  assign n8988 = n8524 ^ x336;
  assign n8989 = n8988 ^ n8452;
  assign n9158 = n7827 ^ n7791;
  assign n9159 = n8989 & n9158;
  assign n9160 = n9159 ^ n7827;
  assign n9162 = n9161 ^ n9160;
  assign n9166 = n9037 ^ n9014;
  assign n8972 = n8521 ^ n8455;
  assign n9163 = n7833 ^ n7797;
  assign n9164 = ~n8972 & ~n9163;
  assign n9165 = n9164 ^ n7833;
  assign n9167 = n9166 ^ n9165;
  assign n9171 = n9034 ^ x375;
  assign n9172 = n9171 ^ n9015;
  assign n8956 = n8518 ^ x338;
  assign n8957 = n8956 ^ n8456;
  assign n9168 = n7805 ^ n7756;
  assign n9169 = ~n8957 & ~n9168;
  assign n9170 = n9169 ^ n7756;
  assign n9173 = n9172 ^ n9170;
  assign n9177 = n9031 ^ x376;
  assign n9178 = n9177 ^ n9017;
  assign n8941 = n8515 ^ n8459;
  assign n9174 = n7811 ^ n7650;
  assign n9175 = n8941 & ~n9174;
  assign n9176 = n9175 ^ n7650;
  assign n9179 = n9178 ^ n9176;
  assign n8900 = n8512 ^ x340;
  assign n8901 = n8900 ^ n8460;
  assign n9181 = n7819 ^ n7594;
  assign n9182 = n8901 & n9181;
  assign n9183 = n9182 ^ n7594;
  assign n9180 = n9028 ^ n9020;
  assign n9184 = n9183 ^ n9180;
  assign n9188 = n9025 ^ x378;
  assign n9189 = n9188 ^ n9021;
  assign n9185 = n7825 ^ n7495;
  assign n9186 = n8738 & ~n9185;
  assign n9187 = n9186 ^ n7495;
  assign n9190 = n9189 ^ n9187;
  assign n9191 = n7832 ^ n7302;
  assign n9192 = n8742 & ~n9191;
  assign n9193 = n9192 ^ n7302;
  assign n8733 = n8732 ^ n8692;
  assign n9194 = n9193 ^ n8733;
  assign n9198 = n8689 ^ x380;
  assign n9199 = n9198 ^ n8677;
  assign n9195 = n7838 ^ n7307;
  assign n9196 = ~n8748 & n9195;
  assign n9197 = n9196 ^ n7307;
  assign n9200 = n9199 ^ n9197;
  assign n9202 = n7847 ^ n7312;
  assign n9203 = ~n8754 & ~n9202;
  assign n9204 = n9203 ^ n7312;
  assign n9201 = n8686 ^ n8680;
  assign n9205 = n9204 ^ n9201;
  assign n9210 = n8673 ^ x383;
  assign n9207 = n7859 ^ n7321;
  assign n9208 = ~n8764 & ~n9207;
  assign n9209 = n9208 ^ n7321;
  assign n9211 = n9210 ^ n9209;
  assign n9410 = n7454 ^ n6340;
  assign n9411 = ~n8121 & ~n9410;
  assign n9412 = n9411 ^ n6340;
  assign n9095 = n8559 ^ n8433;
  assign n9413 = n9412 ^ n9095;
  assign n9414 = n9413 ^ n5731;
  assign n9218 = n7404 ^ n6720;
  assign n9219 = ~n8134 & ~n9218;
  assign n9220 = n9219 ^ n6720;
  assign n9116 = n8550 ^ x328;
  assign n9117 = n9116 ^ n8438;
  assign n9221 = n9220 ^ n9117;
  assign n9225 = n8547 ^ n8441;
  assign n9222 = n7414 ^ n6729;
  assign n9223 = n8140 & n9222;
  assign n9224 = n9223 ^ n6729;
  assign n9226 = n9225 ^ n9224;
  assign n9230 = n8544 ^ x330;
  assign n9231 = n9230 ^ n8442;
  assign n9227 = n7282 ^ n6731;
  assign n9228 = ~n8719 & n9227;
  assign n9229 = n9228 ^ n6731;
  assign n9232 = n9231 ^ n9229;
  assign n9233 = n7249 ^ n6740;
  assign n9234 = n8661 & n9233;
  assign n9235 = n9234 ^ n6740;
  assign n9236 = n9235 ^ n9126;
  assign n9237 = n7778 ^ n7371;
  assign n9238 = n8233 & ~n9237;
  assign n9239 = n9238 ^ n7371;
  assign n9240 = n9239 ^ n9146;
  assign n8984 = n7792 ^ n7245;
  assign n8985 = ~n7769 & ~n8984;
  assign n8986 = n8985 ^ n7245;
  assign n9083 = n8989 ^ n8986;
  assign n8969 = n7799 ^ n7096;
  assign n8970 = ~n7777 & n8969;
  assign n8971 = n8970 ^ n7096;
  assign n8973 = n8972 ^ n8971;
  assign n8953 = n7806 ^ n7078;
  assign n8954 = ~n7783 & n8953;
  assign n8955 = n8954 ^ n7078;
  assign n8958 = n8957 ^ n8955;
  assign n8938 = n7813 ^ n7061;
  assign n8939 = ~n7791 & n8938;
  assign n8940 = n8939 ^ n7061;
  assign n8942 = n8941 ^ n8940;
  assign n8897 = n7820 ^ n7045;
  assign n8898 = ~n7797 & n8897;
  assign n8899 = n8898 ^ n7045;
  assign n8902 = n8901 ^ n8899;
  assign n8893 = n8741 ^ n8738;
  assign n8894 = n8828 ^ n8738;
  assign n8895 = ~n8893 & ~n8894;
  assign n8896 = n8895 ^ n8741;
  assign n8935 = n8901 ^ n8896;
  assign n8936 = n8902 & n8935;
  assign n8937 = n8936 ^ n8899;
  assign n8950 = n8941 ^ n8937;
  assign n8951 = n8942 & ~n8950;
  assign n8952 = n8951 ^ n8940;
  assign n8966 = n8957 ^ n8952;
  assign n8967 = ~n8958 & n8966;
  assign n8968 = n8967 ^ n8955;
  assign n8981 = n8972 ^ n8968;
  assign n8982 = n8973 & n8981;
  assign n8983 = n8982 ^ n8971;
  assign n9084 = n8989 ^ n8983;
  assign n9085 = n9083 & n9084;
  assign n9086 = n9085 ^ n8986;
  assign n9088 = n9087 ^ n9086;
  assign n9080 = n7785 ^ n7278;
  assign n9081 = ~n8221 & ~n9080;
  assign n9082 = n9081 ^ n7278;
  assign n9241 = n9087 ^ n9082;
  assign n9242 = n9088 & n9241;
  assign n9243 = n9242 ^ n9082;
  assign n9244 = n9243 ^ n9239;
  assign n9245 = ~n9240 & ~n9244;
  assign n9246 = n9245 ^ n9146;
  assign n9247 = n9246 ^ n9138;
  assign n9248 = n7771 ^ n7398;
  assign n9249 = ~n8580 & n9248;
  assign n9250 = n9249 ^ n7398;
  assign n9251 = n9250 ^ n9138;
  assign n9252 = n9247 & n9251;
  assign n9253 = n9252 ^ n9250;
  assign n9254 = n9253 ^ n9133;
  assign n9255 = n8112 ^ n7441;
  assign n9256 = n8616 & n9255;
  assign n9257 = n9256 ^ n7441;
  assign n9258 = n9257 ^ n9253;
  assign n9259 = n9254 & n9258;
  assign n9260 = n9259 ^ n9133;
  assign n9261 = n9260 ^ n9126;
  assign n9262 = ~n9236 & ~n9261;
  assign n9263 = n9262 ^ n9235;
  assign n9264 = n9263 ^ n9231;
  assign n9265 = n9232 & ~n9264;
  assign n9266 = n9265 ^ n9229;
  assign n9267 = n9266 ^ n9225;
  assign n9268 = n9226 & ~n9267;
  assign n9269 = n9268 ^ n9224;
  assign n9270 = n9269 ^ n9117;
  assign n9271 = ~n9221 & n9270;
  assign n9272 = n9271 ^ n9220;
  assign n9110 = n8553 ^ n8437;
  assign n9273 = n9272 ^ n9110;
  assign n9215 = n7447 ^ n6777;
  assign n9216 = ~n8132 & ~n9215;
  assign n9217 = n9216 ^ n6777;
  assign n9326 = n9217 ^ n9110;
  assign n9327 = ~n9273 & ~n9326;
  assign n9328 = n9327 ^ n9217;
  assign n9102 = n8556 ^ x326;
  assign n9103 = n9102 ^ n8434;
  assign n9329 = n9328 ^ n9103;
  assign n9323 = n7351 ^ n6342;
  assign n9324 = n8127 & n9323;
  assign n9325 = n9324 ^ n6342;
  assign n9407 = n9325 ^ n9103;
  assign n9408 = n9329 & n9407;
  assign n9409 = n9408 ^ n9325;
  assign n9415 = n9414 ^ n9409;
  assign n9330 = n9329 ^ n9325;
  assign n9274 = n9273 ^ n9217;
  assign n9275 = n9274 ^ n6047;
  assign n9276 = n9269 ^ n9220;
  assign n9277 = n9276 ^ n9117;
  assign n9278 = n9277 ^ n6052;
  assign n9279 = n9266 ^ n9224;
  assign n9280 = n9279 ^ n9225;
  assign n9281 = n9280 ^ n6057;
  assign n9282 = n9263 ^ n9229;
  assign n9283 = n9282 ^ n9231;
  assign n9284 = n9283 ^ n6059;
  assign n9285 = n9260 ^ n9235;
  assign n9286 = n9285 ^ n9126;
  assign n9287 = n9286 ^ n6064;
  assign n9288 = n9257 ^ n9133;
  assign n9289 = n9288 ^ n9253;
  assign n9290 = n9289 ^ n6771;
  assign n9299 = n9250 ^ n9247;
  assign n9291 = n9243 ^ n9240;
  assign n9292 = n9291 ^ n6609;
  assign n9089 = n9088 ^ n9082;
  assign n9090 = n9089 ^ n6592;
  assign n8987 = n8986 ^ n8983;
  assign n8990 = n8989 ^ n8987;
  assign n8991 = n8990 ^ n6538;
  assign n8974 = n8973 ^ n8968;
  assign n8975 = n8974 ^ n6451;
  assign n8959 = n8958 ^ n8952;
  assign n8960 = n8959 ^ n6347;
  assign n8943 = n8942 ^ n8937;
  assign n8944 = n8943 ^ n6353;
  assign n8903 = n8902 ^ n8896;
  assign n8904 = n8903 ^ n6358;
  assign n8890 = n8889 ^ n8830;
  assign n8891 = n8831 & n8890;
  assign n8892 = n8891 ^ n5710;
  assign n8932 = n8903 ^ n8892;
  assign n8933 = n8904 & ~n8932;
  assign n8934 = n8933 ^ n6358;
  assign n8947 = n8943 ^ n8934;
  assign n8948 = ~n8944 & n8947;
  assign n8949 = n8948 ^ n6353;
  assign n8963 = n8959 ^ n8949;
  assign n8964 = n8960 & ~n8963;
  assign n8965 = n8964 ^ n6347;
  assign n8978 = n8974 ^ n8965;
  assign n8979 = ~n8975 & n8978;
  assign n8980 = n8979 ^ n6451;
  assign n9077 = n8990 ^ n8980;
  assign n9078 = n8991 & ~n9077;
  assign n9079 = n9078 ^ n6538;
  assign n9293 = n9089 ^ n9079;
  assign n9294 = n9090 & n9293;
  assign n9295 = n9294 ^ n6592;
  assign n9296 = n9295 ^ n9291;
  assign n9297 = n9292 & ~n9296;
  assign n9298 = n9297 ^ n6609;
  assign n9300 = n9299 ^ n9298;
  assign n9301 = n9299 ^ n6714;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = n9302 ^ n6714;
  assign n9304 = n9303 ^ n9289;
  assign n9305 = n9290 & n9304;
  assign n9306 = n9305 ^ n6771;
  assign n9307 = n9306 ^ n9286;
  assign n9308 = ~n9287 & ~n9307;
  assign n9309 = n9308 ^ n6064;
  assign n9310 = n9309 ^ n9283;
  assign n9311 = ~n9284 & n9310;
  assign n9312 = n9311 ^ n6059;
  assign n9313 = n9312 ^ n9280;
  assign n9314 = ~n9281 & n9313;
  assign n9315 = n9314 ^ n6057;
  assign n9316 = n9315 ^ n9277;
  assign n9317 = n9278 & ~n9316;
  assign n9318 = n9317 ^ n6052;
  assign n9319 = n9318 ^ n9274;
  assign n9320 = n9275 & ~n9319;
  assign n9321 = n9320 ^ n6047;
  assign n9322 = n9321 ^ n5739;
  assign n9331 = n9330 ^ n9322;
  assign n9332 = n9312 ^ n6057;
  assign n9333 = n9332 ^ n9280;
  assign n9334 = n9309 ^ n9284;
  assign n9335 = n9300 ^ n6714;
  assign n9091 = n9090 ^ n9079;
  assign n8905 = n8904 ^ n8892;
  assign n8930 = ~n8928 & n8929;
  assign n8931 = ~n8905 & n8930;
  assign n8945 = n8944 ^ n8934;
  assign n8946 = ~n8931 & ~n8945;
  assign n8961 = n8960 ^ n8949;
  assign n8962 = ~n8946 & ~n8961;
  assign n8976 = n8975 ^ n8965;
  assign n8977 = n8962 & n8976;
  assign n8992 = n8991 ^ n8980;
  assign n9092 = n8977 & ~n8992;
  assign n9336 = ~n9091 & n9092;
  assign n9337 = n9295 ^ n9292;
  assign n9338 = n9336 & n9337;
  assign n9339 = n9335 & ~n9338;
  assign n9340 = n9303 ^ n9290;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = n9306 ^ n9287;
  assign n9343 = ~n9341 & n9342;
  assign n9344 = n9334 & ~n9343;
  assign n9345 = ~n9333 & ~n9344;
  assign n9346 = n9315 ^ n6052;
  assign n9347 = n9346 ^ n9277;
  assign n9348 = n9345 & n9347;
  assign n9349 = n9318 ^ n6047;
  assign n9350 = n9349 ^ n9274;
  assign n9351 = ~n9348 & ~n9350;
  assign n9406 = ~n9331 & ~n9351;
  assign n9416 = n9415 ^ n9406;
  assign n9402 = n9330 ^ n5739;
  assign n9403 = n9330 ^ n9321;
  assign n9404 = ~n9402 & ~n9403;
  assign n9405 = n9404 ^ n5739;
  assign n9417 = n9416 ^ n9405;
  assign n9352 = n9351 ^ n9331;
  assign n9353 = n9352 ^ x353;
  assign n9354 = n9350 ^ n9348;
  assign n9355 = n9354 ^ x354;
  assign n9356 = n9347 ^ n9345;
  assign n9357 = n9356 ^ x355;
  assign n9358 = n9344 ^ n9333;
  assign n9359 = n9358 ^ x356;
  assign n9360 = n9343 ^ n9334;
  assign n9361 = n9360 ^ x357;
  assign n9362 = n9342 ^ n9341;
  assign n9363 = n9362 ^ x358;
  assign n9364 = n9340 ^ n9339;
  assign n9365 = n9364 ^ x359;
  assign n9366 = n9338 ^ n9335;
  assign n9367 = n9366 ^ x360;
  assign n9368 = n9337 ^ n9336;
  assign n9369 = n9368 ^ x361;
  assign n9093 = n9092 ^ n9091;
  assign n9370 = n9093 ^ x362;
  assign n8993 = n8992 ^ n8977;
  assign n8994 = n8993 ^ x363;
  assign n8995 = n8976 ^ n8962;
  assign n8996 = n8995 ^ x364;
  assign n8997 = n8961 ^ n8946;
  assign n8998 = n8997 ^ x365;
  assign n8999 = n8945 ^ n8931;
  assign n9000 = n8999 ^ x366;
  assign n9059 = n8930 ^ n8905;
  assign n9002 = n9001 ^ x368;
  assign n9056 = n9055 ^ n9001;
  assign n9057 = ~n9002 & n9056;
  assign n9058 = n9057 ^ x368;
  assign n9060 = n9059 ^ n9058;
  assign n9061 = n9059 ^ x367;
  assign n9062 = n9060 & ~n9061;
  assign n9063 = n9062 ^ x367;
  assign n9064 = n9063 ^ n8999;
  assign n9065 = ~n9000 & n9064;
  assign n9066 = n9065 ^ x366;
  assign n9067 = n9066 ^ n8997;
  assign n9068 = n8998 & ~n9067;
  assign n9069 = n9068 ^ x365;
  assign n9070 = n9069 ^ n8995;
  assign n9071 = n8996 & ~n9070;
  assign n9072 = n9071 ^ x364;
  assign n9073 = n9072 ^ n8993;
  assign n9074 = ~n8994 & n9073;
  assign n9075 = n9074 ^ x363;
  assign n9371 = n9093 ^ n9075;
  assign n9372 = ~n9370 & n9371;
  assign n9373 = n9372 ^ x362;
  assign n9374 = n9373 ^ n9368;
  assign n9375 = n9369 & ~n9374;
  assign n9376 = n9375 ^ x361;
  assign n9377 = n9376 ^ n9366;
  assign n9378 = n9367 & ~n9377;
  assign n9379 = n9378 ^ x360;
  assign n9380 = n9379 ^ n9364;
  assign n9381 = n9365 & ~n9380;
  assign n9382 = n9381 ^ x359;
  assign n9383 = n9382 ^ n9362;
  assign n9384 = n9363 & ~n9383;
  assign n9385 = n9384 ^ x358;
  assign n9386 = n9385 ^ n9360;
  assign n9387 = ~n9361 & n9386;
  assign n9388 = n9387 ^ x357;
  assign n9389 = n9388 ^ n9358;
  assign n9390 = ~n9359 & n9389;
  assign n9391 = n9390 ^ x356;
  assign n9392 = n9391 ^ n9356;
  assign n9393 = ~n9357 & n9392;
  assign n9394 = n9393 ^ x355;
  assign n9395 = n9394 ^ n9354;
  assign n9396 = n9355 & ~n9395;
  assign n9397 = n9396 ^ x354;
  assign n9398 = n9397 ^ n9352;
  assign n9399 = ~n9353 & n9398;
  assign n9400 = n9399 ^ x353;
  assign n9401 = n9400 ^ x352;
  assign n9418 = n9417 ^ n9401;
  assign n9212 = n7864 ^ n7326;
  assign n9213 = n8769 & n9212;
  assign n9214 = n9213 ^ n7326;
  assign n9419 = n9418 ^ n9214;
  assign n9423 = n9397 ^ x353;
  assign n9424 = n9423 ^ n9352;
  assign n9420 = n7870 ^ n7332;
  assign n9421 = ~n8775 & n9420;
  assign n9422 = n9421 ^ n7332;
  assign n9425 = n9424 ^ n9422;
  assign n9441 = n7875 ^ n7337;
  assign n9442 = ~n8784 & n9441;
  assign n9443 = n9442 ^ n7337;
  assign n9429 = n9391 ^ x355;
  assign n9430 = n9429 ^ n9356;
  assign n9426 = n7881 ^ n7294;
  assign n9427 = ~n8786 & ~n9426;
  assign n9428 = n9427 ^ n7294;
  assign n9431 = n9430 ^ n9428;
  assign n9432 = n7883 ^ n7346;
  assign n9433 = ~n8791 & n9432;
  assign n9434 = n9433 ^ n7346;
  assign n9435 = n9388 ^ x356;
  assign n9436 = n9435 ^ n9358;
  assign n9437 = ~n9434 & ~n9436;
  assign n9438 = n9437 ^ n9430;
  assign n9439 = n9431 & ~n9438;
  assign n9440 = n9439 ^ n9437;
  assign n9444 = n9443 ^ n9440;
  assign n9445 = n9394 ^ x354;
  assign n9446 = n9445 ^ n9354;
  assign n9447 = n9446 ^ n9440;
  assign n9448 = ~n9444 & ~n9447;
  assign n9449 = n9448 ^ n9443;
  assign n9450 = n9449 ^ n9424;
  assign n9451 = ~n9425 & ~n9450;
  assign n9452 = n9451 ^ n9422;
  assign n9453 = n9452 ^ n9418;
  assign n9454 = ~n9419 & ~n9453;
  assign n9455 = n9454 ^ n9214;
  assign n9456 = n9455 ^ n9210;
  assign n9457 = n9211 & n9456;
  assign n9458 = n9457 ^ n9209;
  assign n9206 = n8683 ^ n8682;
  assign n9459 = n9458 ^ n9206;
  assign n9460 = n7853 ^ n7315;
  assign n9461 = n8734 & n9460;
  assign n9462 = n9461 ^ n7315;
  assign n9463 = n9462 ^ n9206;
  assign n9464 = ~n9459 & n9463;
  assign n9465 = n9464 ^ n9462;
  assign n9466 = n9465 ^ n9201;
  assign n9467 = ~n9205 & n9466;
  assign n9468 = n9467 ^ n9204;
  assign n9469 = n9468 ^ n9199;
  assign n9470 = n9200 & n9469;
  assign n9471 = n9470 ^ n9197;
  assign n9472 = n9471 ^ n8733;
  assign n9473 = ~n9194 & n9472;
  assign n9474 = n9473 ^ n9193;
  assign n9475 = n9474 ^ n9189;
  assign n9476 = ~n9190 & ~n9475;
  assign n9477 = n9476 ^ n9187;
  assign n9478 = n9477 ^ n9180;
  assign n9479 = ~n9184 & ~n9478;
  assign n9480 = n9479 ^ n9183;
  assign n9481 = n9480 ^ n9178;
  assign n9482 = ~n9179 & ~n9481;
  assign n9483 = n9482 ^ n9176;
  assign n9484 = n9483 ^ n9172;
  assign n9485 = n9173 & n9484;
  assign n9486 = n9485 ^ n9170;
  assign n9487 = n9486 ^ n9166;
  assign n9488 = ~n9167 & ~n9487;
  assign n9489 = n9488 ^ n9165;
  assign n9490 = n9489 ^ n9161;
  assign n9491 = ~n9162 & ~n9490;
  assign n9492 = n9491 ^ n9160;
  assign n9493 = n9492 ^ n9156;
  assign n9494 = ~n9157 & ~n9493;
  assign n9495 = n9494 ^ n9154;
  assign n9496 = n9495 ^ n9150;
  assign n9497 = ~n9151 & n9496;
  assign n9498 = n9497 ^ n9149;
  assign n9499 = n9498 ^ n9143;
  assign n9500 = ~n9144 & n9499;
  assign n9501 = n9500 ^ n9141;
  assign n9502 = n9501 ^ n9131;
  assign n9503 = n9137 & n9502;
  assign n9504 = n9503 ^ n9136;
  assign n9505 = n9504 ^ n9125;
  assign n9506 = n9130 & ~n9505;
  assign n9507 = n9506 ^ n9129;
  assign n9123 = n9060 ^ x367;
  assign n9508 = n9507 ^ n9123;
  assign n9509 = n8580 ^ n7785;
  assign n9510 = n9231 & ~n9509;
  assign n9511 = n9510 ^ n7785;
  assign n9512 = n9511 ^ n9123;
  assign n9513 = ~n9508 & ~n9512;
  assign n9514 = n9513 ^ n9511;
  assign n9122 = n9063 ^ n9000;
  assign n9515 = n9514 ^ n9122;
  assign n9516 = n8616 ^ n7778;
  assign n9517 = n9225 & n9516;
  assign n9518 = n9517 ^ n7778;
  assign n9519 = n9518 ^ n9122;
  assign n9520 = n9515 & ~n9519;
  assign n9521 = n9520 ^ n9518;
  assign n9118 = n8661 ^ n7771;
  assign n9119 = ~n9117 & ~n9118;
  assign n9120 = n9119 ^ n7771;
  assign n9549 = n9521 ^ n9120;
  assign n9115 = n9066 ^ n8998;
  assign n9550 = n9549 ^ n9115;
  assign n9551 = n9550 ^ n7398;
  assign n9552 = n9518 ^ n9515;
  assign n9553 = n9552 ^ n7371;
  assign n9554 = n9511 ^ n9508;
  assign n9555 = n9554 ^ n7278;
  assign n9556 = n9504 ^ n9130;
  assign n9557 = n9556 ^ n7245;
  assign n9558 = n9501 ^ n9136;
  assign n9559 = n9558 ^ n9131;
  assign n9560 = n9559 ^ n7096;
  assign n9561 = n9498 ^ n9141;
  assign n9562 = n9561 ^ n9143;
  assign n9563 = n9562 ^ n7078;
  assign n9564 = n9495 ^ n9149;
  assign n9565 = n9564 ^ n9150;
  assign n9566 = n9565 ^ n7061;
  assign n9567 = n9492 ^ n9157;
  assign n9568 = n9567 ^ n7045;
  assign n9569 = n9489 ^ n9160;
  assign n9570 = n9569 ^ n9161;
  assign n9571 = n9570 ^ n7028;
  assign n9572 = n9486 ^ n9167;
  assign n9573 = n9572 ^ n7011;
  assign n9574 = n9483 ^ n9170;
  assign n9575 = n9574 ^ n9172;
  assign n9576 = n9575 ^ n6996;
  assign n9577 = n9480 ^ n9179;
  assign n9578 = n9577 ^ n6933;
  assign n9579 = n9477 ^ n9183;
  assign n9580 = n9579 ^ n9180;
  assign n9581 = n9580 ^ n6824;
  assign n9582 = n9474 ^ n9190;
  assign n9583 = n9582 ^ n6267;
  assign n9584 = n9471 ^ n9193;
  assign n9585 = n9584 ^ n8733;
  assign n9586 = n9585 ^ n6274;
  assign n9587 = n9468 ^ n9200;
  assign n9588 = n9587 ^ n6281;
  assign n9589 = n9465 ^ n9204;
  assign n9590 = n9589 ^ n9201;
  assign n9591 = n9590 ^ n6287;
  assign n9592 = n9462 ^ n9459;
  assign n9593 = n9592 ^ n6290;
  assign n9594 = n9455 ^ n9209;
  assign n9595 = n9594 ^ n9210;
  assign n9596 = n9595 ^ n6302;
  assign n9597 = n9452 ^ n9214;
  assign n9598 = n9597 ^ n9418;
  assign n9599 = n9598 ^ n6304;
  assign n9600 = n9449 ^ n9425;
  assign n9601 = n9600 ^ n6316;
  assign n9602 = n9446 ^ n9444;
  assign n9603 = n9602 ^ n6318;
  assign n9604 = n9436 ^ n9434;
  assign n9605 = ~n6335 & n9604;
  assign n9606 = n9605 ^ n6330;
  assign n9607 = n9437 ^ n9428;
  assign n9608 = n9607 ^ n9430;
  assign n9609 = n9608 ^ n9605;
  assign n9610 = ~n9606 & n9609;
  assign n9611 = n9610 ^ n6330;
  assign n9612 = n9611 ^ n9602;
  assign n9613 = ~n9603 & ~n9612;
  assign n9614 = n9613 ^ n6318;
  assign n9615 = n9614 ^ n9600;
  assign n9616 = n9601 & ~n9615;
  assign n9617 = n9616 ^ n6316;
  assign n9618 = n9617 ^ n9598;
  assign n9619 = n9599 & n9618;
  assign n9620 = n9619 ^ n6304;
  assign n9621 = n9620 ^ n9595;
  assign n9622 = ~n9596 & ~n9621;
  assign n9623 = n9622 ^ n6302;
  assign n9624 = n9623 ^ n9592;
  assign n9625 = ~n9593 & ~n9624;
  assign n9626 = n9625 ^ n6290;
  assign n9627 = n9626 ^ n9590;
  assign n9628 = ~n9591 & ~n9627;
  assign n9629 = n9628 ^ n6287;
  assign n9630 = n9629 ^ n9587;
  assign n9631 = n9588 & ~n9630;
  assign n9632 = n9631 ^ n6281;
  assign n9633 = n9632 ^ n9585;
  assign n9634 = n9586 & ~n9633;
  assign n9635 = n9634 ^ n6274;
  assign n9636 = n9635 ^ n9582;
  assign n9637 = n9583 & ~n9636;
  assign n9638 = n9637 ^ n6267;
  assign n9639 = n9638 ^ n9580;
  assign n9640 = ~n9581 & n9639;
  assign n9641 = n9640 ^ n6824;
  assign n9642 = n9641 ^ n9577;
  assign n9643 = ~n9578 & ~n9642;
  assign n9644 = n9643 ^ n6933;
  assign n9645 = n9644 ^ n9575;
  assign n9646 = ~n9576 & n9645;
  assign n9647 = n9646 ^ n6996;
  assign n9648 = n9647 ^ n9572;
  assign n9649 = n9573 & n9648;
  assign n9650 = n9649 ^ n7011;
  assign n9651 = n9650 ^ n9570;
  assign n9652 = n9571 & n9651;
  assign n9653 = n9652 ^ n7028;
  assign n9654 = n9653 ^ n9567;
  assign n9655 = n9568 & n9654;
  assign n9656 = n9655 ^ n7045;
  assign n9657 = n9656 ^ n9565;
  assign n9658 = ~n9566 & n9657;
  assign n9659 = n9658 ^ n7061;
  assign n9660 = n9659 ^ n9562;
  assign n9661 = ~n9563 & n9660;
  assign n9662 = n9661 ^ n7078;
  assign n9663 = n9662 ^ n9559;
  assign n9664 = ~n9560 & ~n9663;
  assign n9665 = n9664 ^ n7096;
  assign n9666 = n9665 ^ n9556;
  assign n9667 = ~n9557 & ~n9666;
  assign n9668 = n9667 ^ n7245;
  assign n9669 = n9668 ^ n9554;
  assign n9670 = ~n9555 & ~n9669;
  assign n9671 = n9670 ^ n7278;
  assign n9672 = n9671 ^ n9552;
  assign n9673 = n9553 & ~n9672;
  assign n9674 = n9673 ^ n7371;
  assign n9675 = n9674 ^ n9550;
  assign n9676 = n9551 & ~n9675;
  assign n9677 = n9676 ^ n7398;
  assign n9121 = n9120 ^ n9115;
  assign n9522 = n9521 ^ n9115;
  assign n9523 = ~n9121 & ~n9522;
  assign n9524 = n9523 ^ n9120;
  assign n9111 = n8719 ^ n8112;
  assign n9112 = n9110 & ~n9111;
  assign n9113 = n9112 ^ n8112;
  assign n9108 = n9069 ^ x364;
  assign n9109 = n9108 ^ n8995;
  assign n9114 = n9113 ^ n9109;
  assign n9547 = n9524 ^ n9114;
  assign n9548 = n9547 ^ n7441;
  assign n9706 = n9677 ^ n9548;
  assign n9707 = n9671 ^ n9553;
  assign n9708 = n9668 ^ n9555;
  assign n9709 = n9665 ^ n9557;
  assign n9710 = n9656 ^ n9566;
  assign n9711 = n9653 ^ n9568;
  assign n9712 = n9650 ^ n9571;
  assign n9713 = n9644 ^ n9576;
  assign n9714 = n9635 ^ n9583;
  assign n9715 = n9632 ^ n6274;
  assign n9716 = n9715 ^ n9585;
  assign n9717 = n9629 ^ n9588;
  assign n9718 = n9611 ^ n6318;
  assign n9719 = n9718 ^ n9602;
  assign n9720 = n9604 ^ n6335;
  assign n9721 = n9608 ^ n9606;
  assign n9722 = ~n9720 & n9721;
  assign n9723 = n9719 & n9722;
  assign n9724 = n9614 ^ n6316;
  assign n9725 = n9724 ^ n9600;
  assign n9726 = ~n9723 & ~n9725;
  assign n9727 = n9617 ^ n6304;
  assign n9728 = n9727 ^ n9598;
  assign n9729 = n9726 & ~n9728;
  assign n9730 = n9620 ^ n6302;
  assign n9731 = n9730 ^ n9595;
  assign n9732 = ~n9729 & n9731;
  assign n9733 = n9623 ^ n6290;
  assign n9734 = n9733 ^ n9592;
  assign n9735 = n9732 & ~n9734;
  assign n9736 = n9626 ^ n9591;
  assign n9737 = ~n9735 & ~n9736;
  assign n9738 = ~n9717 & n9737;
  assign n9739 = n9716 & ~n9738;
  assign n9740 = n9714 & n9739;
  assign n9741 = n9638 ^ n9581;
  assign n9742 = ~n9740 & n9741;
  assign n9743 = n9641 ^ n9578;
  assign n9744 = n9742 & n9743;
  assign n9745 = ~n9713 & n9744;
  assign n9746 = n9647 ^ n9573;
  assign n9747 = n9745 & n9746;
  assign n9748 = n9712 & ~n9747;
  assign n9749 = ~n9711 & n9748;
  assign n9750 = n9710 & ~n9749;
  assign n9751 = n9659 ^ n9563;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = n9662 ^ n7096;
  assign n9754 = n9753 ^ n9559;
  assign n9755 = n9752 & ~n9754;
  assign n9756 = n9709 & n9755;
  assign n9757 = ~n9708 & n9756;
  assign n9758 = ~n9707 & n9757;
  assign n9759 = n9674 ^ n7398;
  assign n9760 = n9759 ^ n9550;
  assign n9761 = ~n9758 & n9760;
  assign n9762 = n9706 & ~n9761;
  assign n9678 = n9677 ^ n9547;
  assign n9679 = ~n9548 & ~n9678;
  assign n9680 = n9679 ^ n7441;
  assign n9525 = n9524 ^ n9109;
  assign n9526 = n9114 & n9525;
  assign n9527 = n9526 ^ n9113;
  assign n9104 = n8140 ^ n7249;
  assign n9105 = n9103 & n9104;
  assign n9106 = n9105 ^ n7249;
  assign n9544 = n9527 ^ n9106;
  assign n9100 = n9072 ^ x363;
  assign n9101 = n9100 ^ n8993;
  assign n9545 = n9544 ^ n9101;
  assign n9546 = n9545 ^ n6740;
  assign n9763 = n9680 ^ n9546;
  assign n9764 = ~n9762 & n9763;
  assign n9681 = n9680 ^ n9545;
  assign n9682 = ~n9546 & n9681;
  assign n9683 = n9682 ^ n6740;
  assign n9107 = n9106 ^ n9101;
  assign n9528 = n9527 ^ n9101;
  assign n9529 = ~n9107 & n9528;
  assign n9530 = n9529 ^ n9106;
  assign n9096 = n8134 ^ n7282;
  assign n9097 = ~n9095 & ~n9096;
  assign n9098 = n9097 ^ n7282;
  assign n9541 = n9530 ^ n9098;
  assign n9076 = n9075 ^ x362;
  assign n9094 = n9093 ^ n9076;
  assign n9542 = n9541 ^ n9094;
  assign n9543 = n9542 ^ n6731;
  assign n9705 = n9683 ^ n9543;
  assign n9808 = n9764 ^ n9705;
  assign n9809 = n9808 ^ x389;
  assign n9810 = n9763 ^ n9762;
  assign n9811 = n9810 ^ x390;
  assign n9928 = n9761 ^ n9706;
  assign n9812 = n9760 ^ n9758;
  assign n9813 = n9812 ^ x392;
  assign n9814 = n9757 ^ n9707;
  assign n9815 = n9814 ^ x393;
  assign n9816 = n9756 ^ n9708;
  assign n9817 = n9816 ^ x394;
  assign n9818 = n9755 ^ n9709;
  assign n9819 = n9818 ^ x395;
  assign n9820 = n9754 ^ n9752;
  assign n9821 = n9820 ^ x396;
  assign n9822 = n9751 ^ n9750;
  assign n9823 = n9822 ^ x397;
  assign n9824 = n9749 ^ n9710;
  assign n9825 = n9824 ^ x398;
  assign n9902 = n9748 ^ n9711;
  assign n9826 = n9747 ^ n9712;
  assign n9827 = n9826 ^ x400;
  assign n9828 = n9746 ^ n9745;
  assign n9829 = n9828 ^ x401;
  assign n9830 = n9744 ^ n9713;
  assign n9831 = n9830 ^ x402;
  assign n9832 = n9743 ^ n9742;
  assign n9833 = n9832 ^ x403;
  assign n9834 = n9741 ^ n9740;
  assign n9835 = n9834 ^ x404;
  assign n9836 = n9739 ^ n9714;
  assign n9837 = n9836 ^ x405;
  assign n9838 = n9738 ^ n9716;
  assign n9839 = n9838 ^ x406;
  assign n9840 = n9737 ^ n9717;
  assign n9841 = n9840 ^ x407;
  assign n9842 = n9736 ^ n9735;
  assign n9843 = n9842 ^ x408;
  assign n9844 = n9734 ^ n9732;
  assign n9845 = n9844 ^ x409;
  assign n9846 = n9731 ^ n9729;
  assign n9847 = n9846 ^ x410;
  assign n9848 = n9728 ^ n9726;
  assign n9849 = n9848 ^ x411;
  assign n9850 = n9725 ^ n9723;
  assign n9851 = n9850 ^ x412;
  assign n9852 = n9722 ^ n9719;
  assign n9853 = n9852 ^ x413;
  assign n9854 = x415 & n9720;
  assign n9855 = n9854 ^ x414;
  assign n9856 = n9721 ^ n9720;
  assign n9857 = n9856 ^ n9854;
  assign n9858 = n9855 & n9857;
  assign n9859 = n9858 ^ x414;
  assign n9860 = n9859 ^ n9852;
  assign n9861 = n9853 & ~n9860;
  assign n9862 = n9861 ^ x413;
  assign n9863 = n9862 ^ n9850;
  assign n9864 = ~n9851 & n9863;
  assign n9865 = n9864 ^ x412;
  assign n9866 = n9865 ^ n9848;
  assign n9867 = n9849 & ~n9866;
  assign n9868 = n9867 ^ x411;
  assign n9869 = n9868 ^ n9846;
  assign n9870 = ~n9847 & n9869;
  assign n9871 = n9870 ^ x410;
  assign n9872 = n9871 ^ n9844;
  assign n9873 = ~n9845 & n9872;
  assign n9874 = n9873 ^ x409;
  assign n9875 = n9874 ^ n9842;
  assign n9876 = ~n9843 & n9875;
  assign n9877 = n9876 ^ x408;
  assign n9878 = n9877 ^ n9840;
  assign n9879 = n9841 & ~n9878;
  assign n9880 = n9879 ^ x407;
  assign n9881 = n9880 ^ n9838;
  assign n9882 = ~n9839 & n9881;
  assign n9883 = n9882 ^ x406;
  assign n9884 = n9883 ^ n9836;
  assign n9885 = n9837 & ~n9884;
  assign n9886 = n9885 ^ x405;
  assign n9887 = n9886 ^ n9834;
  assign n9888 = n9835 & ~n9887;
  assign n9889 = n9888 ^ x404;
  assign n9890 = n9889 ^ n9832;
  assign n9891 = ~n9833 & n9890;
  assign n9892 = n9891 ^ x403;
  assign n9893 = n9892 ^ n9830;
  assign n9894 = n9831 & ~n9893;
  assign n9895 = n9894 ^ x402;
  assign n9896 = n9895 ^ n9828;
  assign n9897 = ~n9829 & n9896;
  assign n9898 = n9897 ^ x401;
  assign n9899 = n9898 ^ n9826;
  assign n9900 = ~n9827 & n9899;
  assign n9901 = n9900 ^ x400;
  assign n9903 = n9902 ^ n9901;
  assign n9904 = n9902 ^ x399;
  assign n9905 = n9903 & ~n9904;
  assign n9906 = n9905 ^ x399;
  assign n9907 = n9906 ^ n9824;
  assign n9908 = n9825 & ~n9907;
  assign n9909 = n9908 ^ x398;
  assign n9910 = n9909 ^ n9822;
  assign n9911 = n9823 & ~n9910;
  assign n9912 = n9911 ^ x397;
  assign n9913 = n9912 ^ n9820;
  assign n9914 = ~n9821 & n9913;
  assign n9915 = n9914 ^ x396;
  assign n9916 = n9915 ^ n9818;
  assign n9917 = n9819 & ~n9916;
  assign n9918 = n9917 ^ x395;
  assign n9919 = n9918 ^ n9816;
  assign n9920 = ~n9817 & n9919;
  assign n9921 = n9920 ^ x394;
  assign n9922 = n9921 ^ n9814;
  assign n9923 = ~n9815 & n9922;
  assign n9924 = n9923 ^ x393;
  assign n9925 = n9924 ^ n9812;
  assign n9926 = n9813 & ~n9925;
  assign n9927 = n9926 ^ x392;
  assign n9929 = n9928 ^ n9927;
  assign n9930 = n9928 ^ x391;
  assign n9931 = n9929 & ~n9930;
  assign n9932 = n9931 ^ x391;
  assign n9933 = n9932 ^ n9810;
  assign n9934 = n9811 & ~n9933;
  assign n9935 = n9934 ^ x390;
  assign n9936 = n9935 ^ n9808;
  assign n9937 = n9809 & ~n9936;
  assign n9938 = n9937 ^ x389;
  assign n9986 = n9938 ^ x388;
  assign n9765 = ~n9705 & ~n9764;
  assign n9684 = n9683 ^ n9542;
  assign n9685 = ~n9543 & n9684;
  assign n9686 = n9685 ^ n6731;
  assign n9703 = n9686 ^ n6729;
  assign n9538 = n9373 ^ n9369;
  assign n9534 = n8132 ^ n7414;
  assign n9535 = ~n8589 & ~n9534;
  assign n9536 = n9535 ^ n7414;
  assign n9099 = n9098 ^ n9094;
  assign n9531 = n9530 ^ n9094;
  assign n9532 = ~n9099 & n9531;
  assign n9533 = n9532 ^ n9098;
  assign n9537 = n9536 ^ n9533;
  assign n9539 = n9538 ^ n9537;
  assign n9704 = n9703 ^ n9539;
  assign n9806 = n9765 ^ n9704;
  assign n9987 = n9986 ^ n9806;
  assign n9983 = n8784 ^ n7883;
  assign n9984 = n9210 & n9983;
  assign n9985 = n9984 ^ n7883;
  assign n10022 = n9987 ^ n9985;
  assign n10058 = n10022 ^ n7346;
  assign n10817 = n10058 ^ x447;
  assign n10105 = n9859 ^ n9853;
  assign n11308 = n10105 ^ n9201;
  assign n11309 = n10817 & ~n11308;
  assign n11310 = n11309 ^ n9201;
  assign n10388 = n9918 ^ x394;
  assign n10389 = n10388 ^ n9816;
  assign n9699 = n9376 ^ x360;
  assign n9700 = n9699 ^ n9366;
  assign n10736 = n9700 ^ n9117;
  assign n10737 = ~n10389 & ~n10736;
  assign n10738 = n10737 ^ n9117;
  assign n10205 = n8989 ^ n7805;
  assign n10206 = ~n9143 & n10205;
  assign n10207 = n10206 ^ n7805;
  assign n10204 = n9877 ^ n9841;
  assign n10208 = n10207 ^ n10204;
  assign n10211 = n8972 ^ n7811;
  assign n10212 = ~n9150 & n10211;
  assign n10213 = n10212 ^ n7811;
  assign n10209 = n9874 ^ x408;
  assign n10210 = n10209 ^ n9842;
  assign n10214 = n10213 ^ n10210;
  assign n10217 = n8957 ^ n7819;
  assign n10218 = ~n9156 & n10217;
  assign n10219 = n10218 ^ n7819;
  assign n10215 = n9871 ^ x409;
  assign n10216 = n10215 ^ n9844;
  assign n10220 = n10219 ^ n10216;
  assign n10223 = n8941 ^ n7825;
  assign n10224 = n9161 & ~n10223;
  assign n10225 = n10224 ^ n7825;
  assign n10221 = n9868 ^ x410;
  assign n10222 = n10221 ^ n9846;
  assign n10226 = n10225 ^ n10222;
  assign n10228 = n8901 ^ n7832;
  assign n10229 = ~n9166 & n10228;
  assign n10230 = n10229 ^ n7832;
  assign n10227 = n9865 ^ n9849;
  assign n10231 = n10230 ^ n10227;
  assign n10131 = n9862 ^ x412;
  assign n10132 = n10131 ^ n9850;
  assign n10128 = n8738 ^ n7838;
  assign n10129 = ~n9172 & ~n10128;
  assign n10130 = n10129 ^ n7838;
  assign n10133 = n10132 ^ n10130;
  assign n10047 = n8748 ^ n7853;
  assign n10048 = n9180 & ~n10047;
  assign n10049 = n10048 ^ n7853;
  assign n10046 = n9856 ^ n9855;
  assign n10050 = n10049 ^ n10046;
  assign n10011 = n9720 ^ x415;
  assign n10007 = n8754 ^ n7859;
  assign n10008 = ~n9189 & n10007;
  assign n10009 = n10008 ^ n7859;
  assign n10042 = n10011 ^ n10009;
  assign n9963 = n9385 ^ n9361;
  assign n9960 = n7454 ^ n7292;
  assign n9961 = ~n8725 & n9960;
  assign n9962 = n9961 ^ n7454;
  assign n9964 = n9963 ^ n9962;
  assign n9965 = n9964 ^ n6340;
  assign n9796 = n9382 ^ n9363;
  assign n9793 = n7892 ^ n7351;
  assign n9794 = n8667 & n9793;
  assign n9795 = n9794 ^ n7351;
  assign n9797 = n9796 ^ n9795;
  assign n9695 = n8127 ^ n7404;
  assign n9696 = n8586 & ~n9695;
  assign n9697 = n9696 ^ n7404;
  assign n9777 = n9700 ^ n9697;
  assign n9691 = n9538 ^ n9536;
  assign n9692 = n9538 ^ n9533;
  assign n9693 = n9691 & ~n9692;
  assign n9694 = n9693 ^ n9536;
  assign n9778 = n9700 ^ n9694;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = n9779 ^ n9697;
  assign n9776 = n9379 ^ n9365;
  assign n9781 = n9780 ^ n9776;
  assign n9773 = n8121 ^ n7447;
  assign n9774 = ~n8622 & ~n9773;
  assign n9775 = n9774 ^ n7447;
  assign n9790 = n9776 ^ n9775;
  assign n9791 = n9781 & n9790;
  assign n9792 = n9791 ^ n9775;
  assign n9957 = n9796 ^ n9792;
  assign n9958 = n9797 & ~n9957;
  assign n9959 = n9958 ^ n9795;
  assign n9966 = n9965 ^ n9959;
  assign n9698 = n9697 ^ n9694;
  assign n9701 = n9700 ^ n9698;
  assign n9540 = n9539 ^ n6729;
  assign n9687 = n9686 ^ n9539;
  assign n9688 = n9540 & ~n9687;
  assign n9689 = n9688 ^ n6729;
  assign n9690 = n9689 ^ n6720;
  assign n9702 = n9701 ^ n9690;
  assign n9766 = ~n9704 & ~n9765;
  assign n9767 = n9702 & n9766;
  assign n9782 = n9781 ^ n9775;
  assign n9768 = n9701 ^ n6720;
  assign n9769 = n9701 ^ n9689;
  assign n9770 = ~n9768 & n9769;
  assign n9771 = n9770 ^ n6720;
  assign n9772 = n9771 ^ n6777;
  assign n9783 = n9782 ^ n9772;
  assign n9784 = ~n9767 & n9783;
  assign n9798 = n9797 ^ n9792;
  assign n9785 = n9782 ^ n6777;
  assign n9786 = n9782 ^ n9771;
  assign n9787 = n9785 & n9786;
  assign n9788 = n9787 ^ n6777;
  assign n9789 = n9788 ^ n6342;
  assign n9799 = n9798 ^ n9789;
  assign n9956 = ~n9784 & n9799;
  assign n9967 = n9966 ^ n9956;
  assign n9952 = n9798 ^ n6342;
  assign n9953 = n9798 ^ n9788;
  assign n9954 = n9952 & n9953;
  assign n9955 = n9954 ^ n6342;
  assign n9968 = n9967 ^ n9955;
  assign n9800 = n9799 ^ n9784;
  assign n9801 = n9800 ^ x385;
  assign n9802 = n9783 ^ n9767;
  assign n9803 = n9802 ^ x386;
  assign n9804 = n9766 ^ n9702;
  assign n9805 = n9804 ^ x387;
  assign n9807 = n9806 ^ x388;
  assign n9939 = n9938 ^ n9806;
  assign n9940 = ~n9807 & n9939;
  assign n9941 = n9940 ^ x388;
  assign n9942 = n9941 ^ n9804;
  assign n9943 = ~n9805 & n9942;
  assign n9944 = n9943 ^ x387;
  assign n9945 = n9944 ^ n9802;
  assign n9946 = ~n9803 & n9945;
  assign n9947 = n9946 ^ x386;
  assign n9948 = n9947 ^ n9800;
  assign n9949 = n9801 & ~n9948;
  assign n9950 = n9949 ^ x385;
  assign n9951 = n9950 ^ x384;
  assign n9969 = n9968 ^ n9951;
  assign n8735 = n8734 ^ n7864;
  assign n8736 = n8733 & ~n8735;
  assign n8737 = n8736 ^ n7864;
  assign n9970 = n9969 ^ n8737;
  assign n9974 = n9947 ^ x385;
  assign n9975 = n9974 ^ n9800;
  assign n9971 = n8764 ^ n7870;
  assign n9972 = ~n9199 & ~n9971;
  assign n9973 = n9972 ^ n7870;
  assign n9976 = n9975 ^ n9973;
  assign n9992 = n8769 ^ n7875;
  assign n9993 = ~n9201 & ~n9992;
  assign n9994 = n9993 ^ n7875;
  assign n9980 = n9941 ^ x387;
  assign n9981 = n9980 ^ n9804;
  assign n9977 = n8775 ^ n7881;
  assign n9978 = n9206 & n9977;
  assign n9979 = n9978 ^ n7881;
  assign n9982 = n9981 ^ n9979;
  assign n9988 = ~n9985 & ~n9987;
  assign n9989 = n9988 ^ n9981;
  assign n9990 = ~n9982 & ~n9989;
  assign n9991 = n9990 ^ n9988;
  assign n9995 = n9994 ^ n9991;
  assign n9996 = n9944 ^ x386;
  assign n9997 = n9996 ^ n9802;
  assign n9998 = n9997 ^ n9991;
  assign n9999 = ~n9995 & n9998;
  assign n10000 = n9999 ^ n9994;
  assign n10001 = n10000 ^ n9975;
  assign n10002 = n9976 & n10001;
  assign n10003 = n10002 ^ n9973;
  assign n10004 = n10003 ^ n9969;
  assign n10005 = n9970 & n10004;
  assign n10006 = n10005 ^ n8737;
  assign n10043 = n10011 ^ n10006;
  assign n10044 = ~n10042 & n10043;
  assign n10045 = n10044 ^ n10009;
  assign n10107 = n10046 ^ n10045;
  assign n10108 = ~n10050 & ~n10107;
  assign n10109 = n10108 ^ n10049;
  assign n10124 = n10109 ^ n10105;
  assign n10102 = n8742 ^ n7847;
  assign n10103 = ~n9178 & ~n10102;
  assign n10104 = n10103 ^ n7847;
  assign n10125 = n10109 ^ n10104;
  assign n10126 = n10124 & n10125;
  assign n10127 = n10126 ^ n10105;
  assign n10232 = n10132 ^ n10127;
  assign n10233 = n10133 & n10232;
  assign n10234 = n10233 ^ n10130;
  assign n10235 = n10234 ^ n10227;
  assign n10236 = n10231 & n10235;
  assign n10237 = n10236 ^ n10230;
  assign n10238 = n10237 ^ n10222;
  assign n10239 = n10226 & n10238;
  assign n10240 = n10239 ^ n10225;
  assign n10241 = n10240 ^ n10216;
  assign n10242 = n10220 & ~n10241;
  assign n10243 = n10242 ^ n10219;
  assign n10244 = n10243 ^ n10210;
  assign n10245 = n10214 & ~n10244;
  assign n10246 = n10245 ^ n10213;
  assign n10247 = n10246 ^ n10204;
  assign n10248 = n10208 & n10247;
  assign n10249 = n10248 ^ n10207;
  assign n10200 = n9087 ^ n7797;
  assign n10201 = ~n9131 & n10200;
  assign n10202 = n10201 ^ n7797;
  assign n10199 = n9880 ^ n9839;
  assign n10203 = n10202 ^ n10199;
  assign n10315 = n10249 ^ n10203;
  assign n10316 = n10315 ^ n7833;
  assign n10317 = n10246 ^ n10208;
  assign n10318 = n10317 ^ n7756;
  assign n10319 = n10243 ^ n10214;
  assign n10320 = n10319 ^ n7650;
  assign n10321 = n10240 ^ n10220;
  assign n10322 = n10321 ^ n7594;
  assign n10323 = n10237 ^ n10226;
  assign n10324 = n10323 ^ n7495;
  assign n10325 = n10234 ^ n10231;
  assign n10326 = n10325 ^ n7302;
  assign n10134 = n10133 ^ n10127;
  assign n10135 = n10134 ^ n7307;
  assign n10051 = n10050 ^ n10045;
  assign n10052 = n10051 ^ n7315;
  assign n10010 = n10009 ^ n10006;
  assign n10012 = n10011 ^ n10010;
  assign n10013 = n10012 ^ n7321;
  assign n10014 = n10003 ^ n8737;
  assign n10015 = n10014 ^ n9969;
  assign n10016 = n10015 ^ n7326;
  assign n10017 = n10000 ^ n9973;
  assign n10018 = n10017 ^ n9975;
  assign n10019 = n10018 ^ n7332;
  assign n10020 = n9997 ^ n9995;
  assign n10021 = n10020 ^ n7337;
  assign n10023 = ~n7346 & n10022;
  assign n10024 = n10023 ^ n7294;
  assign n10025 = n9988 ^ n9979;
  assign n10026 = n10025 ^ n9981;
  assign n10027 = n10026 ^ n10023;
  assign n10028 = n10024 & ~n10027;
  assign n10029 = n10028 ^ n7294;
  assign n10030 = n10029 ^ n10020;
  assign n10031 = ~n10021 & ~n10030;
  assign n10032 = n10031 ^ n7337;
  assign n10033 = n10032 ^ n10018;
  assign n10034 = ~n10019 & ~n10033;
  assign n10035 = n10034 ^ n7332;
  assign n10036 = n10035 ^ n10015;
  assign n10037 = ~n10016 & ~n10036;
  assign n10038 = n10037 ^ n7326;
  assign n10039 = n10038 ^ n10012;
  assign n10040 = n10013 & n10039;
  assign n10041 = n10040 ^ n7321;
  assign n10112 = n10051 ^ n10041;
  assign n10113 = n10052 & ~n10112;
  assign n10114 = n10113 ^ n7315;
  assign n10120 = n10114 ^ n7312;
  assign n10106 = n10105 ^ n10104;
  assign n10110 = n10109 ^ n10106;
  assign n10121 = n10114 ^ n10110;
  assign n10122 = n10120 & n10121;
  assign n10123 = n10122 ^ n7312;
  assign n10327 = n10134 ^ n10123;
  assign n10328 = ~n10135 & ~n10327;
  assign n10329 = n10328 ^ n7307;
  assign n10330 = n10329 ^ n10325;
  assign n10331 = n10326 & ~n10330;
  assign n10332 = n10331 ^ n7302;
  assign n10333 = n10332 ^ n10323;
  assign n10334 = n10324 & n10333;
  assign n10335 = n10334 ^ n7495;
  assign n10336 = n10335 ^ n10321;
  assign n10337 = n10322 & n10336;
  assign n10338 = n10337 ^ n7594;
  assign n10339 = n10338 ^ n10319;
  assign n10340 = ~n10320 & ~n10339;
  assign n10341 = n10340 ^ n7650;
  assign n10342 = n10341 ^ n10317;
  assign n10343 = n10318 & n10342;
  assign n10344 = n10343 ^ n7756;
  assign n10345 = n10344 ^ n10315;
  assign n10346 = n10316 & n10345;
  assign n10347 = n10346 ^ n7833;
  assign n10250 = n10249 ^ n10199;
  assign n10251 = n10203 & n10250;
  assign n10252 = n10251 ^ n10202;
  assign n10195 = n9146 ^ n7791;
  assign n10196 = ~n9125 & ~n10195;
  assign n10197 = n10196 ^ n7791;
  assign n10141 = n9883 ^ n9837;
  assign n10198 = n10197 ^ n10141;
  assign n10313 = n10252 ^ n10198;
  assign n10314 = n10313 ^ n7827;
  assign n10401 = n10347 ^ n10314;
  assign n10402 = n10344 ^ n10316;
  assign n10136 = n10135 ^ n10123;
  assign n10053 = n10052 ^ n10041;
  assign n10054 = n10038 ^ n7321;
  assign n10055 = n10054 ^ n10012;
  assign n10056 = n10032 ^ n7332;
  assign n10057 = n10056 ^ n10018;
  assign n10059 = n10026 ^ n10024;
  assign n10060 = ~n10058 & n10059;
  assign n10061 = n10029 ^ n7337;
  assign n10062 = n10061 ^ n10020;
  assign n10063 = n10060 & ~n10062;
  assign n10064 = ~n10057 & ~n10063;
  assign n10065 = n10035 ^ n7326;
  assign n10066 = n10065 ^ n10015;
  assign n10067 = n10064 & n10066;
  assign n10068 = ~n10055 & ~n10067;
  assign n10101 = n10053 & n10068;
  assign n10111 = n10110 ^ n7312;
  assign n10115 = n10114 ^ n10111;
  assign n10137 = ~n10101 & n10115;
  assign n10403 = n10136 & n10137;
  assign n10404 = n10329 ^ n10326;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = n10332 ^ n10324;
  assign n10407 = n10405 & ~n10406;
  assign n10408 = n10335 ^ n10322;
  assign n10409 = ~n10407 & ~n10408;
  assign n10410 = n10338 ^ n10320;
  assign n10411 = n10409 & ~n10410;
  assign n10412 = n10341 ^ n10318;
  assign n10413 = n10411 & ~n10412;
  assign n10414 = n10402 & n10413;
  assign n10415 = ~n10401 & ~n10414;
  assign n10348 = n10347 ^ n10313;
  assign n10349 = ~n10314 & ~n10348;
  assign n10350 = n10349 ^ n7827;
  assign n10253 = n10252 ^ n10141;
  assign n10254 = ~n10198 & n10253;
  assign n10255 = n10254 ^ n10197;
  assign n10191 = n9138 ^ n7783;
  assign n10192 = ~n9123 & n10191;
  assign n10193 = n10192 ^ n7783;
  assign n10310 = n10255 ^ n10193;
  assign n10189 = n9886 ^ x404;
  assign n10190 = n10189 ^ n9834;
  assign n10311 = n10310 ^ n10190;
  assign n10312 = n10311 ^ n7820;
  assign n10400 = n10350 ^ n10312;
  assign n10488 = n10415 ^ n10400;
  assign n10450 = n10414 ^ n10401;
  assign n10451 = n10450 ^ x432;
  assign n10452 = n10413 ^ n10402;
  assign n10453 = n10452 ^ x433;
  assign n10454 = n10412 ^ n10411;
  assign n10455 = n10454 ^ x434;
  assign n10456 = n10410 ^ n10409;
  assign n10457 = n10456 ^ x435;
  assign n10458 = n10408 ^ n10407;
  assign n10459 = n10458 ^ x436;
  assign n10460 = n10406 ^ n10405;
  assign n10461 = n10460 ^ x437;
  assign n10462 = n10404 ^ n10403;
  assign n10463 = n10462 ^ x438;
  assign n10138 = n10137 ^ n10136;
  assign n10139 = n10138 ^ x439;
  assign n10069 = n10068 ^ n10053;
  assign n10070 = n10069 ^ x441;
  assign n10071 = n10067 ^ n10055;
  assign n10072 = n10071 ^ x442;
  assign n10073 = n10066 ^ n10064;
  assign n10074 = n10073 ^ x443;
  assign n10075 = n10063 ^ n10057;
  assign n10076 = n10075 ^ x444;
  assign n10077 = n10062 ^ n10060;
  assign n10078 = n10077 ^ x445;
  assign n10079 = x447 & n10058;
  assign n10080 = n10079 ^ x446;
  assign n10081 = n10059 ^ n10058;
  assign n10082 = n10081 ^ n10079;
  assign n10083 = n10080 & n10082;
  assign n10084 = n10083 ^ x446;
  assign n10085 = n10084 ^ n10077;
  assign n10086 = ~n10078 & n10085;
  assign n10087 = n10086 ^ x445;
  assign n10088 = n10087 ^ n10075;
  assign n10089 = ~n10076 & n10088;
  assign n10090 = n10089 ^ x444;
  assign n10091 = n10090 ^ n10073;
  assign n10092 = ~n10074 & n10091;
  assign n10093 = n10092 ^ x443;
  assign n10094 = n10093 ^ n10071;
  assign n10095 = n10072 & ~n10094;
  assign n10096 = n10095 ^ x442;
  assign n10097 = n10096 ^ n10069;
  assign n10098 = n10070 & ~n10097;
  assign n10099 = n10098 ^ x441;
  assign n10100 = n10099 ^ x440;
  assign n10116 = n10115 ^ n10101;
  assign n10117 = n10116 ^ n10099;
  assign n10118 = n10100 & ~n10117;
  assign n10119 = n10118 ^ x440;
  assign n10464 = n10138 ^ n10119;
  assign n10465 = ~n10139 & n10464;
  assign n10466 = n10465 ^ x439;
  assign n10467 = n10466 ^ n10462;
  assign n10468 = n10463 & ~n10467;
  assign n10469 = n10468 ^ x438;
  assign n10470 = n10469 ^ n10460;
  assign n10471 = ~n10461 & n10470;
  assign n10472 = n10471 ^ x437;
  assign n10473 = n10472 ^ n10458;
  assign n10474 = ~n10459 & n10473;
  assign n10475 = n10474 ^ x436;
  assign n10476 = n10475 ^ n10456;
  assign n10477 = n10457 & ~n10476;
  assign n10478 = n10477 ^ x435;
  assign n10479 = n10478 ^ n10454;
  assign n10480 = n10455 & ~n10479;
  assign n10481 = n10480 ^ x434;
  assign n10482 = n10481 ^ n10452;
  assign n10483 = ~n10453 & n10482;
  assign n10484 = n10483 ^ x433;
  assign n10485 = n10484 ^ n10450;
  assign n10486 = n10451 & ~n10485;
  assign n10487 = n10486 ^ x432;
  assign n10489 = n10488 ^ n10487;
  assign n10735 = n10489 ^ x431;
  assign n10739 = n10738 ^ n10735;
  assign n10289 = n9915 ^ n9819;
  assign n10742 = n9538 ^ n9225;
  assign n10743 = n10289 & n10742;
  assign n10744 = n10743 ^ n9225;
  assign n10740 = n10484 ^ x432;
  assign n10741 = n10740 ^ n10450;
  assign n10745 = n10744 ^ n10741;
  assign n10154 = n9912 ^ x396;
  assign n10155 = n10154 ^ n9820;
  assign n10747 = n9231 ^ n9094;
  assign n10748 = ~n10155 & ~n10747;
  assign n10749 = n10748 ^ n9231;
  assign n10746 = n10481 ^ n10453;
  assign n10750 = n10749 ^ n10746;
  assign n10160 = n9909 ^ n9823;
  assign n10753 = n9126 ^ n9101;
  assign n10754 = n10160 & n10753;
  assign n10755 = n10754 ^ n9126;
  assign n10751 = n10478 ^ x434;
  assign n10752 = n10751 ^ n10454;
  assign n10756 = n10755 ^ n10752;
  assign n10274 = n9906 ^ x398;
  assign n10275 = n10274 ^ n9824;
  assign n10758 = n9133 ^ n9109;
  assign n10759 = n10275 & ~n10758;
  assign n10760 = n10759 ^ n9133;
  assign n10757 = n10475 ^ n10457;
  assign n10761 = n10760 ^ n10757;
  assign n10165 = n9903 ^ x399;
  assign n10764 = n9138 ^ n9115;
  assign n10765 = ~n10165 & ~n10764;
  assign n10766 = n10765 ^ n9138;
  assign n10762 = n10472 ^ x436;
  assign n10763 = n10762 ^ n10458;
  assign n10767 = n10766 ^ n10763;
  assign n10170 = n9898 ^ x400;
  assign n10171 = n10170 ^ n9826;
  assign n10769 = n9146 ^ n9122;
  assign n10770 = ~n10171 & ~n10769;
  assign n10771 = n10770 ^ n9146;
  assign n10768 = n10469 ^ n10461;
  assign n10772 = n10771 ^ n10768;
  assign n10776 = n10466 ^ n10463;
  assign n10176 = n9895 ^ n9829;
  assign n10773 = n9123 ^ n9087;
  assign n10774 = ~n10176 & n10773;
  assign n10775 = n10774 ^ n9087;
  assign n10777 = n10776 ^ n10775;
  assign n10181 = n9892 ^ x402;
  assign n10182 = n10181 ^ n9830;
  assign n10778 = n9125 ^ n8989;
  assign n10779 = n10182 & ~n10778;
  assign n10780 = n10779 ^ n8989;
  assign n10140 = n10139 ^ n10119;
  assign n10781 = n10780 ^ n10140;
  assign n10187 = n9889 ^ n9833;
  assign n10782 = n9131 ^ n8972;
  assign n10783 = ~n10187 & n10782;
  assign n10784 = n10783 ^ n8972;
  assign n10672 = n10116 ^ n10100;
  assign n10785 = n10784 ^ n10672;
  assign n10786 = n9143 ^ n8957;
  assign n10787 = n10190 & n10786;
  assign n10788 = n10787 ^ n8957;
  assign n10679 = n10096 ^ n10070;
  assign n10789 = n10788 ^ n10679;
  assign n10790 = n9150 ^ n8941;
  assign n10791 = n10141 & ~n10790;
  assign n10792 = n10791 ^ n8941;
  assign n10685 = n10093 ^ x442;
  assign n10686 = n10685 ^ n10071;
  assign n10793 = n10792 ^ n10686;
  assign n10794 = n9156 ^ n8901;
  assign n10795 = ~n10199 & ~n10794;
  assign n10796 = n10795 ^ n8901;
  assign n10691 = n10090 ^ n10074;
  assign n10797 = n10796 ^ n10691;
  assign n10801 = n10087 ^ x444;
  assign n10802 = n10801 ^ n10075;
  assign n10798 = n9161 ^ n8738;
  assign n10799 = n10204 & n10798;
  assign n10800 = n10799 ^ n8738;
  assign n10803 = n10802 ^ n10800;
  assign n10805 = n9166 ^ n8742;
  assign n10806 = ~n10210 & ~n10805;
  assign n10807 = n10806 ^ n8742;
  assign n10804 = n10084 ^ n10078;
  assign n10808 = n10807 ^ n10804;
  assign n10810 = n9172 ^ n8748;
  assign n10811 = ~n10216 & n10810;
  assign n10812 = n10811 ^ n8748;
  assign n10809 = n10081 ^ n10080;
  assign n10813 = n10812 ^ n10809;
  assign n10814 = n9178 ^ n8754;
  assign n10815 = ~n10222 & n10814;
  assign n10816 = n10815 ^ n8754;
  assign n10818 = n10817 ^ n10816;
  assign n10841 = n9180 ^ n8734;
  assign n10842 = n10227 & n10841;
  assign n10843 = n10842 ^ n8734;
  assign n10832 = n8786 ^ n7292;
  assign n10833 = n9418 & n10832;
  assign n10834 = n10833 ^ n7292;
  assign n10712 = n9935 ^ n9809;
  assign n10835 = n10834 ^ n10712;
  assign n10836 = n10835 ^ n7454;
  assign n10602 = n9929 ^ x391;
  assign n10568 = n9924 ^ x392;
  assign n10569 = n10568 ^ n9812;
  assign n10564 = n8667 ^ n8127;
  assign n10565 = ~n9430 & n10564;
  assign n10566 = n10565 ^ n8127;
  assign n10598 = n10569 ^ n10566;
  assign n10536 = n9921 ^ x393;
  assign n10537 = n10536 ^ n9814;
  assign n10532 = n8622 ^ n8132;
  assign n10533 = ~n9436 & n10532;
  assign n10534 = n10533 ^ n8132;
  assign n10560 = n10537 ^ n10534;
  assign n10384 = n8586 ^ n8134;
  assign n10385 = ~n9963 & ~n10384;
  assign n10386 = n10385 ^ n8134;
  assign n10528 = n10389 ^ n10386;
  assign n10151 = n9095 ^ n8719;
  assign n10152 = n9776 & n10151;
  assign n10153 = n10152 ^ n8719;
  assign n10156 = n10155 ^ n10153;
  assign n10157 = n9103 ^ n8661;
  assign n10158 = n9700 & n10157;
  assign n10159 = n10158 ^ n8661;
  assign n10161 = n10160 ^ n10159;
  assign n10162 = n9117 ^ n8580;
  assign n10163 = ~n9094 & n10162;
  assign n10164 = n10163 ^ n8580;
  assign n10166 = n10165 ^ n10164;
  assign n10167 = n9225 ^ n8233;
  assign n10168 = ~n9101 & n10167;
  assign n10169 = n10168 ^ n8233;
  assign n10172 = n10171 ^ n10169;
  assign n10173 = n9231 ^ n8221;
  assign n10174 = n9109 & ~n10173;
  assign n10175 = n10174 ^ n8221;
  assign n10177 = n10176 ^ n10175;
  assign n10178 = n9126 ^ n7769;
  assign n10179 = n9115 & n10178;
  assign n10180 = n10179 ^ n7769;
  assign n10183 = n10182 ^ n10180;
  assign n10184 = n9133 ^ n7777;
  assign n10185 = ~n9122 & n10184;
  assign n10186 = n10185 ^ n7777;
  assign n10188 = n10187 ^ n10186;
  assign n10194 = n10193 ^ n10190;
  assign n10256 = n10255 ^ n10190;
  assign n10257 = ~n10194 & n10256;
  assign n10258 = n10257 ^ n10193;
  assign n10259 = n10258 ^ n10187;
  assign n10260 = n10188 & ~n10259;
  assign n10261 = n10260 ^ n10186;
  assign n10262 = n10261 ^ n10182;
  assign n10263 = ~n10183 & n10262;
  assign n10264 = n10263 ^ n10180;
  assign n10265 = n10264 ^ n10176;
  assign n10266 = n10177 & ~n10265;
  assign n10267 = n10266 ^ n10175;
  assign n10268 = n10267 ^ n10171;
  assign n10269 = ~n10172 & ~n10268;
  assign n10270 = n10269 ^ n10169;
  assign n10271 = n10270 ^ n10165;
  assign n10272 = n10166 & n10271;
  assign n10273 = n10272 ^ n10164;
  assign n10276 = n10275 ^ n10273;
  assign n10277 = n9110 ^ n8616;
  assign n10278 = n9538 & n10277;
  assign n10279 = n10278 ^ n8616;
  assign n10280 = n10279 ^ n10275;
  assign n10281 = n10276 & n10280;
  assign n10282 = n10281 ^ n10279;
  assign n10283 = n10282 ^ n10160;
  assign n10284 = n10161 & ~n10283;
  assign n10285 = n10284 ^ n10159;
  assign n10286 = n10285 ^ n10155;
  assign n10287 = n10156 & n10286;
  assign n10288 = n10287 ^ n10153;
  assign n10290 = n10289 ^ n10288;
  assign n10148 = n8589 ^ n8140;
  assign n10149 = n9796 & ~n10148;
  assign n10150 = n10149 ^ n8140;
  assign n10381 = n10289 ^ n10150;
  assign n10382 = n10290 & n10381;
  assign n10383 = n10382 ^ n10150;
  assign n10529 = n10389 ^ n10383;
  assign n10530 = n10528 & n10529;
  assign n10531 = n10530 ^ n10386;
  assign n10561 = n10537 ^ n10531;
  assign n10562 = n10560 & ~n10561;
  assign n10563 = n10562 ^ n10534;
  assign n10599 = n10569 ^ n10563;
  assign n10600 = n10598 & n10599;
  assign n10601 = n10600 ^ n10566;
  assign n10603 = n10602 ^ n10601;
  assign n10595 = n8725 ^ n8121;
  assign n10596 = n9446 & n10595;
  assign n10597 = n10596 ^ n8121;
  assign n10657 = n10602 ^ n10597;
  assign n10658 = n10603 & n10657;
  assign n10659 = n10658 ^ n10597;
  assign n10655 = n9932 ^ x390;
  assign n10656 = n10655 ^ n9810;
  assign n10660 = n10659 ^ n10656;
  assign n10652 = n8791 ^ n7892;
  assign n10653 = ~n9424 & ~n10652;
  assign n10654 = n10653 ^ n7892;
  assign n10829 = n10656 ^ n10654;
  assign n10830 = n10660 & n10829;
  assign n10831 = n10830 ^ n10654;
  assign n10837 = n10836 ^ n10831;
  assign n10661 = n10660 ^ n10654;
  assign n10604 = n10603 ^ n10597;
  assign n10647 = n10604 ^ n7447;
  assign n10567 = n10566 ^ n10563;
  assign n10570 = n10569 ^ n10567;
  assign n10590 = n10570 ^ n7404;
  assign n10535 = n10534 ^ n10531;
  assign n10538 = n10537 ^ n10535;
  assign n10555 = n10538 ^ n7414;
  assign n10387 = n10386 ^ n10383;
  assign n10390 = n10389 ^ n10387;
  assign n10391 = n10390 ^ n7282;
  assign n10291 = n10290 ^ n10150;
  assign n10292 = n10291 ^ n7249;
  assign n10293 = n10285 ^ n10156;
  assign n10294 = n10293 ^ n8112;
  assign n10295 = n10282 ^ n10159;
  assign n10296 = n10295 ^ n10160;
  assign n10297 = n10296 ^ n7771;
  assign n10298 = n10279 ^ n10276;
  assign n10299 = n10298 ^ n7778;
  assign n10300 = n10270 ^ n10166;
  assign n10301 = n10300 ^ n7785;
  assign n10302 = n10267 ^ n10172;
  assign n10303 = n10302 ^ n7792;
  assign n10304 = n10264 ^ n10177;
  assign n10305 = n10304 ^ n7799;
  assign n10306 = n10261 ^ n10183;
  assign n10307 = n10306 ^ n7806;
  assign n10308 = n10258 ^ n10188;
  assign n10309 = n10308 ^ n7813;
  assign n10351 = n10350 ^ n10311;
  assign n10352 = n10312 & n10351;
  assign n10353 = n10352 ^ n7820;
  assign n10354 = n10353 ^ n10308;
  assign n10355 = ~n10309 & n10354;
  assign n10356 = n10355 ^ n7813;
  assign n10357 = n10356 ^ n10306;
  assign n10358 = n10307 & ~n10357;
  assign n10359 = n10358 ^ n7806;
  assign n10360 = n10359 ^ n10304;
  assign n10361 = n10305 & n10360;
  assign n10362 = n10361 ^ n7799;
  assign n10363 = n10362 ^ n10302;
  assign n10364 = ~n10303 & n10363;
  assign n10365 = n10364 ^ n7792;
  assign n10366 = n10365 ^ n10300;
  assign n10367 = n10301 & n10366;
  assign n10368 = n10367 ^ n7785;
  assign n10369 = n10368 ^ n10298;
  assign n10370 = ~n10299 & n10369;
  assign n10371 = n10370 ^ n7778;
  assign n10372 = n10371 ^ n10296;
  assign n10373 = ~n10297 & ~n10372;
  assign n10374 = n10373 ^ n7771;
  assign n10375 = n10374 ^ n10293;
  assign n10376 = n10294 & n10375;
  assign n10377 = n10376 ^ n8112;
  assign n10378 = n10377 ^ n10291;
  assign n10379 = ~n10292 & n10378;
  assign n10380 = n10379 ^ n7249;
  assign n10524 = n10390 ^ n10380;
  assign n10525 = n10391 & ~n10524;
  assign n10526 = n10525 ^ n7282;
  assign n10556 = n10538 ^ n10526;
  assign n10557 = ~n10555 & n10556;
  assign n10558 = n10557 ^ n7414;
  assign n10591 = n10570 ^ n10558;
  assign n10592 = n10590 & n10591;
  assign n10593 = n10592 ^ n7404;
  assign n10648 = n10604 ^ n10593;
  assign n10649 = n10647 & n10648;
  assign n10650 = n10649 ^ n7447;
  assign n10651 = n10650 ^ n7351;
  assign n10662 = n10661 ^ n10651;
  assign n10559 = n10558 ^ n7404;
  assign n10571 = n10570 ^ n10559;
  assign n10527 = n10526 ^ n7414;
  assign n10539 = n10538 ^ n10527;
  assign n10392 = n10391 ^ n10380;
  assign n10393 = n10377 ^ n10292;
  assign n10394 = n10374 ^ n10294;
  assign n10395 = n10368 ^ n10299;
  assign n10396 = n10365 ^ n10301;
  assign n10397 = n10362 ^ n10303;
  assign n10398 = n10359 ^ n7799;
  assign n10399 = n10398 ^ n10304;
  assign n10416 = ~n10400 & n10415;
  assign n10417 = n10353 ^ n10309;
  assign n10418 = ~n10416 & n10417;
  assign n10419 = n10356 ^ n10307;
  assign n10420 = ~n10418 & n10419;
  assign n10421 = n10399 & n10420;
  assign n10422 = n10397 & n10421;
  assign n10423 = ~n10396 & n10422;
  assign n10424 = ~n10395 & n10423;
  assign n10425 = n10371 ^ n7771;
  assign n10426 = n10425 ^ n10296;
  assign n10427 = ~n10424 & n10426;
  assign n10428 = ~n10394 & ~n10427;
  assign n10429 = n10393 & ~n10428;
  assign n10540 = n10392 & ~n10429;
  assign n10572 = n10539 & ~n10540;
  assign n10589 = ~n10571 & n10572;
  assign n10594 = n10593 ^ n7447;
  assign n10605 = n10604 ^ n10594;
  assign n10663 = ~n10589 & ~n10605;
  assign n10828 = n10662 & ~n10663;
  assign n10838 = n10837 ^ n10828;
  assign n10824 = n10661 ^ n7351;
  assign n10825 = n10661 ^ n10650;
  assign n10826 = ~n10824 & n10825;
  assign n10827 = n10826 ^ n7351;
  assign n10839 = n10838 ^ n10827;
  assign n10664 = n10663 ^ n10662;
  assign n10819 = n10664 ^ x417;
  assign n10606 = n10605 ^ n10589;
  assign n10642 = n10606 ^ x418;
  assign n10573 = n10572 ^ n10571;
  assign n10584 = n10573 ^ x419;
  assign n10541 = n10540 ^ n10539;
  assign n10550 = n10541 ^ x420;
  assign n10430 = n10429 ^ n10392;
  assign n10431 = n10430 ^ x421;
  assign n10432 = n10428 ^ n10393;
  assign n10433 = n10432 ^ x422;
  assign n10434 = n10427 ^ n10394;
  assign n10435 = n10434 ^ x423;
  assign n10436 = n10426 ^ n10424;
  assign n10437 = n10436 ^ x424;
  assign n10438 = n10423 ^ n10395;
  assign n10439 = n10438 ^ x425;
  assign n10440 = n10422 ^ n10396;
  assign n10441 = n10440 ^ x426;
  assign n10442 = n10421 ^ n10397;
  assign n10443 = n10442 ^ x427;
  assign n10444 = n10420 ^ n10399;
  assign n10445 = n10444 ^ x428;
  assign n10446 = n10419 ^ n10418;
  assign n10447 = n10446 ^ x429;
  assign n10448 = n10417 ^ n10416;
  assign n10449 = n10448 ^ x430;
  assign n10490 = n10488 ^ x431;
  assign n10491 = n10489 & ~n10490;
  assign n10492 = n10491 ^ x431;
  assign n10493 = n10492 ^ n10448;
  assign n10494 = n10449 & ~n10493;
  assign n10495 = n10494 ^ x430;
  assign n10496 = n10495 ^ n10446;
  assign n10497 = ~n10447 & n10496;
  assign n10498 = n10497 ^ x429;
  assign n10499 = n10498 ^ n10444;
  assign n10500 = n10445 & ~n10499;
  assign n10501 = n10500 ^ x428;
  assign n10502 = n10501 ^ n10442;
  assign n10503 = n10443 & ~n10502;
  assign n10504 = n10503 ^ x427;
  assign n10505 = n10504 ^ n10440;
  assign n10506 = ~n10441 & n10505;
  assign n10507 = n10506 ^ x426;
  assign n10508 = n10507 ^ n10438;
  assign n10509 = ~n10439 & n10508;
  assign n10510 = n10509 ^ x425;
  assign n10511 = n10510 ^ n10436;
  assign n10512 = n10437 & ~n10511;
  assign n10513 = n10512 ^ x424;
  assign n10514 = n10513 ^ n10434;
  assign n10515 = n10435 & ~n10514;
  assign n10516 = n10515 ^ x423;
  assign n10517 = n10516 ^ n10432;
  assign n10518 = n10433 & ~n10517;
  assign n10519 = n10518 ^ x422;
  assign n10520 = n10519 ^ n10430;
  assign n10521 = ~n10431 & n10520;
  assign n10522 = n10521 ^ x421;
  assign n10551 = n10541 ^ n10522;
  assign n10552 = n10550 & ~n10551;
  assign n10553 = n10552 ^ x420;
  assign n10585 = n10573 ^ n10553;
  assign n10586 = n10584 & ~n10585;
  assign n10587 = n10586 ^ x419;
  assign n10643 = n10606 ^ n10587;
  assign n10644 = n10642 & ~n10643;
  assign n10645 = n10644 ^ x418;
  assign n10820 = n10664 ^ n10645;
  assign n10821 = n10819 & ~n10820;
  assign n10822 = n10821 ^ x417;
  assign n10823 = n10822 ^ x416;
  assign n10840 = n10839 ^ n10823;
  assign n10844 = n10843 ^ n10840;
  assign n10646 = n10645 ^ x417;
  assign n10665 = n10664 ^ n10646;
  assign n10638 = n9189 ^ n8764;
  assign n10639 = ~n10132 & n10638;
  assign n10640 = n10639 ^ n8764;
  assign n10845 = n10665 ^ n10640;
  assign n10612 = n8769 ^ n8733;
  assign n10613 = n10105 & n10612;
  assign n10614 = n10613 ^ n8769;
  assign n10554 = n10553 ^ x419;
  assign n10574 = n10573 ^ n10554;
  assign n10546 = n9199 ^ n8775;
  assign n10547 = ~n10046 & n10546;
  assign n10548 = n10547 ^ n8775;
  assign n10608 = n10574 ^ n10548;
  assign n10145 = n9201 ^ n8784;
  assign n10146 = n10011 & n10145;
  assign n10147 = n10146 ^ n8784;
  assign n10523 = n10522 ^ x420;
  assign n10542 = n10541 ^ n10523;
  assign n10545 = ~n10147 & n10542;
  assign n10609 = n10574 ^ n10545;
  assign n10610 = n10608 & n10609;
  assign n10611 = n10610 ^ n10545;
  assign n10615 = n10614 ^ n10611;
  assign n10588 = n10587 ^ x418;
  assign n10607 = n10606 ^ n10588;
  assign n10635 = n10611 ^ n10607;
  assign n10636 = n10615 & ~n10635;
  assign n10637 = n10636 ^ n10614;
  assign n10846 = n10665 ^ n10637;
  assign n10847 = ~n10845 & ~n10846;
  assign n10848 = n10847 ^ n10640;
  assign n10849 = n10848 ^ n10840;
  assign n10850 = ~n10844 & ~n10849;
  assign n10851 = n10850 ^ n10843;
  assign n10852 = n10851 ^ n10817;
  assign n10853 = ~n10818 & ~n10852;
  assign n10854 = n10853 ^ n10816;
  assign n10855 = n10854 ^ n10809;
  assign n10856 = n10813 & ~n10855;
  assign n10857 = n10856 ^ n10812;
  assign n10858 = n10857 ^ n10804;
  assign n10859 = ~n10808 & ~n10858;
  assign n10860 = n10859 ^ n10807;
  assign n10861 = n10860 ^ n10802;
  assign n10862 = ~n10803 & n10861;
  assign n10863 = n10862 ^ n10800;
  assign n10864 = n10863 ^ n10691;
  assign n10865 = ~n10797 & n10864;
  assign n10866 = n10865 ^ n10796;
  assign n10867 = n10866 ^ n10686;
  assign n10868 = n10793 & ~n10867;
  assign n10869 = n10868 ^ n10792;
  assign n10870 = n10869 ^ n10679;
  assign n10871 = ~n10789 & ~n10870;
  assign n10872 = n10871 ^ n10788;
  assign n10873 = n10872 ^ n10672;
  assign n10874 = ~n10785 & n10873;
  assign n10875 = n10874 ^ n10784;
  assign n10876 = n10875 ^ n10140;
  assign n10877 = ~n10781 & ~n10876;
  assign n10878 = n10877 ^ n10780;
  assign n10879 = n10878 ^ n10776;
  assign n10880 = ~n10777 & ~n10879;
  assign n10881 = n10880 ^ n10775;
  assign n10882 = n10881 ^ n10768;
  assign n10883 = ~n10772 & ~n10882;
  assign n10884 = n10883 ^ n10771;
  assign n10885 = n10884 ^ n10763;
  assign n10886 = n10767 & n10885;
  assign n10887 = n10886 ^ n10766;
  assign n10888 = n10887 ^ n10757;
  assign n10889 = ~n10761 & n10888;
  assign n10890 = n10889 ^ n10760;
  assign n10891 = n10890 ^ n10752;
  assign n10892 = ~n10756 & n10891;
  assign n10893 = n10892 ^ n10755;
  assign n10894 = n10893 ^ n10746;
  assign n10895 = ~n10750 & ~n10894;
  assign n10896 = n10895 ^ n10749;
  assign n10897 = n10896 ^ n10741;
  assign n10898 = n10745 & ~n10897;
  assign n10899 = n10898 ^ n10744;
  assign n10900 = n10899 ^ n10735;
  assign n10901 = n10739 & n10900;
  assign n10902 = n10901 ^ n10738;
  assign n10733 = n10492 ^ x430;
  assign n10734 = n10733 ^ n10448;
  assign n10903 = n10902 ^ n10734;
  assign n10904 = n9776 ^ n9110;
  assign n10905 = ~n10537 & n10904;
  assign n10906 = n10905 ^ n9110;
  assign n10907 = n10906 ^ n10734;
  assign n10908 = n10903 & n10907;
  assign n10909 = n10908 ^ n10906;
  assign n10729 = n9796 ^ n9103;
  assign n10730 = n10569 & n10729;
  assign n10731 = n10730 ^ n9103;
  assign n10945 = n10909 ^ n10731;
  assign n10728 = n10495 ^ n10447;
  assign n10946 = n10945 ^ n10728;
  assign n10947 = n10946 ^ n8661;
  assign n10948 = n10906 ^ n10903;
  assign n10949 = n10948 ^ n8616;
  assign n10950 = n10899 ^ n10739;
  assign n10951 = n10950 ^ n8580;
  assign n10952 = n10896 ^ n10745;
  assign n10953 = n10952 ^ n8233;
  assign n10954 = n10893 ^ n10750;
  assign n10955 = n10954 ^ n8221;
  assign n10956 = n10890 ^ n10756;
  assign n10957 = n10956 ^ n7769;
  assign n10958 = n10887 ^ n10761;
  assign n10959 = n10958 ^ n7777;
  assign n10960 = n10884 ^ n10767;
  assign n10961 = n10960 ^ n7783;
  assign n10962 = n10881 ^ n10772;
  assign n10963 = n10962 ^ n7791;
  assign n10964 = n10878 ^ n10777;
  assign n10965 = n10964 ^ n7797;
  assign n10966 = n10875 ^ n10781;
  assign n10967 = n10966 ^ n7805;
  assign n10968 = n10872 ^ n10785;
  assign n10969 = n10968 ^ n7811;
  assign n10970 = n10869 ^ n10789;
  assign n10971 = n10970 ^ n7819;
  assign n10972 = n10866 ^ n10793;
  assign n10973 = n10972 ^ n7825;
  assign n10974 = n10863 ^ n10797;
  assign n10975 = n10974 ^ n7832;
  assign n10976 = n10860 ^ n10803;
  assign n10977 = n10976 ^ n7838;
  assign n10978 = n10857 ^ n10808;
  assign n10979 = n10978 ^ n7847;
  assign n10980 = n10854 ^ n10813;
  assign n10981 = n10980 ^ n7853;
  assign n10982 = n10851 ^ n10816;
  assign n10983 = n10982 ^ n10817;
  assign n10984 = n10983 ^ n7859;
  assign n10985 = n10848 ^ n10843;
  assign n10986 = n10985 ^ n10840;
  assign n10987 = n10986 ^ n7864;
  assign n10641 = n10640 ^ n10637;
  assign n10666 = n10665 ^ n10641;
  assign n10667 = n10666 ^ n7870;
  assign n10616 = n10615 ^ n10607;
  assign n10631 = n10616 ^ n7875;
  assign n10543 = n10542 ^ n10147;
  assign n10576 = ~n7883 & ~n10543;
  assign n10577 = n10576 ^ n7881;
  assign n10549 = n10548 ^ n10545;
  assign n10575 = n10574 ^ n10549;
  assign n10580 = n10576 ^ n10575;
  assign n10581 = ~n10577 & n10580;
  assign n10582 = n10581 ^ n7881;
  assign n10632 = n10616 ^ n10582;
  assign n10633 = ~n10631 & n10632;
  assign n10634 = n10633 ^ n7875;
  assign n10988 = n10666 ^ n10634;
  assign n10989 = ~n10667 & ~n10988;
  assign n10990 = n10989 ^ n7870;
  assign n10991 = n10990 ^ n10986;
  assign n10992 = ~n10987 & ~n10991;
  assign n10993 = n10992 ^ n7864;
  assign n10994 = n10993 ^ n10983;
  assign n10995 = n10984 & ~n10994;
  assign n10996 = n10995 ^ n7859;
  assign n10997 = n10996 ^ n10980;
  assign n10998 = ~n10981 & ~n10997;
  assign n10999 = n10998 ^ n7853;
  assign n11000 = n10999 ^ n10978;
  assign n11001 = ~n10979 & ~n11000;
  assign n11002 = n11001 ^ n7847;
  assign n11003 = n11002 ^ n10976;
  assign n11004 = n10977 & ~n11003;
  assign n11005 = n11004 ^ n7838;
  assign n11006 = n11005 ^ n10974;
  assign n11007 = ~n10975 & ~n11006;
  assign n11008 = n11007 ^ n7832;
  assign n11009 = n11008 ^ n10972;
  assign n11010 = ~n10973 & ~n11009;
  assign n11011 = n11010 ^ n7825;
  assign n11012 = n11011 ^ n10970;
  assign n11013 = n10971 & ~n11012;
  assign n11014 = n11013 ^ n7819;
  assign n11015 = n11014 ^ n10968;
  assign n11016 = ~n10969 & n11015;
  assign n11017 = n11016 ^ n7811;
  assign n11018 = n11017 ^ n10966;
  assign n11019 = n10967 & n11018;
  assign n11020 = n11019 ^ n7805;
  assign n11021 = n11020 ^ n10964;
  assign n11022 = n10965 & n11021;
  assign n11023 = n11022 ^ n7797;
  assign n11024 = n11023 ^ n10962;
  assign n11025 = ~n10963 & n11024;
  assign n11026 = n11025 ^ n7791;
  assign n11027 = n11026 ^ n10960;
  assign n11028 = ~n10961 & n11027;
  assign n11029 = n11028 ^ n7783;
  assign n11030 = n11029 ^ n10958;
  assign n11031 = ~n10959 & n11030;
  assign n11032 = n11031 ^ n7777;
  assign n11033 = n11032 ^ n10956;
  assign n11034 = ~n10957 & n11033;
  assign n11035 = n11034 ^ n7769;
  assign n11036 = n11035 ^ n10954;
  assign n11037 = ~n10955 & n11036;
  assign n11038 = n11037 ^ n8221;
  assign n11039 = n11038 ^ n10952;
  assign n11040 = n10953 & n11039;
  assign n11041 = n11040 ^ n8233;
  assign n11042 = n11041 ^ n10950;
  assign n11043 = ~n10951 & ~n11042;
  assign n11044 = n11043 ^ n8580;
  assign n11045 = n11044 ^ n10948;
  assign n11046 = ~n10949 & ~n11045;
  assign n11047 = n11046 ^ n8616;
  assign n11048 = n11047 ^ n10946;
  assign n11049 = ~n10947 & n11048;
  assign n11050 = n11049 ^ n8661;
  assign n10732 = n10731 ^ n10728;
  assign n10910 = n10909 ^ n10728;
  assign n10911 = ~n10732 & n10910;
  assign n10912 = n10911 ^ n10731;
  assign n10724 = n9963 ^ n9095;
  assign n10725 = ~n10602 & n10724;
  assign n10726 = n10725 ^ n9095;
  assign n10722 = n10498 ^ x428;
  assign n10723 = n10722 ^ n10444;
  assign n10727 = n10726 ^ n10723;
  assign n10943 = n10912 ^ n10727;
  assign n10944 = n10943 ^ n8719;
  assign n11084 = n11050 ^ n10944;
  assign n11085 = n11044 ^ n10949;
  assign n11086 = n11038 ^ n10953;
  assign n11087 = n11032 ^ n10957;
  assign n11088 = n11014 ^ n10969;
  assign n11089 = n11011 ^ n10971;
  assign n10544 = n10543 ^ n7883;
  assign n10578 = n10577 ^ n10575;
  assign n10579 = n10544 & n10578;
  assign n10583 = n10582 ^ n7875;
  assign n10617 = n10616 ^ n10583;
  assign n10630 = n10579 & n10617;
  assign n10668 = n10667 ^ n10634;
  assign n11090 = ~n10630 & ~n10668;
  assign n11091 = n10990 ^ n10987;
  assign n11092 = n11090 & n11091;
  assign n11093 = n10993 ^ n10984;
  assign n11094 = ~n11092 & ~n11093;
  assign n11095 = n10996 ^ n10981;
  assign n11096 = n11094 & n11095;
  assign n11097 = n10999 ^ n10979;
  assign n11098 = ~n11096 & n11097;
  assign n11099 = n11002 ^ n10977;
  assign n11100 = n11098 & n11099;
  assign n11101 = n11005 ^ n10975;
  assign n11102 = ~n11100 & n11101;
  assign n11103 = n11008 ^ n10973;
  assign n11104 = n11102 & ~n11103;
  assign n11105 = n11089 & ~n11104;
  assign n11106 = ~n11088 & n11105;
  assign n11107 = n11017 ^ n10967;
  assign n11108 = n11106 & n11107;
  assign n11109 = n11020 ^ n10965;
  assign n11110 = n11108 & ~n11109;
  assign n11111 = n11023 ^ n10963;
  assign n11112 = ~n11110 & n11111;
  assign n11113 = n11026 ^ n10961;
  assign n11114 = n11112 & n11113;
  assign n11115 = n11029 ^ n10959;
  assign n11116 = ~n11114 & ~n11115;
  assign n11117 = n11087 & ~n11116;
  assign n11118 = n11035 ^ n10955;
  assign n11119 = n11117 & n11118;
  assign n11120 = ~n11086 & n11119;
  assign n11121 = n11041 ^ n10951;
  assign n11122 = n11120 & ~n11121;
  assign n11123 = n11085 & n11122;
  assign n11124 = n11047 ^ n8661;
  assign n11125 = n11124 ^ n10946;
  assign n11126 = ~n11123 & n11125;
  assign n11127 = n11084 & ~n11126;
  assign n11051 = n11050 ^ n10943;
  assign n11052 = n10944 & n11051;
  assign n11053 = n11052 ^ n8719;
  assign n10913 = n10912 ^ n10723;
  assign n10914 = ~n10727 & ~n10913;
  assign n10915 = n10914 ^ n10726;
  assign n10718 = n9436 ^ n8589;
  assign n10719 = n10656 & n10718;
  assign n10720 = n10719 ^ n8589;
  assign n10940 = n10915 ^ n10720;
  assign n10717 = n10501 ^ n10443;
  assign n10941 = n10940 ^ n10717;
  assign n10942 = n10941 ^ n8140;
  assign n11128 = n11053 ^ n10942;
  assign n11129 = ~n11127 & n11128;
  assign n11054 = n11053 ^ n10941;
  assign n11055 = n10942 & n11054;
  assign n11056 = n11055 ^ n8140;
  assign n10721 = n10720 ^ n10717;
  assign n10916 = n10915 ^ n10717;
  assign n10917 = ~n10721 & n10916;
  assign n10918 = n10917 ^ n10720;
  assign n10713 = n9430 ^ n8586;
  assign n10714 = n10712 & ~n10713;
  assign n10715 = n10714 ^ n8586;
  assign n10937 = n10918 ^ n10715;
  assign n10710 = n10504 ^ x426;
  assign n10711 = n10710 ^ n10440;
  assign n10938 = n10937 ^ n10711;
  assign n10939 = n10938 ^ n8134;
  assign n11083 = n11056 ^ n10939;
  assign n11143 = n11129 ^ n11083;
  assign n11144 = n11143 ^ x453;
  assign n11145 = n11128 ^ n11127;
  assign n11146 = n11145 ^ x454;
  assign n11147 = n11126 ^ n11084;
  assign n11148 = n11147 ^ x455;
  assign n11149 = n11125 ^ n11123;
  assign n11150 = n11149 ^ x456;
  assign n11151 = n11122 ^ n11085;
  assign n11152 = n11151 ^ x457;
  assign n11153 = n11121 ^ n11120;
  assign n11154 = n11153 ^ x458;
  assign n11155 = n11119 ^ n11086;
  assign n11156 = n11155 ^ x459;
  assign n11157 = n11118 ^ n11117;
  assign n11158 = n11157 ^ x460;
  assign n11159 = n11116 ^ n11087;
  assign n11160 = n11159 ^ x461;
  assign n11161 = n11115 ^ n11114;
  assign n11162 = n11161 ^ x462;
  assign n11227 = n11113 ^ n11112;
  assign n11163 = n11111 ^ n11110;
  assign n11164 = n11163 ^ x464;
  assign n11165 = n11109 ^ n11108;
  assign n11166 = n11165 ^ x465;
  assign n11167 = n11107 ^ n11106;
  assign n11168 = n11167 ^ x466;
  assign n11169 = n11105 ^ n11088;
  assign n11170 = n11169 ^ x467;
  assign n11171 = n11104 ^ n11089;
  assign n11172 = n11171 ^ x468;
  assign n11173 = n11103 ^ n11102;
  assign n11174 = n11173 ^ x469;
  assign n11175 = n11101 ^ n11100;
  assign n11176 = n11175 ^ x470;
  assign n11177 = n11099 ^ n11098;
  assign n11178 = n11177 ^ x471;
  assign n11179 = n11097 ^ n11096;
  assign n11180 = n11179 ^ x472;
  assign n11181 = n11095 ^ n11094;
  assign n11182 = n11181 ^ x473;
  assign n11183 = n11093 ^ n11092;
  assign n11184 = n11183 ^ x474;
  assign n11185 = n11091 ^ n11090;
  assign n11186 = n11185 ^ x475;
  assign n10669 = n10668 ^ n10630;
  assign n11187 = n10669 ^ x476;
  assign n10618 = n10617 ^ n10579;
  assign n10619 = n10618 ^ x477;
  assign n10620 = x479 & ~n10544;
  assign n10621 = n10620 ^ x478;
  assign n10622 = n10578 ^ n10544;
  assign n10623 = n10622 ^ n10620;
  assign n10624 = n10621 & ~n10623;
  assign n10625 = n10624 ^ x478;
  assign n10626 = n10625 ^ n10618;
  assign n10627 = n10619 & ~n10626;
  assign n10628 = n10627 ^ x477;
  assign n11188 = n10669 ^ n10628;
  assign n11189 = ~n11187 & n11188;
  assign n11190 = n11189 ^ x476;
  assign n11191 = n11190 ^ n11185;
  assign n11192 = ~n11186 & n11191;
  assign n11193 = n11192 ^ x475;
  assign n11194 = n11193 ^ n11183;
  assign n11195 = n11184 & ~n11194;
  assign n11196 = n11195 ^ x474;
  assign n11197 = n11196 ^ n11181;
  assign n11198 = n11182 & ~n11197;
  assign n11199 = n11198 ^ x473;
  assign n11200 = n11199 ^ n11179;
  assign n11201 = n11180 & ~n11200;
  assign n11202 = n11201 ^ x472;
  assign n11203 = n11202 ^ n11177;
  assign n11204 = ~n11178 & n11203;
  assign n11205 = n11204 ^ x471;
  assign n11206 = n11205 ^ n11175;
  assign n11207 = ~n11176 & n11206;
  assign n11208 = n11207 ^ x470;
  assign n11209 = n11208 ^ n11173;
  assign n11210 = ~n11174 & n11209;
  assign n11211 = n11210 ^ x469;
  assign n11212 = n11211 ^ n11171;
  assign n11213 = n11172 & ~n11212;
  assign n11214 = n11213 ^ x468;
  assign n11215 = n11214 ^ n11169;
  assign n11216 = n11170 & ~n11215;
  assign n11217 = n11216 ^ x467;
  assign n11218 = n11217 ^ n11167;
  assign n11219 = ~n11168 & n11218;
  assign n11220 = n11219 ^ x466;
  assign n11221 = n11220 ^ n11165;
  assign n11222 = n11166 & ~n11221;
  assign n11223 = n11222 ^ x465;
  assign n11224 = n11223 ^ n11163;
  assign n11225 = ~n11164 & n11224;
  assign n11226 = n11225 ^ x464;
  assign n11228 = n11227 ^ n11226;
  assign n11229 = n11227 ^ x463;
  assign n11230 = ~n11228 & n11229;
  assign n11231 = n11230 ^ x463;
  assign n11232 = n11231 ^ n11161;
  assign n11233 = ~n11162 & n11232;
  assign n11234 = n11233 ^ x462;
  assign n11235 = n11234 ^ n11159;
  assign n11236 = ~n11160 & n11235;
  assign n11237 = n11236 ^ x461;
  assign n11238 = n11237 ^ n11157;
  assign n11239 = n11158 & ~n11238;
  assign n11240 = n11239 ^ x460;
  assign n11241 = n11240 ^ n11155;
  assign n11242 = ~n11156 & n11241;
  assign n11243 = n11242 ^ x459;
  assign n11244 = n11243 ^ n11153;
  assign n11245 = ~n11154 & n11244;
  assign n11246 = n11245 ^ x458;
  assign n11247 = n11246 ^ n11151;
  assign n11248 = n11152 & ~n11247;
  assign n11249 = n11248 ^ x457;
  assign n11250 = n11249 ^ n11149;
  assign n11251 = n11150 & ~n11250;
  assign n11252 = n11251 ^ x456;
  assign n11253 = n11252 ^ n11147;
  assign n11254 = ~n11148 & n11253;
  assign n11255 = n11254 ^ x455;
  assign n11256 = n11255 ^ n11145;
  assign n11257 = n11146 & ~n11256;
  assign n11258 = n11257 ^ x454;
  assign n11259 = n11258 ^ n11143;
  assign n11260 = n11144 & ~n11259;
  assign n11261 = n11260 ^ x453;
  assign n11306 = n11261 ^ x452;
  assign n11130 = ~n11083 & ~n11129;
  assign n11057 = n11056 ^ n10938;
  assign n11058 = ~n10939 & ~n11057;
  assign n11059 = n11058 ^ n8134;
  assign n10716 = n10715 ^ n10711;
  assign n10919 = n10918 ^ n10711;
  assign n10920 = ~n10716 & ~n10919;
  assign n10921 = n10920 ^ n10715;
  assign n10706 = n9446 ^ n8622;
  assign n10707 = ~n9987 & ~n10706;
  assign n10708 = n10707 ^ n8622;
  assign n10934 = n10921 ^ n10708;
  assign n10705 = n10507 ^ n10439;
  assign n10935 = n10934 ^ n10705;
  assign n10936 = n10935 ^ n8132;
  assign n11082 = n11059 ^ n10936;
  assign n11141 = n11130 ^ n11082;
  assign n11307 = n11306 ^ n11141;
  assign n11364 = n11310 ^ n11307;
  assign n11414 = n11364 ^ n8784;
  assign n11990 = n11414 ^ x511;
  assign n10676 = n10625 ^ n10619;
  assign n12606 = n10804 ^ n10676;
  assign n12607 = n11990 & ~n12606;
  assign n12608 = n12607 ^ n10804;
  assign n11764 = n11249 ^ x456;
  assign n11765 = n11764 ^ n11149;
  assign n11076 = n10516 ^ x422;
  assign n11077 = n11076 ^ n10432;
  assign n12099 = n11077 ^ n10656;
  assign n12100 = n11765 & n12099;
  assign n12101 = n12100 ^ n10656;
  assign n11488 = n11196 ^ n11182;
  assign n11485 = n10182 ^ n9143;
  assign n11486 = ~n10763 & ~n11485;
  assign n11487 = n11486 ^ n9143;
  assign n11489 = n11488 ^ n11487;
  assign n11402 = n11193 ^ x474;
  assign n11403 = n11402 ^ n11183;
  assign n11399 = n10187 ^ n9150;
  assign n11400 = ~n10768 & n11399;
  assign n11401 = n11400 ^ n9150;
  assign n11404 = n11403 ^ n11401;
  assign n11345 = n11190 ^ n11186;
  assign n11342 = n10190 ^ n9156;
  assign n11343 = n10776 & ~n11342;
  assign n11344 = n11343 ^ n9156;
  assign n11346 = n11345 ^ n11344;
  assign n10629 = n10628 ^ x476;
  assign n10670 = n10669 ^ n10629;
  assign n10142 = n10141 ^ n9161;
  assign n10143 = ~n10140 & n10142;
  assign n10144 = n10143 ^ n9161;
  assign n10671 = n10670 ^ n10144;
  assign n10673 = n10199 ^ n9166;
  assign n10674 = n10672 & n10673;
  assign n10675 = n10674 ^ n9166;
  assign n10677 = n10676 ^ n10675;
  assign n10680 = n10204 ^ n9172;
  assign n10681 = n10679 & ~n10680;
  assign n10682 = n10681 ^ n9172;
  assign n10678 = n10622 ^ n10621;
  assign n10683 = n10682 ^ n10678;
  assign n10687 = n10210 ^ n9178;
  assign n10688 = n10686 & n10687;
  assign n10689 = n10688 ^ n9178;
  assign n10684 = n10544 ^ x479;
  assign n10690 = n10689 ^ n10684;
  assign n11286 = n10519 ^ n10431;
  assign n11283 = n9206 ^ n8786;
  assign n11284 = ~n9969 & ~n11283;
  assign n11285 = n11284 ^ n8786;
  assign n11287 = n11286 ^ n11285;
  assign n11288 = n11287 ^ n7292;
  assign n10701 = n9424 ^ n8667;
  assign n10702 = ~n9981 & ~n10701;
  assign n10703 = n10702 ^ n8667;
  assign n10699 = n10510 ^ x424;
  assign n10700 = n10699 ^ n10436;
  assign n10704 = n10703 ^ n10700;
  assign n10709 = n10708 ^ n10705;
  assign n10922 = n10921 ^ n10705;
  assign n10923 = n10709 & n10922;
  assign n10924 = n10923 ^ n10708;
  assign n10925 = n10924 ^ n10700;
  assign n10926 = n10704 & n10925;
  assign n10927 = n10926 ^ n10703;
  assign n10698 = n10513 ^ n10435;
  assign n10928 = n10927 ^ n10698;
  assign n10695 = n9418 ^ n8725;
  assign n10696 = ~n9997 & ~n10695;
  assign n10697 = n10696 ^ n8725;
  assign n11073 = n10698 ^ n10697;
  assign n11074 = ~n10928 & ~n11073;
  assign n11075 = n11074 ^ n10697;
  assign n11078 = n11077 ^ n11075;
  assign n11070 = n9210 ^ n8791;
  assign n11071 = n9975 & ~n11070;
  assign n11072 = n11071 ^ n8791;
  assign n11280 = n11077 ^ n11072;
  assign n11281 = n11078 & ~n11280;
  assign n11282 = n11281 ^ n11072;
  assign n11289 = n11288 ^ n11282;
  assign n11079 = n11078 ^ n11072;
  assign n10929 = n10928 ^ n10697;
  assign n10930 = n10929 ^ n8121;
  assign n10931 = n10924 ^ n10703;
  assign n10932 = n10931 ^ n10700;
  assign n10933 = n10932 ^ n8127;
  assign n11060 = n11059 ^ n10935;
  assign n11061 = ~n10936 & n11060;
  assign n11062 = n11061 ^ n8132;
  assign n11063 = n11062 ^ n10932;
  assign n11064 = ~n10933 & ~n11063;
  assign n11065 = n11064 ^ n8127;
  assign n11066 = n11065 ^ n10929;
  assign n11067 = n10930 & n11066;
  assign n11068 = n11067 ^ n8121;
  assign n11069 = n11068 ^ n7892;
  assign n11080 = n11079 ^ n11069;
  assign n11081 = n11065 ^ n10930;
  assign n11131 = ~n11082 & ~n11130;
  assign n11132 = n11062 ^ n10933;
  assign n11133 = n11131 & ~n11132;
  assign n11134 = n11081 & ~n11133;
  assign n11279 = n11080 & ~n11134;
  assign n11290 = n11289 ^ n11279;
  assign n11275 = n11079 ^ n7892;
  assign n11276 = n11079 ^ n11068;
  assign n11277 = n11275 & n11276;
  assign n11278 = n11277 ^ n7892;
  assign n11291 = n11290 ^ n11278;
  assign n11135 = n11134 ^ n11080;
  assign n11136 = n11135 ^ x449;
  assign n11137 = n11133 ^ n11081;
  assign n11138 = n11137 ^ x450;
  assign n11139 = n11132 ^ n11131;
  assign n11140 = n11139 ^ x451;
  assign n11142 = n11141 ^ x452;
  assign n11262 = n11261 ^ n11141;
  assign n11263 = ~n11142 & n11262;
  assign n11264 = n11263 ^ x452;
  assign n11265 = n11264 ^ n11139;
  assign n11266 = n11140 & ~n11265;
  assign n11267 = n11266 ^ x451;
  assign n11268 = n11267 ^ n11137;
  assign n11269 = ~n11138 & n11268;
  assign n11270 = n11269 ^ x450;
  assign n11271 = n11270 ^ n11135;
  assign n11272 = n11136 & ~n11271;
  assign n11273 = n11272 ^ x449;
  assign n11274 = n11273 ^ x448;
  assign n11292 = n11291 ^ n11274;
  assign n10692 = n10216 ^ n9180;
  assign n10693 = ~n10691 & ~n10692;
  assign n10694 = n10693 ^ n9180;
  assign n11293 = n11292 ^ n10694;
  assign n11318 = n10222 ^ n9189;
  assign n11319 = ~n10802 & n11318;
  assign n11320 = n11319 ^ n9189;
  assign n11296 = n10227 ^ n8733;
  assign n11297 = ~n10804 & n11296;
  assign n11298 = n11297 ^ n8733;
  assign n11294 = n11267 ^ x450;
  assign n11295 = n11294 ^ n11137;
  assign n11299 = n11298 ^ n11295;
  assign n11302 = n10132 ^ n9199;
  assign n11303 = ~n10809 & n11302;
  assign n11304 = n11303 ^ n9199;
  assign n11300 = n11264 ^ x451;
  assign n11301 = n11300 ^ n11139;
  assign n11305 = n11304 ^ n11301;
  assign n11311 = ~n11307 & ~n11310;
  assign n11312 = n11311 ^ n11301;
  assign n11313 = n11305 & n11312;
  assign n11314 = n11313 ^ n11311;
  assign n11315 = n11314 ^ n11295;
  assign n11316 = ~n11299 & n11315;
  assign n11317 = n11316 ^ n11298;
  assign n11321 = n11320 ^ n11317;
  assign n11322 = n11270 ^ x449;
  assign n11323 = n11322 ^ n11135;
  assign n11324 = n11323 ^ n11317;
  assign n11325 = ~n11321 & ~n11324;
  assign n11326 = n11325 ^ n11320;
  assign n11327 = n11326 ^ n11292;
  assign n11328 = ~n11293 & ~n11327;
  assign n11329 = n11328 ^ n10694;
  assign n11330 = n11329 ^ n10684;
  assign n11331 = n10690 & n11330;
  assign n11332 = n11331 ^ n10689;
  assign n11333 = n11332 ^ n10678;
  assign n11334 = ~n10683 & n11333;
  assign n11335 = n11334 ^ n10682;
  assign n11336 = n11335 ^ n10676;
  assign n11337 = ~n10677 & n11336;
  assign n11338 = n11337 ^ n10675;
  assign n11339 = n11338 ^ n10670;
  assign n11340 = ~n10671 & ~n11339;
  assign n11341 = n11340 ^ n10144;
  assign n11396 = n11345 ^ n11341;
  assign n11397 = n11346 & n11396;
  assign n11398 = n11397 ^ n11344;
  assign n11482 = n11403 ^ n11398;
  assign n11483 = ~n11404 & n11482;
  assign n11484 = n11483 ^ n11401;
  assign n11490 = n11489 ^ n11484;
  assign n11491 = n11490 ^ n8957;
  assign n11405 = n11404 ^ n11398;
  assign n11406 = n11405 ^ n8941;
  assign n11347 = n11346 ^ n11341;
  assign n11348 = n11347 ^ n8901;
  assign n11349 = n11338 ^ n10671;
  assign n11350 = n11349 ^ n8738;
  assign n11351 = n11335 ^ n10677;
  assign n11352 = n11351 ^ n8742;
  assign n11353 = n11332 ^ n10683;
  assign n11354 = n11353 ^ n8748;
  assign n11355 = n11329 ^ n10690;
  assign n11356 = n11355 ^ n8754;
  assign n11357 = n11326 ^ n11293;
  assign n11358 = n11357 ^ n8734;
  assign n11359 = n11323 ^ n11321;
  assign n11360 = n11359 ^ n8764;
  assign n11361 = n11314 ^ n11298;
  assign n11362 = n11361 ^ n11295;
  assign n11363 = n11362 ^ n8769;
  assign n11365 = ~n8784 & n11364;
  assign n11366 = n11365 ^ n8775;
  assign n11367 = n11311 ^ n11304;
  assign n11368 = n11367 ^ n11301;
  assign n11369 = n11368 ^ n11365;
  assign n11370 = ~n11366 & n11369;
  assign n11371 = n11370 ^ n8775;
  assign n11372 = n11371 ^ n11362;
  assign n11373 = ~n11363 & ~n11372;
  assign n11374 = n11373 ^ n8769;
  assign n11375 = n11374 ^ n11359;
  assign n11376 = n11360 & n11375;
  assign n11377 = n11376 ^ n8764;
  assign n11378 = n11377 ^ n11357;
  assign n11379 = n11358 & n11378;
  assign n11380 = n11379 ^ n8734;
  assign n11381 = n11380 ^ n11355;
  assign n11382 = ~n11356 & ~n11381;
  assign n11383 = n11382 ^ n8754;
  assign n11384 = n11383 ^ n11353;
  assign n11385 = ~n11354 & n11384;
  assign n11386 = n11385 ^ n8748;
  assign n11387 = n11386 ^ n11351;
  assign n11388 = n11352 & n11387;
  assign n11389 = n11388 ^ n8742;
  assign n11390 = n11389 ^ n11349;
  assign n11391 = n11350 & ~n11390;
  assign n11392 = n11391 ^ n8738;
  assign n11393 = n11392 ^ n11347;
  assign n11394 = n11348 & ~n11393;
  assign n11395 = n11394 ^ n8901;
  assign n11479 = n11405 ^ n11395;
  assign n11480 = n11406 & ~n11479;
  assign n11481 = n11480 ^ n8941;
  assign n11492 = n11491 ^ n11481;
  assign n11407 = n11406 ^ n11395;
  assign n11408 = n11386 ^ n11352;
  assign n11409 = n11383 ^ n11354;
  assign n11410 = n11380 ^ n11356;
  assign n11411 = n11377 ^ n11358;
  assign n11412 = n11374 ^ n11360;
  assign n11413 = n11371 ^ n11363;
  assign n11415 = n11368 ^ n11366;
  assign n11416 = ~n11414 & n11415;
  assign n11417 = n11413 & n11416;
  assign n11418 = ~n11412 & ~n11417;
  assign n11419 = n11411 & n11418;
  assign n11420 = ~n11410 & ~n11419;
  assign n11421 = n11409 & n11420;
  assign n11422 = n11408 & ~n11421;
  assign n11423 = n11389 ^ n11350;
  assign n11424 = n11422 & ~n11423;
  assign n11425 = n11392 ^ n11348;
  assign n11426 = ~n11424 & n11425;
  assign n11493 = n11407 & n11426;
  assign n11714 = n11492 & ~n11493;
  assign n11653 = n11490 ^ n11481;
  assign n11654 = ~n11491 & ~n11653;
  assign n11655 = n11654 ^ n8957;
  assign n11574 = n11488 ^ n11484;
  assign n11575 = ~n11489 & n11574;
  assign n11576 = n11575 ^ n11487;
  assign n11571 = n11199 ^ x472;
  assign n11572 = n11571 ^ n11179;
  assign n11568 = n10176 ^ n9131;
  assign n11569 = n10757 & n11568;
  assign n11570 = n11569 ^ n9131;
  assign n11573 = n11572 ^ n11570;
  assign n11651 = n11576 ^ n11573;
  assign n11652 = n11651 ^ n8972;
  assign n11715 = n11655 ^ n11652;
  assign n11716 = n11714 & ~n11715;
  assign n11656 = n11655 ^ n11651;
  assign n11657 = ~n11652 & n11656;
  assign n11658 = n11657 ^ n8972;
  assign n11577 = n11576 ^ n11572;
  assign n11578 = ~n11573 & n11577;
  assign n11579 = n11578 ^ n11570;
  assign n11565 = n11202 ^ x471;
  assign n11566 = n11565 ^ n11177;
  assign n11562 = n10171 ^ n9125;
  assign n11563 = n10752 & n11562;
  assign n11564 = n11563 ^ n9125;
  assign n11567 = n11566 ^ n11564;
  assign n11649 = n11579 ^ n11567;
  assign n11650 = n11649 ^ n8989;
  assign n11717 = n11658 ^ n11650;
  assign n11718 = n11716 & ~n11717;
  assign n11659 = n11658 ^ n11649;
  assign n11660 = ~n11650 & ~n11659;
  assign n11661 = n11660 ^ n8989;
  assign n11580 = n11579 ^ n11566;
  assign n11581 = n11567 & ~n11580;
  assign n11582 = n11581 ^ n11564;
  assign n11558 = n10165 ^ n9123;
  assign n11559 = ~n10746 & n11558;
  assign n11560 = n11559 ^ n9123;
  assign n11557 = n11205 ^ n11176;
  assign n11561 = n11560 ^ n11557;
  assign n11647 = n11582 ^ n11561;
  assign n11648 = n11647 ^ n9087;
  assign n11719 = n11661 ^ n11648;
  assign n11720 = n11718 & ~n11719;
  assign n11662 = n11661 ^ n11647;
  assign n11663 = n11648 & n11662;
  assign n11664 = n11663 ^ n9087;
  assign n11583 = n11582 ^ n11557;
  assign n11584 = n11561 & ~n11583;
  assign n11585 = n11584 ^ n11560;
  assign n11555 = n11208 ^ n11174;
  assign n11552 = n10275 ^ n9122;
  assign n11553 = n10741 & ~n11552;
  assign n11554 = n11553 ^ n9122;
  assign n11556 = n11555 ^ n11554;
  assign n11645 = n11585 ^ n11556;
  assign n11646 = n11645 ^ n9146;
  assign n11721 = n11664 ^ n11646;
  assign n11722 = ~n11720 & n11721;
  assign n11665 = n11664 ^ n11645;
  assign n11666 = ~n11646 & ~n11665;
  assign n11667 = n11666 ^ n9146;
  assign n11586 = n11585 ^ n11555;
  assign n11587 = n11556 & ~n11586;
  assign n11588 = n11587 ^ n11554;
  assign n11549 = n11211 ^ x468;
  assign n11550 = n11549 ^ n11171;
  assign n11546 = n10160 ^ n9115;
  assign n11547 = ~n10735 & n11546;
  assign n11548 = n11547 ^ n9115;
  assign n11551 = n11550 ^ n11548;
  assign n11643 = n11588 ^ n11551;
  assign n11644 = n11643 ^ n9138;
  assign n11723 = n11667 ^ n11644;
  assign n11724 = n11722 & n11723;
  assign n11668 = n11667 ^ n11643;
  assign n11669 = n11644 & n11668;
  assign n11670 = n11669 ^ n9138;
  assign n11589 = n11588 ^ n11550;
  assign n11590 = n11551 & n11589;
  assign n11591 = n11590 ^ n11548;
  assign n11542 = n10155 ^ n9109;
  assign n11543 = n10734 & ~n11542;
  assign n11544 = n11543 ^ n9109;
  assign n11640 = n11591 ^ n11544;
  assign n11541 = n11214 ^ n11170;
  assign n11641 = n11640 ^ n11541;
  assign n11642 = n11641 ^ n9133;
  assign n11713 = n11670 ^ n11642;
  assign n11792 = n11724 ^ n11713;
  assign n11793 = n11792 ^ x494;
  assign n11818 = n11723 ^ n11722;
  assign n11794 = n11721 ^ n11720;
  assign n11795 = n11794 ^ x496;
  assign n11796 = n11719 ^ n11718;
  assign n11797 = n11796 ^ x497;
  assign n11798 = n11717 ^ n11716;
  assign n11799 = n11798 ^ x498;
  assign n11800 = n11715 ^ n11714;
  assign n11801 = n11800 ^ x499;
  assign n11494 = n11493 ^ n11492;
  assign n11802 = n11494 ^ x500;
  assign n11427 = n11426 ^ n11407;
  assign n11428 = n11427 ^ x501;
  assign n11429 = n11425 ^ n11424;
  assign n11430 = n11429 ^ x502;
  assign n11431 = n11423 ^ n11422;
  assign n11432 = n11431 ^ x503;
  assign n11433 = n11421 ^ n11408;
  assign n11434 = n11433 ^ x504;
  assign n11435 = n11420 ^ n11409;
  assign n11436 = n11435 ^ x505;
  assign n11437 = n11419 ^ n11410;
  assign n11438 = n11437 ^ x506;
  assign n11439 = n11418 ^ n11411;
  assign n11440 = n11439 ^ x507;
  assign n11441 = n11417 ^ n11412;
  assign n11442 = n11441 ^ x508;
  assign n11443 = n11416 ^ n11413;
  assign n11444 = n11443 ^ x509;
  assign n11445 = x511 & n11414;
  assign n11446 = n11445 ^ x510;
  assign n11447 = n11415 ^ n11414;
  assign n11448 = n11447 ^ n11445;
  assign n11449 = n11446 & n11448;
  assign n11450 = n11449 ^ x510;
  assign n11451 = n11450 ^ n11443;
  assign n11452 = n11444 & ~n11451;
  assign n11453 = n11452 ^ x509;
  assign n11454 = n11453 ^ n11441;
  assign n11455 = ~n11442 & n11454;
  assign n11456 = n11455 ^ x508;
  assign n11457 = n11456 ^ n11439;
  assign n11458 = ~n11440 & n11457;
  assign n11459 = n11458 ^ x507;
  assign n11460 = n11459 ^ n11437;
  assign n11461 = n11438 & ~n11460;
  assign n11462 = n11461 ^ x506;
  assign n11463 = n11462 ^ n11435;
  assign n11464 = n11436 & ~n11463;
  assign n11465 = n11464 ^ x505;
  assign n11466 = n11465 ^ n11433;
  assign n11467 = n11434 & ~n11466;
  assign n11468 = n11467 ^ x504;
  assign n11469 = n11468 ^ n11431;
  assign n11470 = n11432 & ~n11469;
  assign n11471 = n11470 ^ x503;
  assign n11472 = n11471 ^ n11429;
  assign n11473 = ~n11430 & n11472;
  assign n11474 = n11473 ^ x502;
  assign n11475 = n11474 ^ n11427;
  assign n11476 = n11428 & ~n11475;
  assign n11477 = n11476 ^ x501;
  assign n11803 = n11494 ^ n11477;
  assign n11804 = n11802 & ~n11803;
  assign n11805 = n11804 ^ x500;
  assign n11806 = n11805 ^ n11800;
  assign n11807 = n11801 & ~n11806;
  assign n11808 = n11807 ^ x499;
  assign n11809 = n11808 ^ n11798;
  assign n11810 = n11799 & ~n11809;
  assign n11811 = n11810 ^ x498;
  assign n11812 = n11811 ^ n11796;
  assign n11813 = n11797 & ~n11812;
  assign n11814 = n11813 ^ x497;
  assign n11815 = n11814 ^ n11794;
  assign n11816 = ~n11795 & n11815;
  assign n11817 = n11816 ^ x496;
  assign n11819 = n11818 ^ n11817;
  assign n11820 = n11818 ^ x495;
  assign n11821 = ~n11819 & n11820;
  assign n11822 = n11821 ^ x495;
  assign n11823 = n11822 ^ n11792;
  assign n11824 = ~n11793 & n11823;
  assign n11825 = n11824 ^ x494;
  assign n11725 = ~n11713 & ~n11724;
  assign n11671 = n11670 ^ n11641;
  assign n11672 = ~n11642 & n11671;
  assign n11673 = n11672 ^ n9133;
  assign n11545 = n11544 ^ n11541;
  assign n11592 = n11591 ^ n11541;
  assign n11593 = n11545 & ~n11592;
  assign n11594 = n11593 ^ n11544;
  assign n11537 = n10289 ^ n9101;
  assign n11538 = ~n10728 & ~n11537;
  assign n11539 = n11538 ^ n9101;
  assign n11637 = n11594 ^ n11539;
  assign n11496 = n11217 ^ x466;
  assign n11497 = n11496 ^ n11167;
  assign n11638 = n11637 ^ n11497;
  assign n11639 = n11638 ^ n9126;
  assign n11712 = n11673 ^ n11639;
  assign n11790 = n11725 ^ n11712;
  assign n11791 = n11790 ^ x493;
  assign n12098 = n11825 ^ n11791;
  assign n12102 = n12101 ^ n12098;
  assign n11749 = n11246 ^ n11152;
  assign n12105 = n10698 ^ n10602;
  assign n12106 = n11749 & ~n12105;
  assign n12107 = n12106 ^ n10602;
  assign n12103 = n11822 ^ x494;
  assign n12104 = n12103 ^ n11792;
  assign n12108 = n12107 ^ n12104;
  assign n11704 = n11243 ^ x458;
  assign n11705 = n11704 ^ n11153;
  assign n12110 = n10700 ^ n10569;
  assign n12111 = ~n11705 & n12110;
  assign n12112 = n12111 ^ n10569;
  assign n12109 = n11819 ^ x495;
  assign n12113 = n12112 ^ n12109;
  assign n11619 = n11240 ^ n11156;
  assign n12116 = n10705 ^ n10537;
  assign n12117 = ~n11619 & n12116;
  assign n12118 = n12117 ^ n10537;
  assign n12114 = n11814 ^ x496;
  assign n12115 = n12114 ^ n11794;
  assign n12119 = n12118 ^ n12115;
  assign n11507 = n11237 ^ x460;
  assign n11508 = n11507 ^ n11157;
  assign n12121 = n10711 ^ n10389;
  assign n12122 = n11508 & n12121;
  assign n12123 = n12122 ^ n10389;
  assign n12120 = n11811 ^ n11797;
  assign n12124 = n12123 ^ n12120;
  assign n12128 = n11808 ^ x498;
  assign n12129 = n12128 ^ n11798;
  assign n11513 = n11234 ^ n11160;
  assign n12125 = n10717 ^ n10289;
  assign n12126 = ~n11513 & n12125;
  assign n12127 = n12126 ^ n10289;
  assign n12130 = n12129 ^ n12127;
  assign n12134 = n11805 ^ n11801;
  assign n11518 = n11231 ^ x462;
  assign n11519 = n11518 ^ n11161;
  assign n12131 = n10723 ^ n10155;
  assign n12132 = ~n11519 & ~n12131;
  assign n12133 = n12132 ^ n10155;
  assign n12135 = n12134 ^ n12133;
  assign n11524 = n11228 ^ x463;
  assign n12136 = n10728 ^ n10160;
  assign n12137 = n11524 & ~n12136;
  assign n12138 = n12137 ^ n10160;
  assign n11478 = n11477 ^ x500;
  assign n11495 = n11494 ^ n11478;
  assign n12139 = n12138 ^ n11495;
  assign n11526 = n11223 ^ x464;
  assign n11527 = n11526 ^ n11163;
  assign n12140 = n10734 ^ n10275;
  assign n12141 = ~n11527 & n12140;
  assign n12142 = n12141 ^ n10275;
  assign n12040 = n11474 ^ n11428;
  assign n12143 = n12142 ^ n12040;
  assign n11532 = n11220 ^ n11166;
  assign n12144 = n10735 ^ n10165;
  assign n12145 = n11532 & n12144;
  assign n12146 = n12145 ^ n10165;
  assign n12046 = n11471 ^ n11430;
  assign n12147 = n12146 ^ n12046;
  assign n12148 = n10741 ^ n10171;
  assign n12149 = ~n11497 & ~n12148;
  assign n12150 = n12149 ^ n10171;
  assign n12052 = n11468 ^ x503;
  assign n12053 = n12052 ^ n11431;
  assign n12151 = n12150 ^ n12053;
  assign n12152 = n10746 ^ n10176;
  assign n12153 = n11541 & n12152;
  assign n12154 = n12153 ^ n10176;
  assign n12060 = n11465 ^ x504;
  assign n12061 = n12060 ^ n11433;
  assign n12155 = n12154 ^ n12061;
  assign n12159 = n11462 ^ n11436;
  assign n12156 = n10752 ^ n10182;
  assign n12157 = n11550 & n12156;
  assign n12158 = n12157 ^ n10182;
  assign n12160 = n12159 ^ n12158;
  assign n12161 = n10757 ^ n10187;
  assign n12162 = ~n11555 & ~n12161;
  assign n12163 = n12162 ^ n10187;
  assign n12067 = n11459 ^ x506;
  assign n12068 = n12067 ^ n11437;
  assign n12164 = n12163 ^ n12068;
  assign n12168 = n11456 ^ n11440;
  assign n12165 = n10763 ^ n10190;
  assign n12166 = ~n11557 & ~n12165;
  assign n12167 = n12166 ^ n10190;
  assign n12169 = n12168 ^ n12167;
  assign n12173 = n11453 ^ x508;
  assign n12174 = n12173 ^ n11441;
  assign n12170 = n10768 ^ n10141;
  assign n12171 = ~n11566 & ~n12170;
  assign n12172 = n12171 ^ n10141;
  assign n12175 = n12174 ^ n12172;
  assign n12179 = n11450 ^ x509;
  assign n12180 = n12179 ^ n11443;
  assign n12176 = n10776 ^ n10199;
  assign n12177 = n11572 & ~n12176;
  assign n12178 = n12177 ^ n10199;
  assign n12181 = n12180 ^ n12178;
  assign n12030 = n11447 ^ n11446;
  assign n12027 = n10204 ^ n10140;
  assign n12028 = n11488 & ~n12027;
  assign n12029 = n12028 ^ n10204;
  assign n12031 = n12030 ^ n12029;
  assign n11987 = n10672 ^ n10210;
  assign n11988 = n11403 & ~n11987;
  assign n11989 = n11988 ^ n10210;
  assign n11991 = n11990 ^ n11989;
  assign n11960 = n10046 ^ n9206;
  assign n11961 = ~n10840 & ~n11960;
  assign n11962 = n11961 ^ n9206;
  assign n11959 = n11258 ^ n11144;
  assign n11963 = n11962 ^ n11959;
  assign n11964 = n11963 ^ n8786;
  assign n11870 = n11252 ^ n11148;
  assign n11761 = n9975 ^ n9424;
  assign n11762 = n10574 & ~n11761;
  assign n11763 = n11762 ^ n9424;
  assign n11766 = n11765 ^ n11763;
  assign n11746 = n9997 ^ n9446;
  assign n11747 = n10542 & ~n11746;
  assign n11748 = n11747 ^ n9446;
  assign n11750 = n11749 ^ n11748;
  assign n11701 = n9981 ^ n9430;
  assign n11702 = ~n11286 & n11701;
  assign n11703 = n11702 ^ n9430;
  assign n11706 = n11705 ^ n11703;
  assign n11616 = n9987 ^ n9436;
  assign n11617 = n11077 & n11616;
  assign n11618 = n11617 ^ n9436;
  assign n11620 = n11619 ^ n11618;
  assign n11504 = n10712 ^ n9963;
  assign n11505 = n10698 & ~n11504;
  assign n11506 = n11505 ^ n9963;
  assign n11509 = n11508 ^ n11506;
  assign n11510 = n10656 ^ n9796;
  assign n11511 = n10700 & n11510;
  assign n11512 = n11511 ^ n9796;
  assign n11514 = n11513 ^ n11512;
  assign n11515 = n10602 ^ n9776;
  assign n11516 = ~n10705 & ~n11515;
  assign n11517 = n11516 ^ n9776;
  assign n11520 = n11519 ^ n11517;
  assign n11521 = n10569 ^ n9700;
  assign n11522 = ~n10711 & n11521;
  assign n11523 = n11522 ^ n9700;
  assign n11525 = n11524 ^ n11523;
  assign n11528 = n10537 ^ n9538;
  assign n11529 = n10717 & ~n11528;
  assign n11530 = n11529 ^ n9538;
  assign n11531 = n11530 ^ n11527;
  assign n11533 = n10389 ^ n9094;
  assign n11534 = n10723 & n11533;
  assign n11535 = n11534 ^ n9094;
  assign n11536 = n11535 ^ n11532;
  assign n11540 = n11539 ^ n11497;
  assign n11595 = n11594 ^ n11497;
  assign n11596 = n11540 & n11595;
  assign n11597 = n11596 ^ n11539;
  assign n11598 = n11597 ^ n11532;
  assign n11599 = ~n11536 & n11598;
  assign n11600 = n11599 ^ n11535;
  assign n11601 = n11600 ^ n11527;
  assign n11602 = ~n11531 & ~n11601;
  assign n11603 = n11602 ^ n11530;
  assign n11604 = n11603 ^ n11524;
  assign n11605 = n11525 & ~n11604;
  assign n11606 = n11605 ^ n11523;
  assign n11607 = n11606 ^ n11519;
  assign n11608 = ~n11520 & n11607;
  assign n11609 = n11608 ^ n11517;
  assign n11610 = n11609 ^ n11513;
  assign n11611 = ~n11514 & n11610;
  assign n11612 = n11611 ^ n11512;
  assign n11613 = n11612 ^ n11508;
  assign n11614 = ~n11509 & ~n11613;
  assign n11615 = n11614 ^ n11506;
  assign n11698 = n11619 ^ n11615;
  assign n11699 = n11620 & ~n11698;
  assign n11700 = n11699 ^ n11618;
  assign n11743 = n11705 ^ n11700;
  assign n11744 = n11706 & ~n11743;
  assign n11745 = n11744 ^ n11703;
  assign n11758 = n11749 ^ n11745;
  assign n11759 = n11750 & n11758;
  assign n11760 = n11759 ^ n11748;
  assign n11867 = n11765 ^ n11760;
  assign n11868 = ~n11766 & ~n11867;
  assign n11869 = n11868 ^ n11763;
  assign n11871 = n11870 ^ n11869;
  assign n11864 = n9969 ^ n9418;
  assign n11865 = n10607 & ~n11864;
  assign n11866 = n11865 ^ n9418;
  assign n11913 = n11870 ^ n11866;
  assign n11914 = ~n11871 & ~n11913;
  assign n11915 = n11914 ^ n11866;
  assign n11911 = n11255 ^ x454;
  assign n11912 = n11911 ^ n11145;
  assign n11916 = n11915 ^ n11912;
  assign n11908 = n10011 ^ n9210;
  assign n11909 = n10665 & n11908;
  assign n11910 = n11909 ^ n9210;
  assign n11956 = n11912 ^ n11910;
  assign n11957 = ~n11916 & n11956;
  assign n11958 = n11957 ^ n11910;
  assign n11965 = n11964 ^ n11958;
  assign n11707 = n11706 ^ n11700;
  assign n11708 = n11707 ^ n8586;
  assign n11621 = n11620 ^ n11615;
  assign n11622 = n11621 ^ n8589;
  assign n11623 = n11612 ^ n11509;
  assign n11624 = n11623 ^ n9095;
  assign n11625 = n11609 ^ n11514;
  assign n11626 = n11625 ^ n9103;
  assign n11627 = n11606 ^ n11520;
  assign n11628 = n11627 ^ n9110;
  assign n11629 = n11603 ^ n11525;
  assign n11630 = n11629 ^ n9117;
  assign n11631 = n11600 ^ n11530;
  assign n11632 = n11631 ^ n11527;
  assign n11633 = n11632 ^ n9225;
  assign n11634 = n11597 ^ n11535;
  assign n11635 = n11634 ^ n11532;
  assign n11636 = n11635 ^ n9231;
  assign n11674 = n11673 ^ n11638;
  assign n11675 = ~n11639 & n11674;
  assign n11676 = n11675 ^ n9126;
  assign n11677 = n11676 ^ n11635;
  assign n11678 = n11636 & n11677;
  assign n11679 = n11678 ^ n9231;
  assign n11680 = n11679 ^ n11632;
  assign n11681 = n11633 & ~n11680;
  assign n11682 = n11681 ^ n9225;
  assign n11683 = n11682 ^ n11629;
  assign n11684 = ~n11630 & ~n11683;
  assign n11685 = n11684 ^ n9117;
  assign n11686 = n11685 ^ n11627;
  assign n11687 = ~n11628 & ~n11686;
  assign n11688 = n11687 ^ n9110;
  assign n11689 = n11688 ^ n11625;
  assign n11690 = ~n11626 & n11689;
  assign n11691 = n11690 ^ n9103;
  assign n11692 = n11691 ^ n11623;
  assign n11693 = n11624 & n11692;
  assign n11694 = n11693 ^ n9095;
  assign n11695 = n11694 ^ n11621;
  assign n11696 = n11622 & ~n11695;
  assign n11697 = n11696 ^ n8589;
  assign n11709 = n11708 ^ n11697;
  assign n11710 = n11682 ^ n11630;
  assign n11711 = n11679 ^ n11633;
  assign n11726 = n11712 & ~n11725;
  assign n11727 = n11676 ^ n11636;
  assign n11728 = n11726 & ~n11727;
  assign n11729 = n11711 & n11728;
  assign n11730 = ~n11710 & n11729;
  assign n11731 = n11685 ^ n11628;
  assign n11732 = n11730 & n11731;
  assign n11733 = n11688 ^ n11626;
  assign n11734 = ~n11732 & n11733;
  assign n11735 = n11691 ^ n11624;
  assign n11736 = ~n11734 & n11735;
  assign n11737 = n11694 ^ n11622;
  assign n11738 = ~n11736 & n11737;
  assign n11739 = n11709 & ~n11738;
  assign n11751 = n11750 ^ n11745;
  assign n11752 = n11751 ^ n8622;
  assign n11740 = n11707 ^ n11697;
  assign n11741 = ~n11708 & ~n11740;
  assign n11742 = n11741 ^ n8586;
  assign n11753 = n11752 ^ n11742;
  assign n11754 = ~n11739 & ~n11753;
  assign n11767 = n11766 ^ n11760;
  assign n11768 = n11767 ^ n8667;
  assign n11755 = n11751 ^ n11742;
  assign n11756 = n11752 & n11755;
  assign n11757 = n11756 ^ n8622;
  assign n11769 = n11768 ^ n11757;
  assign n11860 = n11754 & ~n11769;
  assign n11872 = n11871 ^ n11866;
  assign n11873 = n11872 ^ n8725;
  assign n11861 = n11767 ^ n11757;
  assign n11862 = ~n11768 & ~n11861;
  assign n11863 = n11862 ^ n8667;
  assign n11874 = n11873 ^ n11863;
  assign n11903 = ~n11860 & ~n11874;
  assign n11917 = n11916 ^ n11910;
  assign n11904 = n11872 ^ n11863;
  assign n11905 = ~n11873 & ~n11904;
  assign n11906 = n11905 ^ n8725;
  assign n11907 = n11906 ^ n8791;
  assign n11918 = n11917 ^ n11907;
  assign n11955 = ~n11903 & ~n11918;
  assign n11966 = n11965 ^ n11955;
  assign n11951 = n11917 ^ n8791;
  assign n11952 = n11917 ^ n11906;
  assign n11953 = ~n11951 & n11952;
  assign n11954 = n11953 ^ n8791;
  assign n11967 = n11966 ^ n11954;
  assign n11919 = n11918 ^ n11903;
  assign n11946 = n11919 ^ x481;
  assign n11875 = n11874 ^ n11860;
  assign n11898 = n11875 ^ x482;
  assign n11770 = n11769 ^ n11754;
  assign n11771 = n11770 ^ x483;
  assign n11772 = n11753 ^ n11739;
  assign n11773 = n11772 ^ x484;
  assign n11774 = n11738 ^ n11709;
  assign n11775 = n11774 ^ x485;
  assign n11776 = n11737 ^ n11736;
  assign n11777 = n11776 ^ x486;
  assign n11778 = n11735 ^ n11734;
  assign n11779 = n11778 ^ x487;
  assign n11780 = n11733 ^ n11732;
  assign n11781 = n11780 ^ x488;
  assign n11782 = n11731 ^ n11730;
  assign n11783 = n11782 ^ x489;
  assign n11784 = n11729 ^ n11710;
  assign n11785 = n11784 ^ x490;
  assign n11786 = n11728 ^ n11711;
  assign n11787 = n11786 ^ x491;
  assign n11788 = n11727 ^ n11726;
  assign n11789 = n11788 ^ x492;
  assign n11826 = n11825 ^ n11790;
  assign n11827 = ~n11791 & n11826;
  assign n11828 = n11827 ^ x493;
  assign n11829 = n11828 ^ n11788;
  assign n11830 = ~n11789 & n11829;
  assign n11831 = n11830 ^ x492;
  assign n11832 = n11831 ^ n11786;
  assign n11833 = n11787 & ~n11832;
  assign n11834 = n11833 ^ x491;
  assign n11835 = n11834 ^ n11784;
  assign n11836 = ~n11785 & n11835;
  assign n11837 = n11836 ^ x490;
  assign n11838 = n11837 ^ n11782;
  assign n11839 = n11783 & ~n11838;
  assign n11840 = n11839 ^ x489;
  assign n11841 = n11840 ^ n11780;
  assign n11842 = n11781 & ~n11841;
  assign n11843 = n11842 ^ x488;
  assign n11844 = n11843 ^ n11778;
  assign n11845 = ~n11779 & n11844;
  assign n11846 = n11845 ^ x487;
  assign n11847 = n11846 ^ n11776;
  assign n11848 = n11777 & ~n11847;
  assign n11849 = n11848 ^ x486;
  assign n11850 = n11849 ^ n11774;
  assign n11851 = ~n11775 & n11850;
  assign n11852 = n11851 ^ x485;
  assign n11853 = n11852 ^ n11772;
  assign n11854 = ~n11773 & n11853;
  assign n11855 = n11854 ^ x484;
  assign n11856 = n11855 ^ n11770;
  assign n11857 = n11771 & ~n11856;
  assign n11858 = n11857 ^ x483;
  assign n11899 = n11875 ^ n11858;
  assign n11900 = n11898 & ~n11899;
  assign n11901 = n11900 ^ x482;
  assign n11947 = n11919 ^ n11901;
  assign n11948 = ~n11946 & n11947;
  assign n11949 = n11948 ^ x481;
  assign n11950 = n11949 ^ x480;
  assign n11968 = n11967 ^ n11950;
  assign n11943 = n10679 ^ n10216;
  assign n11944 = ~n11345 & ~n11943;
  assign n11945 = n11944 ^ n10216;
  assign n11969 = n11968 ^ n11945;
  assign n11902 = n11901 ^ x481;
  assign n11920 = n11919 ^ n11902;
  assign n11895 = n10686 ^ n10222;
  assign n11896 = ~n10670 & ~n11895;
  assign n11897 = n11896 ^ n10222;
  assign n11921 = n11920 ^ n11897;
  assign n11859 = n11858 ^ x482;
  assign n11876 = n11875 ^ n11859;
  assign n11501 = n10691 ^ n10227;
  assign n11502 = n10676 & ~n11501;
  assign n11503 = n11502 ^ n10227;
  assign n11877 = n11876 ^ n11503;
  assign n11881 = n11855 ^ n11771;
  assign n11878 = n10802 ^ n10132;
  assign n11879 = n10678 & n11878;
  assign n11880 = n11879 ^ n10132;
  assign n11882 = n11881 ^ n11880;
  assign n11883 = n10804 ^ n10105;
  assign n11884 = ~n10684 & ~n11883;
  assign n11885 = n11884 ^ n10105;
  assign n11886 = n11852 ^ x484;
  assign n11887 = n11886 ^ n11772;
  assign n11888 = n11885 & ~n11887;
  assign n11889 = n11888 ^ n11881;
  assign n11890 = n11882 & n11889;
  assign n11891 = n11890 ^ n11888;
  assign n11892 = n11891 ^ n11876;
  assign n11893 = n11877 & ~n11892;
  assign n11894 = n11893 ^ n11503;
  assign n11940 = n11920 ^ n11894;
  assign n11941 = n11921 & n11940;
  assign n11942 = n11941 ^ n11897;
  assign n11984 = n11968 ^ n11942;
  assign n11985 = n11969 & ~n11984;
  assign n11986 = n11985 ^ n11945;
  assign n12024 = n11990 ^ n11986;
  assign n12025 = ~n11991 & n12024;
  assign n12026 = n12025 ^ n11989;
  assign n12182 = n12030 ^ n12026;
  assign n12183 = ~n12031 & ~n12182;
  assign n12184 = n12183 ^ n12029;
  assign n12185 = n12184 ^ n12180;
  assign n12186 = ~n12181 & ~n12185;
  assign n12187 = n12186 ^ n12178;
  assign n12188 = n12187 ^ n12174;
  assign n12189 = ~n12175 & ~n12188;
  assign n12190 = n12189 ^ n12172;
  assign n12191 = n12190 ^ n12168;
  assign n12192 = ~n12169 & n12191;
  assign n12193 = n12192 ^ n12167;
  assign n12194 = n12193 ^ n12068;
  assign n12195 = ~n12164 & ~n12194;
  assign n12196 = n12195 ^ n12163;
  assign n12197 = n12196 ^ n12159;
  assign n12198 = n12160 & n12197;
  assign n12199 = n12198 ^ n12158;
  assign n12200 = n12199 ^ n12061;
  assign n12201 = ~n12155 & ~n12200;
  assign n12202 = n12201 ^ n12154;
  assign n12203 = n12202 ^ n12053;
  assign n12204 = ~n12151 & n12203;
  assign n12205 = n12204 ^ n12150;
  assign n12206 = n12205 ^ n12046;
  assign n12207 = n12147 & ~n12206;
  assign n12208 = n12207 ^ n12146;
  assign n12209 = n12208 ^ n12040;
  assign n12210 = n12143 & n12209;
  assign n12211 = n12210 ^ n12142;
  assign n12212 = n12211 ^ n11495;
  assign n12213 = n12139 & ~n12212;
  assign n12214 = n12213 ^ n12138;
  assign n12215 = n12214 ^ n12134;
  assign n12216 = ~n12135 & ~n12215;
  assign n12217 = n12216 ^ n12133;
  assign n12218 = n12217 ^ n12129;
  assign n12219 = n12130 & n12218;
  assign n12220 = n12219 ^ n12127;
  assign n12221 = n12220 ^ n12120;
  assign n12222 = ~n12124 & ~n12221;
  assign n12223 = n12222 ^ n12123;
  assign n12224 = n12223 ^ n12115;
  assign n12225 = n12119 & ~n12224;
  assign n12226 = n12225 ^ n12118;
  assign n12227 = n12226 ^ n12109;
  assign n12228 = n12113 & n12227;
  assign n12229 = n12228 ^ n12112;
  assign n12230 = n12229 ^ n12104;
  assign n12231 = n12108 & n12230;
  assign n12232 = n12231 ^ n12107;
  assign n12233 = n12232 ^ n12098;
  assign n12234 = ~n12102 & ~n12233;
  assign n12235 = n12234 ^ n12101;
  assign n12094 = n11286 ^ n10712;
  assign n12095 = ~n11870 & ~n12094;
  assign n12096 = n12095 ^ n10712;
  assign n12092 = n11828 ^ x492;
  assign n12093 = n12092 ^ n11788;
  assign n12097 = n12096 ^ n12093;
  assign n12262 = n12235 ^ n12097;
  assign n12263 = n12262 ^ n9963;
  assign n12264 = n12232 ^ n12102;
  assign n12265 = n12264 ^ n9796;
  assign n12266 = n12229 ^ n12108;
  assign n12267 = n12266 ^ n9776;
  assign n12268 = n12226 ^ n12113;
  assign n12269 = n12268 ^ n9700;
  assign n12270 = n12223 ^ n12119;
  assign n12271 = n12270 ^ n9538;
  assign n12272 = n12220 ^ n12124;
  assign n12273 = n12272 ^ n9094;
  assign n12274 = n12217 ^ n12130;
  assign n12275 = n12274 ^ n9101;
  assign n12276 = n12214 ^ n12133;
  assign n12277 = n12276 ^ n12134;
  assign n12278 = n12277 ^ n9109;
  assign n12279 = n12211 ^ n12138;
  assign n12280 = n12279 ^ n11495;
  assign n12281 = n12280 ^ n9115;
  assign n12282 = n12208 ^ n12142;
  assign n12283 = n12282 ^ n12040;
  assign n12284 = n12283 ^ n9122;
  assign n12285 = n12205 ^ n12147;
  assign n12286 = n12285 ^ n9123;
  assign n12287 = n12202 ^ n12151;
  assign n12288 = n12287 ^ n9125;
  assign n12289 = n12199 ^ n12155;
  assign n12290 = n12289 ^ n9131;
  assign n12291 = n12196 ^ n12160;
  assign n12292 = n12291 ^ n9143;
  assign n12293 = n12193 ^ n12164;
  assign n12294 = n12293 ^ n9150;
  assign n12295 = n12190 ^ n12169;
  assign n12296 = n12295 ^ n9156;
  assign n12297 = n12187 ^ n12175;
  assign n12298 = n12297 ^ n9161;
  assign n12299 = n12184 ^ n12181;
  assign n12300 = n12299 ^ n9166;
  assign n12032 = n12031 ^ n12026;
  assign n12033 = n12032 ^ n9172;
  assign n11992 = n11991 ^ n11986;
  assign n11993 = n11992 ^ n9178;
  assign n11970 = n11969 ^ n11942;
  assign n11971 = n11970 ^ n9180;
  assign n11922 = n11921 ^ n11894;
  assign n11923 = n11922 ^ n9189;
  assign n11924 = n11891 ^ n11877;
  assign n11925 = n11924 ^ n8733;
  assign n11926 = n11887 ^ n11885;
  assign n11927 = ~n9201 & ~n11926;
  assign n11928 = n11927 ^ n9199;
  assign n11929 = n11888 ^ n11880;
  assign n11930 = n11929 ^ n11881;
  assign n11931 = n11930 ^ n11927;
  assign n11932 = ~n11928 & n11931;
  assign n11933 = n11932 ^ n9199;
  assign n11934 = n11933 ^ n11924;
  assign n11935 = n11925 & n11934;
  assign n11936 = n11935 ^ n8733;
  assign n11937 = n11936 ^ n11922;
  assign n11938 = ~n11923 & ~n11937;
  assign n11939 = n11938 ^ n9189;
  assign n11981 = n11970 ^ n11939;
  assign n11982 = ~n11971 & ~n11981;
  assign n11983 = n11982 ^ n9180;
  assign n12021 = n11992 ^ n11983;
  assign n12022 = ~n11993 & ~n12021;
  assign n12023 = n12022 ^ n9178;
  assign n12301 = n12032 ^ n12023;
  assign n12302 = ~n12033 & n12301;
  assign n12303 = n12302 ^ n9172;
  assign n12304 = n12303 ^ n12299;
  assign n12305 = n12300 & ~n12304;
  assign n12306 = n12305 ^ n9166;
  assign n12307 = n12306 ^ n12297;
  assign n12308 = n12298 & n12307;
  assign n12309 = n12308 ^ n9161;
  assign n12310 = n12309 ^ n12295;
  assign n12311 = n12296 & n12310;
  assign n12312 = n12311 ^ n9156;
  assign n12313 = n12312 ^ n12293;
  assign n12314 = n12294 & ~n12313;
  assign n12315 = n12314 ^ n9150;
  assign n12316 = n12315 ^ n12291;
  assign n12317 = n12292 & ~n12316;
  assign n12318 = n12317 ^ n9143;
  assign n12319 = n12318 ^ n12289;
  assign n12320 = n12290 & ~n12319;
  assign n12321 = n12320 ^ n9131;
  assign n12322 = n12321 ^ n12287;
  assign n12323 = ~n12288 & n12322;
  assign n12324 = n12323 ^ n9125;
  assign n12325 = n12324 ^ n12285;
  assign n12326 = n12286 & ~n12325;
  assign n12327 = n12326 ^ n9123;
  assign n12328 = n12327 ^ n12283;
  assign n12329 = n12284 & ~n12328;
  assign n12330 = n12329 ^ n9122;
  assign n12331 = n12330 ^ n12280;
  assign n12332 = n12281 & n12331;
  assign n12333 = n12332 ^ n9115;
  assign n12334 = n12333 ^ n12277;
  assign n12335 = ~n12278 & n12334;
  assign n12336 = n12335 ^ n9109;
  assign n12337 = n12336 ^ n12274;
  assign n12338 = n12275 & n12337;
  assign n12339 = n12338 ^ n9101;
  assign n12340 = n12339 ^ n12272;
  assign n12341 = n12273 & ~n12340;
  assign n12342 = n12341 ^ n9094;
  assign n12343 = n12342 ^ n12270;
  assign n12344 = ~n12271 & ~n12343;
  assign n12345 = n12344 ^ n9538;
  assign n12346 = n12345 ^ n12268;
  assign n12347 = ~n12269 & n12346;
  assign n12348 = n12347 ^ n9700;
  assign n12349 = n12348 ^ n12266;
  assign n12350 = n12267 & ~n12349;
  assign n12351 = n12350 ^ n9776;
  assign n12352 = n12351 ^ n12264;
  assign n12353 = n12265 & ~n12352;
  assign n12354 = n12353 ^ n9796;
  assign n12355 = n12354 ^ n12262;
  assign n12356 = n12263 & n12355;
  assign n12357 = n12356 ^ n9963;
  assign n12236 = n12235 ^ n12093;
  assign n12237 = ~n12097 & n12236;
  assign n12238 = n12237 ^ n12096;
  assign n12088 = n10542 ^ n9987;
  assign n12089 = n11912 & ~n12088;
  assign n12090 = n12089 ^ n9987;
  assign n12086 = n11831 ^ x491;
  assign n12087 = n12086 ^ n11786;
  assign n12091 = n12090 ^ n12087;
  assign n12260 = n12238 ^ n12091;
  assign n12261 = n12260 ^ n9436;
  assign n12384 = n12357 ^ n12261;
  assign n12385 = n12324 ^ n12286;
  assign n12386 = n12312 ^ n12294;
  assign n12034 = n12033 ^ n12023;
  assign n11972 = n11971 ^ n11939;
  assign n11973 = n11936 ^ n11923;
  assign n11974 = n11933 ^ n11925;
  assign n11975 = n11926 ^ n9201;
  assign n11976 = n11930 ^ n11928;
  assign n11977 = n11975 & n11976;
  assign n11978 = ~n11974 & n11977;
  assign n11979 = n11973 & ~n11978;
  assign n11980 = ~n11972 & n11979;
  assign n11994 = n11993 ^ n11983;
  assign n12035 = ~n11980 & ~n11994;
  assign n12387 = n12034 & n12035;
  assign n12388 = n12303 ^ n12300;
  assign n12389 = ~n12387 & n12388;
  assign n12390 = n12306 ^ n12298;
  assign n12391 = n12389 & n12390;
  assign n12392 = n12309 ^ n12296;
  assign n12393 = ~n12391 & n12392;
  assign n12394 = ~n12386 & n12393;
  assign n12395 = n12315 ^ n12292;
  assign n12396 = ~n12394 & n12395;
  assign n12397 = n12318 ^ n12290;
  assign n12398 = n12396 & n12397;
  assign n12399 = n12321 ^ n12288;
  assign n12400 = n12398 & ~n12399;
  assign n12401 = n12385 & n12400;
  assign n12402 = n12327 ^ n12284;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = n12330 ^ n12281;
  assign n12405 = n12403 & ~n12404;
  assign n12406 = n12333 ^ n12278;
  assign n12407 = ~n12405 & n12406;
  assign n12408 = n12336 ^ n12275;
  assign n12409 = ~n12407 & n12408;
  assign n12410 = n12339 ^ n12273;
  assign n12411 = n12409 & ~n12410;
  assign n12412 = n12342 ^ n12271;
  assign n12413 = n12411 & n12412;
  assign n12414 = n12345 ^ n12269;
  assign n12415 = n12413 & ~n12414;
  assign n12416 = n12348 ^ n12267;
  assign n12417 = n12415 & n12416;
  assign n12418 = n12351 ^ n12265;
  assign n12419 = ~n12417 & ~n12418;
  assign n12420 = n12354 ^ n12263;
  assign n12421 = ~n12419 & n12420;
  assign n12422 = n12384 & ~n12421;
  assign n12358 = n12357 ^ n12260;
  assign n12359 = n12261 & ~n12358;
  assign n12360 = n12359 ^ n9436;
  assign n12239 = n12238 ^ n12087;
  assign n12240 = ~n12091 & ~n12239;
  assign n12241 = n12240 ^ n12090;
  assign n12082 = n10574 ^ n9981;
  assign n12083 = n11959 & ~n12082;
  assign n12084 = n12083 ^ n9981;
  assign n12257 = n12241 ^ n12084;
  assign n12080 = n11834 ^ x490;
  assign n12081 = n12080 ^ n11784;
  assign n12258 = n12257 ^ n12081;
  assign n12259 = n12258 ^ n9430;
  assign n12383 = n12360 ^ n12259;
  assign n12537 = n12422 ^ n12383;
  assign n12433 = n12421 ^ n12384;
  assign n2265 = x263 ^ x71;
  assign n2266 = n2265 ^ x423;
  assign n2267 = n2266 ^ x7;
  assign n12434 = n12433 ^ n2267;
  assign n12435 = n12420 ^ n12419;
  assign n12436 = n12435 ^ n1213;
  assign n12437 = n12418 ^ n12417;
  assign n12438 = n12437 ^ n1207;
  assign n12523 = n12416 ^ n12415;
  assign n12439 = n12414 ^ n12413;
  assign n12440 = n12439 ^ n896;
  assign n12515 = n12412 ^ n12411;
  assign n12441 = n12410 ^ n12409;
  assign n12442 = n12441 ^ n799;
  assign n12443 = n12408 ^ n12407;
  assign n12444 = n12443 ^ n787;
  assign n12445 = n12406 ^ n12405;
  assign n12446 = n12445 ^ n781;
  assign n12501 = n12404 ^ n12403;
  assign n12447 = n12402 ^ n12401;
  assign n12451 = n12450 ^ n12447;
  assign n12493 = n12400 ^ n12385;
  assign n12452 = n12399 ^ n12398;
  assign n12453 = n12452 ^ n572;
  assign n12485 = n12397 ^ n12396;
  assign n12454 = n12395 ^ n12394;
  assign n12458 = n12457 ^ n12454;
  assign n12477 = n12393 ^ n12386;
  assign n12459 = n12392 ^ n12391;
  assign n12460 = n12459 ^ n2170;
  assign n12469 = n12390 ^ n12389;
  assign n12461 = n12388 ^ n12387;
  assign n12462 = n12461 ^ n1889;
  assign n12036 = n12035 ^ n12034;
  assign n12037 = n12036 ^ n1871;
  assign n11995 = n11994 ^ n11980;
  assign n11996 = n11995 ^ n1691;
  assign n11997 = n11979 ^ n11972;
  assign n11998 = n11997 ^ n1855;
  assign n12010 = n11978 ^ n11973;
  assign n11999 = n11977 ^ n11974;
  assign n12000 = n11999 ^ n1444;
  assign n12001 = n1470 & ~n11975;
  assign n12002 = n12001 ^ n1419;
  assign n12003 = n11976 ^ n11975;
  assign n12004 = n12003 ^ n12001;
  assign n12005 = n12002 & ~n12004;
  assign n12006 = n12005 ^ n1419;
  assign n12007 = n12006 ^ n11999;
  assign n12008 = ~n12000 & n12007;
  assign n12009 = n12008 ^ n1444;
  assign n12011 = n12010 ^ n12009;
  assign n12012 = n12010 ^ n1595;
  assign n12013 = ~n12011 & n12012;
  assign n12014 = n12013 ^ n1595;
  assign n12015 = n12014 ^ n11997;
  assign n12016 = n11998 & ~n12015;
  assign n12017 = n12016 ^ n1855;
  assign n12018 = n12017 ^ n11995;
  assign n12019 = n11996 & ~n12018;
  assign n12020 = n12019 ^ n1691;
  assign n12463 = n12036 ^ n12020;
  assign n12464 = n12037 & ~n12463;
  assign n12465 = n12464 ^ n1871;
  assign n12466 = n12465 ^ n12461;
  assign n12467 = n12462 & ~n12466;
  assign n12468 = n12467 ^ n1889;
  assign n12470 = n12469 ^ n12468;
  assign n12471 = n12469 ^ n2011;
  assign n12472 = n12470 & ~n12471;
  assign n12473 = n12472 ^ n2011;
  assign n12474 = n12473 ^ n12459;
  assign n12475 = ~n12460 & n12474;
  assign n12476 = n12475 ^ n2170;
  assign n12478 = n12477 ^ n12476;
  assign n12479 = n12477 ^ n2162;
  assign n12480 = n12478 & ~n12479;
  assign n12481 = n12480 ^ n2162;
  assign n12482 = n12481 ^ n12454;
  assign n12483 = n12458 & ~n12482;
  assign n12484 = n12483 ^ n12457;
  assign n12486 = n12485 ^ n12484;
  assign n12487 = n12485 ^ n601;
  assign n12488 = n12486 & ~n12487;
  assign n12489 = n12488 ^ n601;
  assign n12490 = n12489 ^ n12452;
  assign n12491 = n12453 & ~n12490;
  assign n12492 = n12491 ^ n572;
  assign n12494 = n12493 ^ n12492;
  assign n12495 = n12493 ^ n522;
  assign n12496 = n12494 & ~n12495;
  assign n12497 = n12496 ^ n522;
  assign n12498 = n12497 ^ n12447;
  assign n12499 = n12451 & ~n12498;
  assign n12500 = n12499 ^ n12450;
  assign n12502 = n12501 ^ n12500;
  assign n12503 = n12501 ^ n533;
  assign n12504 = n12502 & ~n12503;
  assign n12505 = n12504 ^ n533;
  assign n12506 = n12505 ^ n12445;
  assign n12507 = n12446 & ~n12506;
  assign n12508 = n12507 ^ n781;
  assign n12509 = n12508 ^ n12443;
  assign n12510 = ~n12444 & n12509;
  assign n12511 = n12510 ^ n787;
  assign n12512 = n12511 ^ n12441;
  assign n12513 = ~n12442 & n12512;
  assign n12514 = n12513 ^ n799;
  assign n12516 = n12515 ^ n12514;
  assign n12517 = n12515 ^ n881;
  assign n12518 = ~n12516 & n12517;
  assign n12519 = n12518 ^ n881;
  assign n12520 = n12519 ^ n12439;
  assign n12521 = ~n12440 & n12520;
  assign n12522 = n12521 ^ n896;
  assign n12524 = n12523 ^ n12522;
  assign n12525 = n12523 ^ n1037;
  assign n12526 = ~n12524 & n12525;
  assign n12527 = n12526 ^ n1037;
  assign n12528 = n12527 ^ n12437;
  assign n12529 = ~n12438 & n12528;
  assign n12530 = n12529 ^ n1207;
  assign n12531 = n12530 ^ n12435;
  assign n12532 = ~n12436 & n12531;
  assign n12533 = n12532 ^ n1213;
  assign n12534 = n12533 ^ n12433;
  assign n12535 = n12434 & ~n12534;
  assign n12536 = n12535 ^ n2267;
  assign n12538 = n12537 ^ n12536;
  assign n1533 = x422 ^ x70;
  assign n1534 = n1533 ^ x262;
  assign n1535 = n1534 ^ x6;
  assign n12539 = n12537 ^ n1535;
  assign n12540 = ~n12538 & n12539;
  assign n12541 = n12540 ^ n1535;
  assign n12361 = n12360 ^ n12258;
  assign n12362 = n12259 & ~n12361;
  assign n12363 = n12362 ^ n9430;
  assign n12085 = n12084 ^ n12081;
  assign n12242 = n12241 ^ n12081;
  assign n12243 = n12085 & ~n12242;
  assign n12244 = n12243 ^ n12084;
  assign n12076 = n10607 ^ n9997;
  assign n12077 = ~n11307 & ~n12076;
  assign n12078 = n12077 ^ n9997;
  assign n12254 = n12244 ^ n12078;
  assign n12075 = n11837 ^ n11783;
  assign n12255 = n12254 ^ n12075;
  assign n12256 = n12255 ^ n9446;
  assign n12424 = n12363 ^ n12256;
  assign n12423 = ~n12383 & ~n12422;
  assign n12431 = n12424 ^ n12423;
  assign n12432 = n12431 ^ n2360;
  assign n12605 = n12541 ^ n12432;
  assign n12677 = n12608 ^ n12605;
  assign n12718 = n12677 ^ n10105;
  assign n12754 = n12718 & n12753;
  assign n12755 = n12754 ^ n1572;
  assign n12609 = n12605 & ~n12608;
  assign n12601 = n10802 ^ n10670;
  assign n12602 = ~n12030 & n12601;
  assign n12603 = n12602 ^ n10802;
  assign n12680 = n12609 ^ n12603;
  assign n12542 = n12541 ^ n12431;
  assign n12543 = n12432 & ~n12542;
  assign n12544 = n12543 ^ n2360;
  assign n12425 = ~n12423 & n12424;
  assign n12364 = n12363 ^ n12255;
  assign n12365 = n12256 & n12364;
  assign n12366 = n12365 ^ n9446;
  assign n12248 = n10665 ^ n9975;
  assign n12249 = n11301 & n12248;
  assign n12250 = n12249 ^ n9975;
  assign n12079 = n12078 ^ n12075;
  assign n12245 = n12244 ^ n12075;
  assign n12246 = ~n12079 & n12245;
  assign n12247 = n12246 ^ n12078;
  assign n12251 = n12250 ^ n12247;
  assign n12073 = n11840 ^ x488;
  assign n12074 = n12073 ^ n11780;
  assign n12252 = n12251 ^ n12074;
  assign n12253 = n12252 ^ n9424;
  assign n12382 = n12366 ^ n12253;
  assign n12429 = n12425 ^ n12382;
  assign n12430 = n12429 ^ n2522;
  assign n12600 = n12544 ^ n12430;
  assign n12681 = n12680 ^ n12600;
  assign n12678 = n10105 & ~n12677;
  assign n12679 = n12678 ^ n10132;
  assign n12719 = n12681 ^ n12679;
  assign n12756 = n12719 ^ n12718;
  assign n12757 = n12756 ^ n12754;
  assign n12758 = n12755 & n12757;
  assign n12759 = n12758 ^ n1572;
  assign n12720 = ~n12718 & n12719;
  assign n12682 = n12681 ^ n12678;
  assign n12683 = ~n12679 & n12682;
  assign n12684 = n12683 ^ n10132;
  assign n12545 = n12544 ^ n12429;
  assign n12546 = n12430 & ~n12545;
  assign n12547 = n12546 ^ n2522;
  assign n12426 = ~n12382 & n12425;
  assign n12377 = n11843 ^ n11779;
  assign n12373 = n12250 ^ n12074;
  assign n12374 = n12247 ^ n12074;
  assign n12375 = n12373 & n12374;
  assign n12376 = n12375 ^ n12250;
  assign n12378 = n12377 ^ n12376;
  assign n12370 = n10840 ^ n9969;
  assign n12371 = ~n11295 & n12370;
  assign n12372 = n12371 ^ n9969;
  assign n12379 = n12378 ^ n12372;
  assign n12380 = n12379 ^ n9418;
  assign n12367 = n12366 ^ n12252;
  assign n12368 = n12253 & n12367;
  assign n12369 = n12368 ^ n9424;
  assign n12381 = n12380 ^ n12369;
  assign n12427 = n12426 ^ n12381;
  assign n12428 = n12427 ^ n2538;
  assign n12617 = n12547 ^ n12428;
  assign n12613 = n11345 ^ n10691;
  assign n12614 = n12180 & n12613;
  assign n12615 = n12614 ^ n10691;
  assign n12674 = n12617 ^ n12615;
  assign n12604 = n12603 ^ n12600;
  assign n12610 = n12609 ^ n12600;
  assign n12611 = n12604 & n12610;
  assign n12612 = n12611 ^ n12609;
  assign n12675 = n12674 ^ n12612;
  assign n12676 = n12675 ^ n10227;
  assign n12717 = n12684 ^ n12676;
  assign n12749 = n12720 ^ n12717;
  assign n12750 = n12749 ^ n1578;
  assign n13322 = n12759 ^ n12750;
  assign n12900 = n12478 ^ n2162;
  assign n12897 = n11519 ^ n10734;
  assign n12898 = ~n12115 & ~n12897;
  assign n12899 = n12898 ^ n10734;
  assign n12901 = n12900 ^ n12899;
  assign n12905 = n12473 ^ n12460;
  assign n12902 = n11524 ^ n10735;
  assign n12903 = n12120 & ~n12902;
  assign n12904 = n12903 ^ n10735;
  assign n12906 = n12905 ^ n12904;
  assign n12835 = n12470 ^ n2011;
  assign n12832 = n11527 ^ n10741;
  assign n12833 = n12129 & ~n12832;
  assign n12834 = n12833 ^ n10741;
  assign n12836 = n12835 ^ n12834;
  assign n12812 = n12465 ^ n12462;
  assign n12808 = n11532 ^ n10746;
  assign n12809 = n12134 & ~n12808;
  assign n12810 = n12809 ^ n10746;
  assign n12828 = n12812 ^ n12810;
  assign n12044 = n12017 ^ n11996;
  assign n12041 = n11541 ^ n10757;
  assign n12042 = n12040 & n12041;
  assign n12043 = n12042 ^ n10757;
  assign n12045 = n12044 ^ n12043;
  assign n12050 = n12014 ^ n11998;
  assign n12047 = n11550 ^ n10763;
  assign n12048 = ~n12046 & ~n12047;
  assign n12049 = n12048 ^ n10763;
  assign n12051 = n12050 ^ n12049;
  assign n12057 = n12011 ^ n1595;
  assign n12054 = n11555 ^ n10768;
  assign n12055 = n12053 & n12054;
  assign n12056 = n12055 ^ n10768;
  assign n12058 = n12057 ^ n12056;
  assign n12062 = n11557 ^ n10776;
  assign n12063 = n12061 & ~n12062;
  assign n12064 = n12063 ^ n10776;
  assign n12059 = n12006 ^ n12000;
  assign n12065 = n12064 ^ n12059;
  assign n12630 = n12003 ^ n12002;
  assign n12069 = n11572 ^ n10672;
  assign n12070 = n12068 & n12069;
  assign n12071 = n12070 ^ n10672;
  assign n12066 = n11975 ^ n1470;
  assign n12072 = n12071 ^ n12066;
  assign n12591 = n11488 ^ n10679;
  assign n12592 = ~n12168 & n12591;
  assign n12593 = n12592 ^ n10679;
  assign n12584 = n11849 ^ n11775;
  assign n12581 = n10809 ^ n10046;
  assign n12582 = ~n11292 & n12581;
  assign n12583 = n12582 ^ n10046;
  assign n12585 = n12584 ^ n12583;
  assign n12586 = n12585 ^ n9206;
  assign n12561 = n11846 ^ x486;
  assign n12562 = n12561 ^ n11776;
  assign n12558 = n12377 ^ n12372;
  assign n12559 = n12378 & n12558;
  assign n12560 = n12559 ^ n12372;
  assign n12563 = n12562 ^ n12560;
  assign n12555 = n10817 ^ n10011;
  assign n12556 = n11323 & n12555;
  assign n12557 = n12556 ^ n10011;
  assign n12578 = n12562 ^ n12557;
  assign n12579 = n12563 & n12578;
  assign n12580 = n12579 ^ n12557;
  assign n12587 = n12586 ^ n12580;
  assign n12564 = n12563 ^ n12557;
  assign n12551 = n12379 ^ n12369;
  assign n12552 = n12380 & n12551;
  assign n12553 = n12552 ^ n9418;
  assign n12554 = n12553 ^ n9210;
  assign n12565 = n12564 ^ n12554;
  assign n12566 = ~n12381 & ~n12426;
  assign n12577 = n12565 & ~n12566;
  assign n12588 = n12587 ^ n12577;
  assign n12573 = n12564 ^ n9210;
  assign n12574 = n12564 ^ n12553;
  assign n12575 = ~n12573 & n12574;
  assign n12576 = n12575 ^ n9210;
  assign n12589 = n12588 ^ n12576;
  assign n12567 = n12566 ^ n12565;
  assign n12548 = n12547 ^ n12427;
  assign n12549 = n12428 & ~n12548;
  assign n12550 = n12549 ^ n2538;
  assign n12568 = n12567 ^ n12550;
  assign n12569 = n12567 ^ n2625;
  assign n12570 = ~n12568 & n12569;
  assign n12571 = n12570 ^ n2625;
  assign n12572 = n12571 ^ n1487;
  assign n12590 = n12589 ^ n12572;
  assign n12594 = n12593 ^ n12590;
  assign n12598 = n12568 ^ n2625;
  assign n12595 = n11403 ^ n10686;
  assign n12596 = ~n12174 & n12595;
  assign n12597 = n12596 ^ n10686;
  assign n12599 = n12598 ^ n12597;
  assign n12616 = n12615 ^ n12612;
  assign n12618 = n12617 ^ n12612;
  assign n12619 = ~n12616 & ~n12618;
  assign n12620 = n12619 ^ n12615;
  assign n12621 = n12620 ^ n12598;
  assign n12622 = n12599 & n12621;
  assign n12623 = n12622 ^ n12597;
  assign n12624 = n12623 ^ n12590;
  assign n12625 = ~n12594 & n12624;
  assign n12626 = n12625 ^ n12593;
  assign n12627 = n12626 ^ n12066;
  assign n12628 = ~n12072 & n12627;
  assign n12629 = n12628 ^ n12071;
  assign n12631 = n12630 ^ n12629;
  assign n12632 = n11566 ^ n10140;
  assign n12633 = n12159 & n12632;
  assign n12634 = n12633 ^ n10140;
  assign n12635 = n12634 ^ n12630;
  assign n12636 = ~n12631 & ~n12635;
  assign n12637 = n12636 ^ n12634;
  assign n12638 = n12637 ^ n12059;
  assign n12639 = ~n12065 & ~n12638;
  assign n12640 = n12639 ^ n12064;
  assign n12641 = n12640 ^ n12057;
  assign n12642 = ~n12058 & ~n12641;
  assign n12643 = n12642 ^ n12056;
  assign n12644 = n12643 ^ n12050;
  assign n12645 = ~n12051 & n12644;
  assign n12646 = n12645 ^ n12049;
  assign n12647 = n12646 ^ n12044;
  assign n12648 = n12045 & n12647;
  assign n12649 = n12648 ^ n12043;
  assign n12038 = n12037 ^ n12020;
  assign n12804 = n12649 ^ n12038;
  assign n11498 = n11497 ^ n10752;
  assign n11499 = n11495 & ~n11498;
  assign n11500 = n11499 ^ n10752;
  assign n12805 = n12649 ^ n11500;
  assign n12806 = n12804 & ~n12805;
  assign n12807 = n12806 ^ n12038;
  assign n12829 = n12812 ^ n12807;
  assign n12830 = ~n12828 & ~n12829;
  assign n12831 = n12830 ^ n12810;
  assign n12907 = n12835 ^ n12831;
  assign n12908 = ~n12836 & ~n12907;
  assign n12909 = n12908 ^ n12834;
  assign n12910 = n12909 ^ n12905;
  assign n12911 = n12906 & n12910;
  assign n12912 = n12911 ^ n12904;
  assign n12913 = n12912 ^ n12900;
  assign n12914 = ~n12901 & ~n12913;
  assign n12915 = n12914 ^ n12899;
  assign n12892 = n11513 ^ n10728;
  assign n12893 = n12109 & n12892;
  assign n12894 = n12893 ^ n10728;
  assign n12968 = n12915 ^ n12894;
  assign n12895 = n12481 ^ n12458;
  assign n12969 = n12968 ^ n12895;
  assign n12970 = n12969 ^ n10160;
  assign n12971 = n12912 ^ n12899;
  assign n12972 = n12971 ^ n12900;
  assign n12973 = n12972 ^ n10275;
  assign n12974 = n12909 ^ n12906;
  assign n12975 = n12974 ^ n10165;
  assign n12837 = n12836 ^ n12831;
  assign n12838 = n12837 ^ n10171;
  assign n12811 = n12810 ^ n12807;
  assign n12813 = n12812 ^ n12811;
  assign n12814 = n12813 ^ n10176;
  assign n12652 = n12646 ^ n12043;
  assign n12653 = n12652 ^ n12044;
  assign n12654 = n12653 ^ n10187;
  assign n12655 = n12643 ^ n12049;
  assign n12656 = n12655 ^ n12050;
  assign n12657 = n12656 ^ n10190;
  assign n12658 = n12640 ^ n12056;
  assign n12659 = n12658 ^ n12057;
  assign n12660 = n12659 ^ n10141;
  assign n12661 = n12637 ^ n12064;
  assign n12662 = n12661 ^ n12059;
  assign n12663 = n12662 ^ n10199;
  assign n12664 = n12634 ^ n12631;
  assign n12665 = n12664 ^ n10204;
  assign n12666 = n12626 ^ n12071;
  assign n12667 = n12666 ^ n12066;
  assign n12668 = n12667 ^ n10210;
  assign n12669 = n12623 ^ n12593;
  assign n12670 = n12669 ^ n12590;
  assign n12671 = n12670 ^ n10216;
  assign n12672 = n12620 ^ n12599;
  assign n12673 = n12672 ^ n10222;
  assign n12685 = n12684 ^ n12675;
  assign n12686 = ~n12676 & ~n12685;
  assign n12687 = n12686 ^ n10227;
  assign n12688 = n12687 ^ n12672;
  assign n12689 = n12673 & n12688;
  assign n12690 = n12689 ^ n10222;
  assign n12691 = n12690 ^ n12670;
  assign n12692 = n12671 & ~n12691;
  assign n12693 = n12692 ^ n10216;
  assign n12694 = n12693 ^ n12667;
  assign n12695 = n12668 & ~n12694;
  assign n12696 = n12695 ^ n10210;
  assign n12697 = n12696 ^ n12664;
  assign n12698 = ~n12665 & ~n12697;
  assign n12699 = n12698 ^ n10204;
  assign n12700 = n12699 ^ n12662;
  assign n12701 = ~n12663 & ~n12700;
  assign n12702 = n12701 ^ n10199;
  assign n12703 = n12702 ^ n12659;
  assign n12704 = ~n12660 & ~n12703;
  assign n12705 = n12704 ^ n10141;
  assign n12706 = n12705 ^ n12656;
  assign n12707 = n12657 & ~n12706;
  assign n12708 = n12707 ^ n10190;
  assign n12709 = n12708 ^ n12653;
  assign n12710 = n12654 & n12709;
  assign n12711 = n12710 ^ n10187;
  assign n12800 = n12711 ^ n10182;
  assign n12039 = n12038 ^ n11500;
  assign n12650 = n12649 ^ n12039;
  assign n12801 = n12711 ^ n12650;
  assign n12802 = ~n12800 & n12801;
  assign n12803 = n12802 ^ n10182;
  assign n12825 = n12813 ^ n12803;
  assign n12826 = n12814 & n12825;
  assign n12827 = n12826 ^ n10176;
  assign n12976 = n12837 ^ n12827;
  assign n12977 = ~n12838 & n12976;
  assign n12978 = n12977 ^ n10171;
  assign n12979 = n12978 ^ n12974;
  assign n12980 = ~n12975 & n12979;
  assign n12981 = n12980 ^ n10165;
  assign n12982 = n12981 ^ n12972;
  assign n12983 = n12973 & n12982;
  assign n12984 = n12983 ^ n10275;
  assign n12985 = n12984 ^ n12969;
  assign n12986 = ~n12970 & n12985;
  assign n12987 = n12986 ^ n10160;
  assign n12896 = n12895 ^ n12894;
  assign n12916 = n12915 ^ n12895;
  assign n12917 = ~n12896 & ~n12916;
  assign n12918 = n12917 ^ n12894;
  assign n12887 = n11508 ^ n10723;
  assign n12888 = ~n12104 & n12887;
  assign n12889 = n12888 ^ n10723;
  assign n12965 = n12918 ^ n12889;
  assign n12890 = n12486 ^ n601;
  assign n12966 = n12965 ^ n12890;
  assign n12967 = n12966 ^ n10155;
  assign n13037 = n12987 ^ n12967;
  assign n12651 = n12650 ^ n10182;
  assign n12712 = n12711 ^ n12651;
  assign n12713 = n12705 ^ n12657;
  assign n12714 = n12699 ^ n12663;
  assign n12715 = n12696 ^ n12665;
  assign n12716 = n12693 ^ n12668;
  assign n12721 = n12717 & n12720;
  assign n12722 = n12687 ^ n12673;
  assign n12723 = ~n12721 & ~n12722;
  assign n12724 = n12690 ^ n12671;
  assign n12725 = n12723 & n12724;
  assign n12726 = ~n12716 & ~n12725;
  assign n12727 = n12715 & n12726;
  assign n12728 = n12714 & ~n12727;
  assign n12729 = n12702 ^ n12660;
  assign n12730 = n12728 & ~n12729;
  assign n12731 = n12713 & ~n12730;
  assign n12732 = n12708 ^ n12654;
  assign n12733 = n12731 & n12732;
  assign n12799 = n12712 & ~n12733;
  assign n12815 = n12814 ^ n12803;
  assign n12824 = n12799 & ~n12815;
  assign n12839 = n12838 ^ n12827;
  assign n13030 = n12824 & ~n12839;
  assign n13031 = n12978 ^ n12975;
  assign n13032 = n13030 & ~n13031;
  assign n13033 = n12981 ^ n12973;
  assign n13034 = ~n13032 & ~n13033;
  assign n13035 = n12984 ^ n12970;
  assign n13036 = n13034 & ~n13035;
  assign n13101 = n13037 ^ n13036;
  assign n13096 = n13035 ^ n13034;
  assign n13083 = n13033 ^ n13032;
  assign n13084 = n13083 ^ n638;
  assign n13088 = n13031 ^ n13030;
  assign n12840 = n12839 ^ n12824;
  assign n12844 = n12843 ^ n12840;
  assign n12816 = n12815 ^ n12799;
  assign n12734 = n12733 ^ n12712;
  assign n12738 = n12737 ^ n12734;
  assign n12788 = n12732 ^ n12731;
  assign n12739 = n12730 ^ n12713;
  assign n12740 = n12739 ^ n578;
  assign n12780 = n12729 ^ n12728;
  assign n12741 = n12727 ^ n12714;
  assign n12742 = n12741 ^ n1899;
  assign n12743 = n12726 ^ n12715;
  assign n12744 = n12743 ^ n1748;
  assign n12745 = n12725 ^ n12716;
  assign n12746 = n12745 ^ n1751;
  assign n12747 = n12724 ^ n12723;
  assign n12748 = n12747 ^ n1652;
  assign n12763 = n12722 ^ n12721;
  assign n12760 = n12759 ^ n12749;
  assign n12761 = n12750 & ~n12760;
  assign n12762 = n12761 ^ n1578;
  assign n12764 = n12763 ^ n12762;
  assign n12765 = n12763 ^ n1590;
  assign n12766 = n12764 & ~n12765;
  assign n12767 = n12766 ^ n1590;
  assign n12768 = n12767 ^ n12747;
  assign n12769 = ~n12748 & n12768;
  assign n12770 = n12769 ^ n1652;
  assign n12771 = n12770 ^ n12745;
  assign n12772 = n12746 & ~n12771;
  assign n12773 = n12772 ^ n1751;
  assign n12774 = n12773 ^ n12743;
  assign n12775 = n12744 & ~n12774;
  assign n12776 = n12775 ^ n1748;
  assign n12777 = n12776 ^ n12741;
  assign n12778 = n12742 & ~n12777;
  assign n12779 = n12778 ^ n1899;
  assign n12781 = n12780 ^ n12779;
  assign n12782 = n12780 ^ n2130;
  assign n12783 = ~n12781 & n12782;
  assign n12784 = n12783 ^ n2130;
  assign n12785 = n12784 ^ n12739;
  assign n12786 = ~n12740 & n12785;
  assign n12787 = n12786 ^ n578;
  assign n12789 = n12788 ^ n12787;
  assign n12793 = n12792 ^ n12788;
  assign n12794 = ~n12789 & n12793;
  assign n12795 = n12794 ^ n12792;
  assign n12796 = n12795 ^ n12734;
  assign n12797 = n12738 & ~n12796;
  assign n12798 = n12797 ^ n12737;
  assign n12817 = n12816 ^ n12798;
  assign n12821 = n12820 ^ n12816;
  assign n12822 = ~n12817 & n12821;
  assign n12823 = n12822 ^ n12820;
  assign n13085 = n12840 ^ n12823;
  assign n13086 = n12844 & ~n13085;
  assign n13087 = n13086 ^ n12843;
  assign n13089 = n13088 ^ n13087;
  assign n13090 = n13088 ^ n632;
  assign n13091 = ~n13089 & n13090;
  assign n13092 = n13091 ^ n632;
  assign n13093 = n13092 ^ n13083;
  assign n13094 = n13084 & ~n13093;
  assign n13095 = n13094 ^ n638;
  assign n13097 = n13096 ^ n13095;
  assign n13098 = n13096 ^ n547;
  assign n13099 = n13097 & ~n13098;
  assign n13100 = n13099 ^ n547;
  assign n13102 = n13101 ^ n13100;
  assign n13466 = n13102 ^ n553;
  assign n13065 = n12524 ^ n1037;
  assign n13463 = n12377 ^ n11870;
  assign n13464 = n13065 & n13463;
  assign n13465 = n13464 ^ n11870;
  assign n13467 = n13466 ^ n13465;
  assign n13471 = n13097 ^ n547;
  assign n13023 = n12519 ^ n12440;
  assign n13468 = n12074 ^ n11765;
  assign n13469 = ~n13023 & n13468;
  assign n13470 = n13469 ^ n11765;
  assign n13472 = n13471 ^ n13470;
  assign n13476 = n13092 ^ n13084;
  assign n12947 = n12516 ^ n881;
  assign n13473 = n12075 ^ n11749;
  assign n13474 = n12947 & n13473;
  assign n13475 = n13474 ^ n11749;
  assign n13477 = n13476 ^ n13475;
  assign n13481 = n13089 ^ n632;
  assign n12856 = n12511 ^ n12442;
  assign n13478 = n12081 ^ n11705;
  assign n13479 = ~n12856 & n13478;
  assign n13480 = n13479 ^ n11705;
  assign n13482 = n13481 ^ n13480;
  assign n12861 = n12508 ^ n12444;
  assign n13483 = n12087 ^ n11619;
  assign n13484 = ~n12861 & ~n13483;
  assign n13485 = n13484 ^ n11619;
  assign n12845 = n12844 ^ n12823;
  assign n13486 = n13485 ^ n12845;
  assign n12866 = n12505 ^ n12446;
  assign n13487 = n12093 ^ n11508;
  assign n13488 = n12866 & ~n13487;
  assign n13489 = n13488 ^ n11508;
  assign n13388 = n12820 ^ n12817;
  assign n13490 = n13489 ^ n13388;
  assign n12871 = n12502 ^ n533;
  assign n13491 = n12098 ^ n11513;
  assign n13492 = ~n12871 & n13491;
  assign n13493 = n13492 ^ n11513;
  assign n13394 = n12795 ^ n12738;
  assign n13494 = n13493 ^ n13394;
  assign n12846 = n12497 ^ n12451;
  assign n13495 = n12104 ^ n11519;
  assign n13496 = n12846 & n13495;
  assign n13497 = n13496 ^ n11519;
  assign n13400 = n12792 ^ n12789;
  assign n13498 = n13497 ^ n13400;
  assign n12877 = n12494 ^ n522;
  assign n13499 = n12109 ^ n11524;
  assign n13500 = ~n12877 & n13499;
  assign n13501 = n13500 ^ n11524;
  assign n13406 = n12784 ^ n12740;
  assign n13502 = n13501 ^ n13406;
  assign n12882 = n12489 ^ n12453;
  assign n13503 = n12115 ^ n11527;
  assign n13504 = n12882 & n13503;
  assign n13505 = n13504 ^ n11527;
  assign n13412 = n12781 ^ n2130;
  assign n13506 = n13505 ^ n13412;
  assign n13507 = n12120 ^ n11532;
  assign n13508 = ~n12890 & n13507;
  assign n13509 = n13508 ^ n11532;
  assign n13419 = n12776 ^ n12742;
  assign n13510 = n13509 ^ n13419;
  assign n13511 = n12129 ^ n11497;
  assign n13512 = n12895 & ~n13511;
  assign n13513 = n13512 ^ n11497;
  assign n13425 = n12773 ^ n12744;
  assign n13514 = n13513 ^ n13425;
  assign n13515 = n12134 ^ n11541;
  assign n13516 = ~n12900 & n13515;
  assign n13517 = n13516 ^ n11541;
  assign n13431 = n12770 ^ n12746;
  assign n13518 = n13517 ^ n13431;
  assign n13519 = n11550 ^ n11495;
  assign n13520 = ~n12905 & n13519;
  assign n13521 = n13520 ^ n11550;
  assign n13436 = n12767 ^ n12748;
  assign n13522 = n13521 ^ n13436;
  assign n13380 = n12764 ^ n1590;
  assign n13376 = n12040 ^ n11555;
  assign n13377 = ~n12835 & ~n13376;
  assign n13378 = n13377 ^ n11555;
  assign n13523 = n13380 ^ n13378;
  assign n13323 = n12046 ^ n11557;
  assign n13324 = n12812 & n13323;
  assign n13325 = n13324 ^ n11557;
  assign n13326 = n13325 ^ n13322;
  assign n13310 = n12756 ^ n12755;
  assign n13295 = n12753 ^ n12718;
  assign n13291 = n12061 ^ n11572;
  assign n13292 = n12044 & n13291;
  assign n13293 = n13292 ^ n11572;
  assign n13306 = n13295 ^ n13293;
  assign n13277 = n12159 ^ n11488;
  assign n13278 = n12050 & n13277;
  assign n13279 = n13278 ^ n11488;
  assign n13019 = n11301 ^ n10574;
  assign n13020 = ~n12584 & n13019;
  assign n13021 = n13020 ^ n10574;
  assign n12943 = n11307 ^ n10542;
  assign n12944 = n12562 & ~n12943;
  assign n12945 = n12944 ^ n10542;
  assign n13015 = n12947 ^ n12945;
  assign n12853 = n11959 ^ n11286;
  assign n12854 = ~n12377 & ~n12853;
  assign n12855 = n12854 ^ n11286;
  assign n12857 = n12856 ^ n12855;
  assign n12858 = n11912 ^ n11077;
  assign n12859 = n12074 & n12858;
  assign n12860 = n12859 ^ n11077;
  assign n12862 = n12861 ^ n12860;
  assign n12863 = n11870 ^ n10698;
  assign n12864 = n12075 & ~n12863;
  assign n12865 = n12864 ^ n10698;
  assign n12867 = n12866 ^ n12865;
  assign n12868 = n11765 ^ n10700;
  assign n12869 = ~n12081 & n12868;
  assign n12870 = n12869 ^ n10700;
  assign n12872 = n12871 ^ n12870;
  assign n12873 = n11749 ^ n10705;
  assign n12874 = n12087 & ~n12873;
  assign n12875 = n12874 ^ n10705;
  assign n12876 = n12875 ^ n12846;
  assign n12878 = n11705 ^ n10711;
  assign n12879 = ~n12093 & n12878;
  assign n12880 = n12879 ^ n10711;
  assign n12881 = n12880 ^ n12877;
  assign n12883 = n11619 ^ n10717;
  assign n12884 = ~n12098 & ~n12883;
  assign n12885 = n12884 ^ n10717;
  assign n12886 = n12885 ^ n12882;
  assign n12891 = n12890 ^ n12889;
  assign n12919 = n12918 ^ n12890;
  assign n12920 = ~n12891 & ~n12919;
  assign n12921 = n12920 ^ n12889;
  assign n12922 = n12921 ^ n12882;
  assign n12923 = n12886 & ~n12922;
  assign n12924 = n12923 ^ n12885;
  assign n12925 = n12924 ^ n12877;
  assign n12926 = n12881 & n12925;
  assign n12927 = n12926 ^ n12880;
  assign n12928 = n12927 ^ n12846;
  assign n12929 = ~n12876 & n12928;
  assign n12930 = n12929 ^ n12875;
  assign n12931 = n12930 ^ n12871;
  assign n12932 = ~n12872 & ~n12931;
  assign n12933 = n12932 ^ n12870;
  assign n12934 = n12933 ^ n12866;
  assign n12935 = n12867 & ~n12934;
  assign n12936 = n12935 ^ n12865;
  assign n12937 = n12936 ^ n12861;
  assign n12938 = ~n12862 & n12937;
  assign n12939 = n12938 ^ n12860;
  assign n12940 = n12939 ^ n12856;
  assign n12941 = n12857 & n12940;
  assign n12942 = n12941 ^ n12855;
  assign n13016 = n12947 ^ n12942;
  assign n13017 = n13015 & n13016;
  assign n13018 = n13017 ^ n12945;
  assign n13022 = n13021 ^ n13018;
  assign n13024 = n13023 ^ n13022;
  assign n13025 = n13024 ^ n9981;
  assign n12946 = n12945 ^ n12942;
  assign n12948 = n12947 ^ n12946;
  assign n12949 = n12948 ^ n9987;
  assign n12950 = n12939 ^ n12857;
  assign n12951 = n12950 ^ n10712;
  assign n12952 = n12936 ^ n12862;
  assign n12953 = n12952 ^ n10656;
  assign n12954 = n12933 ^ n12867;
  assign n12955 = n12954 ^ n10602;
  assign n12956 = n12930 ^ n12872;
  assign n12957 = n12956 ^ n10569;
  assign n12958 = n12927 ^ n12875;
  assign n12959 = n12958 ^ n12846;
  assign n12960 = n12959 ^ n10537;
  assign n12961 = n12924 ^ n12881;
  assign n12962 = n12961 ^ n10389;
  assign n12963 = n12921 ^ n12886;
  assign n12964 = n12963 ^ n10289;
  assign n12988 = n12987 ^ n12966;
  assign n12989 = ~n12967 & ~n12988;
  assign n12990 = n12989 ^ n10155;
  assign n12991 = n12990 ^ n12963;
  assign n12992 = n12964 & n12991;
  assign n12993 = n12992 ^ n10289;
  assign n12994 = n12993 ^ n12961;
  assign n12995 = ~n12962 & ~n12994;
  assign n12996 = n12995 ^ n10389;
  assign n12997 = n12996 ^ n12959;
  assign n12998 = ~n12960 & n12997;
  assign n12999 = n12998 ^ n10537;
  assign n13000 = n12999 ^ n12956;
  assign n13001 = n12957 & n13000;
  assign n13002 = n13001 ^ n10569;
  assign n13003 = n13002 ^ n12954;
  assign n13004 = ~n12955 & ~n13003;
  assign n13005 = n13004 ^ n10602;
  assign n13006 = n13005 ^ n12952;
  assign n13007 = ~n12953 & ~n13006;
  assign n13008 = n13007 ^ n10656;
  assign n13009 = n13008 ^ n12950;
  assign n13010 = n12951 & ~n13009;
  assign n13011 = n13010 ^ n10712;
  assign n13012 = n13011 ^ n12948;
  assign n13013 = n12949 & n13012;
  assign n13014 = n13013 ^ n9987;
  assign n13026 = n13025 ^ n13014;
  assign n13027 = n13011 ^ n12949;
  assign n13028 = n12999 ^ n12957;
  assign n13029 = n12996 ^ n12960;
  assign n13038 = ~n13036 & n13037;
  assign n13039 = n12990 ^ n12964;
  assign n13040 = ~n13038 & ~n13039;
  assign n13041 = n12993 ^ n12962;
  assign n13042 = n13040 & ~n13041;
  assign n13043 = n13029 & n13042;
  assign n13044 = ~n13028 & n13043;
  assign n13045 = n13002 ^ n12955;
  assign n13046 = n13044 & ~n13045;
  assign n13047 = n13005 ^ n10656;
  assign n13048 = n13047 ^ n12952;
  assign n13049 = ~n13046 & ~n13048;
  assign n13050 = n13008 ^ n12951;
  assign n13051 = ~n13049 & n13050;
  assign n13052 = ~n13027 & ~n13051;
  assign n13053 = ~n13026 & ~n13052;
  assign n13061 = n11295 ^ n10607;
  assign n13062 = ~n11887 & ~n13061;
  assign n13063 = n13062 ^ n10607;
  assign n13057 = n13023 ^ n13021;
  assign n13058 = n13023 ^ n13018;
  assign n13059 = ~n13057 & n13058;
  assign n13060 = n13059 ^ n13021;
  assign n13064 = n13063 ^ n13060;
  assign n13066 = n13065 ^ n13064;
  assign n13067 = n13066 ^ n9997;
  assign n13054 = n13024 ^ n13014;
  assign n13055 = n13025 & ~n13054;
  assign n13056 = n13055 ^ n9981;
  assign n13068 = n13067 ^ n13056;
  assign n13142 = ~n13053 & ~n13068;
  assign n13154 = n13066 ^ n13056;
  assign n13155 = ~n13067 & n13154;
  assign n13156 = n13155 ^ n9997;
  assign n13147 = n13065 ^ n13063;
  assign n13148 = n13065 ^ n13060;
  assign n13149 = n13147 & ~n13148;
  assign n13150 = n13149 ^ n13063;
  assign n13144 = n11323 ^ n10665;
  assign n13145 = n11881 & n13144;
  assign n13146 = n13145 ^ n10665;
  assign n13151 = n13150 ^ n13146;
  assign n13143 = n12527 ^ n12438;
  assign n13152 = n13151 ^ n13143;
  assign n13153 = n13152 ^ n9975;
  assign n13157 = n13156 ^ n13153;
  assign n13191 = n13142 & ~n13157;
  assign n13187 = n13156 ^ n13152;
  assign n13188 = ~n13153 & ~n13187;
  assign n13189 = n13188 ^ n9975;
  assign n13180 = n13146 ^ n13143;
  assign n13181 = n13150 ^ n13143;
  assign n13182 = ~n13180 & n13181;
  assign n13183 = n13182 ^ n13146;
  assign n13179 = n12530 ^ n12436;
  assign n13184 = n13183 ^ n13179;
  assign n13176 = n11292 ^ n10840;
  assign n13177 = n11876 & n13176;
  assign n13178 = n13177 ^ n10840;
  assign n13185 = n13184 ^ n13178;
  assign n13186 = n13185 ^ n9969;
  assign n13190 = n13189 ^ n13186;
  assign n13192 = n13191 ^ n13190;
  assign n13193 = n13192 ^ n2559;
  assign n13158 = n13157 ^ n13142;
  assign n13069 = n13068 ^ n13053;
  assign n2412 = x293 ^ x101;
  assign n2413 = n2412 ^ x453;
  assign n2414 = n2413 ^ x37;
  assign n13070 = n13069 ^ n2414;
  assign n13134 = n13052 ^ n13026;
  assign n13071 = n13051 ^ n13027;
  assign n13072 = n13071 ^ n1335;
  assign n13073 = n13050 ^ n13049;
  assign n13074 = n13073 ^ n1323;
  assign n13075 = n13048 ^ n13046;
  assign n13076 = n13075 ^ n1144;
  assign n13120 = n13045 ^ n13044;
  assign n13077 = n13043 ^ n13028;
  assign n13078 = n13077 ^ n1001;
  assign n13112 = n13042 ^ n13029;
  assign n13079 = n13041 ^ n13040;
  assign n13080 = n13079 ^ n986;
  assign n13081 = n13039 ^ n13038;
  assign n13082 = n13081 ^ n711;
  assign n13103 = n13101 ^ n553;
  assign n13104 = ~n13102 & n13103;
  assign n13105 = n13104 ^ n553;
  assign n13106 = n13105 ^ n13081;
  assign n13107 = n13082 & ~n13106;
  assign n13108 = n13107 ^ n711;
  assign n13109 = n13108 ^ n13079;
  assign n13110 = ~n13080 & n13109;
  assign n13111 = n13110 ^ n986;
  assign n13113 = n13112 ^ n13111;
  assign n13114 = n13112 ^ n812;
  assign n13115 = ~n13113 & n13114;
  assign n13116 = n13115 ^ n812;
  assign n13117 = n13116 ^ n13077;
  assign n13118 = ~n13078 & n13117;
  assign n13119 = n13118 ^ n1001;
  assign n13121 = n13120 ^ n13119;
  assign n13122 = n13120 ^ n1019;
  assign n13123 = n13121 & ~n13122;
  assign n13124 = n13123 ^ n1019;
  assign n13125 = n13124 ^ n13075;
  assign n13126 = ~n13076 & n13125;
  assign n13127 = n13126 ^ n1144;
  assign n13128 = n13127 ^ n13073;
  assign n13129 = ~n13074 & n13128;
  assign n13130 = n13129 ^ n1323;
  assign n13131 = n13130 ^ n13071;
  assign n13132 = ~n13072 & n13131;
  assign n13133 = n13132 ^ n1335;
  assign n13135 = n13134 ^ n13133;
  assign n13136 = n13134 ^ n2314;
  assign n13137 = ~n13135 & n13136;
  assign n13138 = n13137 ^ n2314;
  assign n13139 = n13138 ^ n13069;
  assign n13140 = ~n13070 & n13139;
  assign n13141 = n13140 ^ n2414;
  assign n13159 = n13158 ^ n13141;
  assign n13173 = n13158 ^ n1511;
  assign n13174 = ~n13159 & n13173;
  assign n13175 = n13174 ^ n1511;
  assign n13232 = n13192 ^ n13175;
  assign n13233 = n13193 & ~n13232;
  assign n13234 = n13233 ^ n2559;
  assign n13229 = ~n13190 & ~n13191;
  assign n13223 = n13179 ^ n13178;
  assign n13224 = n13184 & n13223;
  assign n13225 = n13224 ^ n13178;
  assign n13222 = n12533 ^ n12434;
  assign n13226 = n13225 ^ n13222;
  assign n13219 = n10817 ^ n10684;
  assign n13220 = ~n11920 & ~n13219;
  assign n13221 = n13220 ^ n10817;
  assign n13227 = n13226 ^ n13221;
  assign n13215 = n13189 ^ n13185;
  assign n13216 = ~n13186 & ~n13215;
  assign n13217 = n13216 ^ n9969;
  assign n13218 = n13217 ^ n10011;
  assign n13228 = n13227 ^ n13218;
  assign n13230 = n13229 ^ n13228;
  assign n13231 = n13230 ^ n1424;
  assign n13235 = n13234 ^ n13231;
  assign n13212 = n12068 ^ n11403;
  assign n13213 = n12057 & n13212;
  assign n13214 = n13213 ^ n11403;
  assign n13236 = n13235 ^ n13214;
  assign n13194 = n13193 ^ n13175;
  assign n13170 = n12168 ^ n11345;
  assign n13171 = ~n12059 & n13170;
  assign n13172 = n13171 ^ n11345;
  assign n13195 = n13194 ^ n13172;
  assign n13160 = n13159 ^ n1511;
  assign n12850 = n12174 ^ n10670;
  assign n12851 = n12630 & n12850;
  assign n12852 = n12851 ^ n10670;
  assign n13161 = n13160 ^ n12852;
  assign n13162 = n13138 ^ n13070;
  assign n13163 = n12180 ^ n10676;
  assign n13164 = ~n12066 & n13163;
  assign n13165 = n13164 ^ n10676;
  assign n13166 = ~n13162 & n13165;
  assign n13167 = n13166 ^ n13160;
  assign n13168 = n13161 & n13167;
  assign n13169 = n13168 ^ n13166;
  assign n13209 = n13194 ^ n13169;
  assign n13210 = ~n13195 & ~n13209;
  assign n13211 = n13210 ^ n13172;
  assign n13274 = n13235 ^ n13211;
  assign n13275 = ~n13236 & ~n13274;
  assign n13276 = n13275 ^ n13214;
  assign n13280 = n13279 ^ n13276;
  assign n13265 = n10809 ^ n10678;
  assign n13266 = ~n11968 & ~n13265;
  assign n13267 = n13266 ^ n10809;
  assign n13264 = n12538 ^ n1535;
  assign n13268 = n13267 ^ n13264;
  assign n13269 = n13268 ^ n10046;
  assign n13261 = n13222 ^ n13221;
  assign n13262 = n13226 & n13261;
  assign n13263 = n13262 ^ n13221;
  assign n13270 = n13269 ^ n13263;
  assign n13260 = ~n13228 & ~n13229;
  assign n13271 = n13270 ^ n13260;
  assign n13256 = n13227 ^ n10011;
  assign n13257 = n13227 ^ n13217;
  assign n13258 = ~n13256 & ~n13257;
  assign n13259 = n13258 ^ n10011;
  assign n13272 = n13271 ^ n13259;
  assign n13249 = n13234 ^ n13230;
  assign n13250 = ~n13231 & n13249;
  assign n13251 = n13250 ^ n1424;
  assign n13255 = n13254 ^ n13251;
  assign n13273 = n13272 ^ n13255;
  assign n13288 = n13276 ^ n13273;
  assign n13289 = n13280 & n13288;
  assign n13290 = n13289 ^ n13279;
  assign n13307 = n13295 ^ n13290;
  assign n13308 = n13306 & ~n13307;
  assign n13309 = n13308 ^ n13293;
  assign n13311 = n13310 ^ n13309;
  assign n13303 = n12053 ^ n11566;
  assign n13304 = n12038 & ~n13303;
  assign n13305 = n13304 ^ n11566;
  assign n13319 = n13310 ^ n13305;
  assign n13320 = n13311 & n13319;
  assign n13321 = n13320 ^ n13305;
  assign n13373 = n13322 ^ n13321;
  assign n13374 = ~n13326 & n13373;
  assign n13375 = n13374 ^ n13325;
  assign n13524 = n13380 ^ n13375;
  assign n13525 = n13523 & ~n13524;
  assign n13526 = n13525 ^ n13378;
  assign n13527 = n13526 ^ n13436;
  assign n13528 = ~n13522 & ~n13527;
  assign n13529 = n13528 ^ n13521;
  assign n13530 = n13529 ^ n13431;
  assign n13531 = n13518 & ~n13530;
  assign n13532 = n13531 ^ n13517;
  assign n13533 = n13532 ^ n13425;
  assign n13534 = ~n13514 & ~n13533;
  assign n13535 = n13534 ^ n13513;
  assign n13536 = n13535 ^ n13419;
  assign n13537 = n13510 & n13536;
  assign n13538 = n13537 ^ n13509;
  assign n13539 = n13538 ^ n13412;
  assign n13540 = ~n13506 & ~n13539;
  assign n13541 = n13540 ^ n13505;
  assign n13542 = n13541 ^ n13406;
  assign n13543 = ~n13502 & ~n13542;
  assign n13544 = n13543 ^ n13501;
  assign n13545 = n13544 ^ n13400;
  assign n13546 = ~n13498 & ~n13545;
  assign n13547 = n13546 ^ n13497;
  assign n13548 = n13547 ^ n13394;
  assign n13549 = ~n13494 & n13548;
  assign n13550 = n13549 ^ n13493;
  assign n13551 = n13550 ^ n13388;
  assign n13552 = n13490 & n13551;
  assign n13553 = n13552 ^ n13489;
  assign n13554 = n13553 ^ n12845;
  assign n13555 = ~n13486 & ~n13554;
  assign n13556 = n13555 ^ n13485;
  assign n13557 = n13556 ^ n13481;
  assign n13558 = ~n13482 & n13557;
  assign n13559 = n13558 ^ n13480;
  assign n13560 = n13559 ^ n13476;
  assign n13561 = n13477 & n13560;
  assign n13562 = n13561 ^ n13475;
  assign n13563 = n13562 ^ n13471;
  assign n13564 = ~n13472 & n13563;
  assign n13565 = n13564 ^ n13470;
  assign n13566 = n13565 ^ n13466;
  assign n13567 = ~n13467 & ~n13566;
  assign n13568 = n13567 ^ n13465;
  assign n13461 = n13105 ^ n13082;
  assign n13458 = n12562 ^ n11912;
  assign n13459 = ~n13143 & n13458;
  assign n13460 = n13459 ^ n11912;
  assign n13462 = n13461 ^ n13460;
  assign n13594 = n13568 ^ n13462;
  assign n13595 = n13594 ^ n11077;
  assign n13596 = n13565 ^ n13467;
  assign n13597 = n13596 ^ n10698;
  assign n13598 = n13562 ^ n13472;
  assign n13599 = n13598 ^ n10700;
  assign n13600 = n13559 ^ n13477;
  assign n13601 = n13600 ^ n10705;
  assign n13602 = n13556 ^ n13482;
  assign n13603 = n13602 ^ n10711;
  assign n13604 = n13553 ^ n13486;
  assign n13605 = n13604 ^ n10717;
  assign n13606 = n13550 ^ n13490;
  assign n13607 = n13606 ^ n10723;
  assign n13608 = n13547 ^ n13494;
  assign n13609 = n13608 ^ n10728;
  assign n13610 = n13544 ^ n13497;
  assign n13611 = n13610 ^ n13400;
  assign n13612 = n13611 ^ n10734;
  assign n13613 = n13541 ^ n13502;
  assign n13614 = n13613 ^ n10735;
  assign n13615 = n13538 ^ n13506;
  assign n13616 = n13615 ^ n10741;
  assign n13617 = n13535 ^ n13510;
  assign n13618 = n13617 ^ n10746;
  assign n13619 = n13532 ^ n13514;
  assign n13620 = n13619 ^ n10752;
  assign n13621 = n13529 ^ n13517;
  assign n13622 = n13621 ^ n13431;
  assign n13623 = n13622 ^ n10757;
  assign n13624 = n13526 ^ n13521;
  assign n13625 = n13624 ^ n13436;
  assign n13626 = n13625 ^ n10763;
  assign n13379 = n13378 ^ n13375;
  assign n13381 = n13380 ^ n13379;
  assign n13382 = n13381 ^ n10768;
  assign n13327 = n13326 ^ n13321;
  assign n13328 = n13327 ^ n10776;
  assign n13312 = n13311 ^ n13305;
  assign n13313 = n13312 ^ n10140;
  assign n13294 = n13293 ^ n13290;
  assign n13296 = n13295 ^ n13294;
  assign n13281 = n13280 ^ n13273;
  assign n13282 = n13281 ^ n10679;
  assign n13237 = n13236 ^ n13211;
  assign n13238 = n13237 ^ n10686;
  assign n13196 = n13195 ^ n13169;
  assign n13197 = n13196 ^ n10691;
  assign n13198 = n13165 ^ n13162;
  assign n13199 = ~n10804 & ~n13198;
  assign n13200 = n13199 ^ n10802;
  assign n13201 = n13166 ^ n12852;
  assign n13202 = n13201 ^ n13160;
  assign n13203 = n13202 ^ n13199;
  assign n13204 = ~n13200 & n13203;
  assign n13205 = n13204 ^ n10802;
  assign n13206 = n13205 ^ n13196;
  assign n13207 = n13197 & ~n13206;
  assign n13208 = n13207 ^ n10691;
  assign n13246 = n13237 ^ n13208;
  assign n13247 = n13238 & n13246;
  assign n13248 = n13247 ^ n10686;
  assign n13285 = n13281 ^ n13248;
  assign n13286 = ~n13282 & n13285;
  assign n13287 = n13286 ^ n10679;
  assign n13297 = n13296 ^ n13287;
  assign n13300 = n13296 ^ n10672;
  assign n13301 = ~n13297 & n13300;
  assign n13302 = n13301 ^ n10672;
  assign n13316 = n13312 ^ n13302;
  assign n13317 = ~n13313 & ~n13316;
  assign n13318 = n13317 ^ n10140;
  assign n13370 = n13327 ^ n13318;
  assign n13371 = n13328 & n13370;
  assign n13372 = n13371 ^ n10776;
  assign n13627 = n13381 ^ n13372;
  assign n13628 = n13382 & n13627;
  assign n13629 = n13628 ^ n10768;
  assign n13630 = n13629 ^ n13625;
  assign n13631 = ~n13626 & n13630;
  assign n13632 = n13631 ^ n10763;
  assign n13633 = n13632 ^ n13622;
  assign n13634 = n13623 & n13633;
  assign n13635 = n13634 ^ n10757;
  assign n13636 = n13635 ^ n13619;
  assign n13637 = ~n13620 & n13636;
  assign n13638 = n13637 ^ n10752;
  assign n13639 = n13638 ^ n13617;
  assign n13640 = n13618 & n13639;
  assign n13641 = n13640 ^ n10746;
  assign n13642 = n13641 ^ n13615;
  assign n13643 = ~n13616 & ~n13642;
  assign n13644 = n13643 ^ n10741;
  assign n13645 = n13644 ^ n13613;
  assign n13646 = ~n13614 & ~n13645;
  assign n13647 = n13646 ^ n10735;
  assign n13648 = n13647 ^ n13611;
  assign n13649 = ~n13612 & ~n13648;
  assign n13650 = n13649 ^ n10734;
  assign n13651 = n13650 ^ n13608;
  assign n13652 = ~n13609 & ~n13651;
  assign n13653 = n13652 ^ n10728;
  assign n13654 = n13653 ^ n13606;
  assign n13655 = ~n13607 & ~n13654;
  assign n13656 = n13655 ^ n10723;
  assign n13657 = n13656 ^ n13604;
  assign n13658 = ~n13605 & n13657;
  assign n13659 = n13658 ^ n10717;
  assign n13660 = n13659 ^ n13602;
  assign n13661 = ~n13603 & ~n13660;
  assign n13662 = n13661 ^ n10711;
  assign n13663 = n13662 ^ n13600;
  assign n13664 = n13601 & ~n13663;
  assign n13665 = n13664 ^ n10705;
  assign n13666 = n13665 ^ n13598;
  assign n13667 = ~n13599 & ~n13666;
  assign n13668 = n13667 ^ n10700;
  assign n13669 = n13668 ^ n13596;
  assign n13670 = ~n13597 & n13669;
  assign n13671 = n13670 ^ n10698;
  assign n13672 = n13671 ^ n13594;
  assign n13673 = ~n13595 & n13672;
  assign n13674 = n13673 ^ n11077;
  assign n13569 = n13568 ^ n13461;
  assign n13570 = n13462 & n13569;
  assign n13571 = n13570 ^ n13460;
  assign n13456 = n13108 ^ n13080;
  assign n13453 = n12584 ^ n11959;
  assign n13454 = ~n13179 & ~n13453;
  assign n13455 = n13454 ^ n11959;
  assign n13457 = n13456 ^ n13455;
  assign n13592 = n13571 ^ n13457;
  assign n13593 = n13592 ^ n11286;
  assign n13701 = n13674 ^ n13593;
  assign n13702 = n13659 ^ n13603;
  assign n13703 = n13656 ^ n13605;
  assign n13704 = n13638 ^ n13618;
  assign n13705 = n13632 ^ n13623;
  assign n13239 = n13238 ^ n13208;
  assign n13240 = n13205 ^ n13197;
  assign n13241 = n13198 ^ n10804;
  assign n13242 = n13202 ^ n13200;
  assign n13243 = n13241 & n13242;
  assign n13244 = ~n13240 & n13243;
  assign n13245 = n13239 & ~n13244;
  assign n13283 = n13282 ^ n13248;
  assign n13284 = n13245 & n13283;
  assign n13298 = n13297 ^ n10672;
  assign n13299 = ~n13284 & n13298;
  assign n13314 = n13313 ^ n13302;
  assign n13315 = n13299 & ~n13314;
  assign n13329 = n13328 ^ n13318;
  assign n13369 = ~n13315 & n13329;
  assign n13383 = n13382 ^ n13372;
  assign n13706 = n13369 & ~n13383;
  assign n13707 = n13629 ^ n13626;
  assign n13708 = ~n13706 & n13707;
  assign n13709 = ~n13705 & n13708;
  assign n13710 = n13635 ^ n13620;
  assign n13711 = ~n13709 & n13710;
  assign n13712 = ~n13704 & n13711;
  assign n13713 = n13641 ^ n13616;
  assign n13714 = n13712 & ~n13713;
  assign n13715 = n13644 ^ n13614;
  assign n13716 = n13714 & n13715;
  assign n13717 = n13647 ^ n13612;
  assign n13718 = ~n13716 & n13717;
  assign n13719 = n13650 ^ n13609;
  assign n13720 = n13718 & ~n13719;
  assign n13721 = n13653 ^ n13607;
  assign n13722 = ~n13720 & ~n13721;
  assign n13723 = ~n13703 & ~n13722;
  assign n13724 = ~n13702 & n13723;
  assign n13725 = n13662 ^ n13601;
  assign n13726 = n13724 & ~n13725;
  assign n13727 = n13665 ^ n13599;
  assign n13728 = n13726 & n13727;
  assign n13729 = n13668 ^ n13597;
  assign n13730 = n13728 & ~n13729;
  assign n13731 = n13671 ^ n13595;
  assign n13732 = ~n13730 & n13731;
  assign n13733 = n13701 & ~n13732;
  assign n13675 = n13674 ^ n13592;
  assign n13676 = n13593 & n13675;
  assign n13677 = n13676 ^ n11286;
  assign n13572 = n13571 ^ n13456;
  assign n13573 = ~n13457 & n13572;
  assign n13574 = n13573 ^ n13455;
  assign n13451 = n13113 ^ n812;
  assign n13448 = n11887 ^ n11307;
  assign n13449 = n13222 & n13448;
  assign n13450 = n13449 ^ n11307;
  assign n13452 = n13451 ^ n13450;
  assign n13590 = n13574 ^ n13452;
  assign n13591 = n13590 ^ n10542;
  assign n13734 = n13677 ^ n13591;
  assign n13735 = ~n13733 & ~n13734;
  assign n13678 = n13677 ^ n13590;
  assign n13679 = ~n13591 & ~n13678;
  assign n13680 = n13679 ^ n10542;
  assign n13575 = n13574 ^ n13451;
  assign n13576 = ~n13452 & ~n13575;
  assign n13577 = n13576 ^ n13450;
  assign n13446 = n13116 ^ n13078;
  assign n13443 = n11881 ^ n11301;
  assign n13444 = n13264 & n13443;
  assign n13445 = n13444 ^ n11301;
  assign n13447 = n13446 ^ n13445;
  assign n13588 = n13577 ^ n13447;
  assign n13589 = n13588 ^ n10574;
  assign n13700 = n13680 ^ n13589;
  assign n13855 = n13735 ^ n13700;
  assign n13758 = n13734 ^ n13733;
  assign n2374 = x487 ^ x135;
  assign n2375 = n2374 ^ x327;
  assign n2376 = n2375 ^ x71;
  assign n13759 = n13758 ^ n2376;
  assign n13760 = n13732 ^ n13701;
  assign n1200 = x328 ^ x136;
  assign n1201 = n1200 ^ x488;
  assign n1202 = n1201 ^ x72;
  assign n13761 = n13760 ^ n1202;
  assign n13762 = n13731 ^ n13730;
  assign n13763 = n13762 ^ n1272;
  assign n13841 = n13729 ^ n13728;
  assign n13764 = n13727 ^ n13726;
  assign n13765 = n13764 ^ n891;
  assign n13833 = n13725 ^ n13724;
  assign n13766 = n13723 ^ n13702;
  assign n13767 = n13766 ^ n767;
  assign n13768 = n13722 ^ n13703;
  assign n13769 = n13768 ^ n705;
  assign n13822 = n13721 ^ n13720;
  assign n13817 = n13719 ^ n13718;
  assign n13770 = n13717 ^ n13716;
  assign n13774 = n13773 ^ n13770;
  assign n13806 = n13715 ^ n13714;
  assign n13775 = n13713 ^ n13712;
  assign n13776 = n13775 ^ n515;
  assign n13795 = n13711 ^ n13704;
  assign n13777 = n13710 ^ n13709;
  assign n13778 = n13777 ^ n588;
  assign n13787 = n13708 ^ n13705;
  assign n13779 = n13707 ^ n13706;
  assign n13780 = n13779 ^ n2178;
  assign n13384 = n13383 ^ n13369;
  assign n13330 = n13329 ^ n13315;
  assign n13331 = n13330 ^ n1843;
  assign n13332 = n13314 ^ n13299;
  assign n13333 = n13332 ^ n1833;
  assign n13334 = n13298 ^ n13284;
  assign n13335 = n13334 ^ n1735;
  assign n13336 = n13283 ^ n13245;
  assign n13337 = n13336 ^ n1723;
  assign n13352 = n13244 ^ n13239;
  assign n13338 = n13243 ^ n13240;
  assign n13339 = n13338 ^ n1439;
  assign n13340 = n1412 & ~n13241;
  assign n13344 = n13343 ^ n13340;
  assign n13345 = n13242 ^ n13241;
  assign n13346 = n13345 ^ n13340;
  assign n13347 = n13344 & ~n13346;
  assign n13348 = n13347 ^ n13343;
  assign n13349 = n13348 ^ n13338;
  assign n13350 = ~n13339 & n13349;
  assign n13351 = n13350 ^ n1439;
  assign n13353 = n13352 ^ n13351;
  assign n13354 = n13352 ^ n1717;
  assign n13355 = ~n13353 & n13354;
  assign n13356 = n13355 ^ n1717;
  assign n13357 = n13356 ^ n13336;
  assign n13358 = ~n13337 & n13357;
  assign n13359 = n13358 ^ n1723;
  assign n13360 = n13359 ^ n13334;
  assign n13361 = ~n13335 & n13360;
  assign n13362 = n13361 ^ n1735;
  assign n13363 = n13362 ^ n13332;
  assign n13364 = ~n13333 & n13363;
  assign n13365 = n13364 ^ n1833;
  assign n13366 = n13365 ^ n13330;
  assign n13367 = n13331 & ~n13366;
  assign n13368 = n13367 ^ n1843;
  assign n13385 = n13384 ^ n13368;
  assign n13781 = n13384 ^ n1980;
  assign n13782 = ~n13385 & n13781;
  assign n13783 = n13782 ^ n1980;
  assign n13784 = n13783 ^ n13779;
  assign n13785 = ~n13780 & n13784;
  assign n13786 = n13785 ^ n2178;
  assign n13788 = n13787 ^ n13786;
  assign n13789 = n13787 ^ n2165;
  assign n13790 = n13788 & ~n13789;
  assign n13791 = n13790 ^ n2165;
  assign n13792 = n13791 ^ n13777;
  assign n13793 = n13778 & ~n13792;
  assign n13794 = n13793 ^ n588;
  assign n13796 = n13795 ^ n13794;
  assign n13800 = n13799 ^ n13795;
  assign n13801 = ~n13796 & n13800;
  assign n13802 = n13801 ^ n13799;
  assign n13803 = n13802 ^ n13775;
  assign n13804 = n13776 & ~n13803;
  assign n13805 = n13804 ^ n515;
  assign n13807 = n13806 ^ n13805;
  assign n13811 = n13810 ^ n13806;
  assign n13812 = n13807 & ~n13811;
  assign n13813 = n13812 ^ n13810;
  assign n13814 = n13813 ^ n13770;
  assign n13815 = ~n13774 & n13814;
  assign n13816 = n13815 ^ n13773;
  assign n13818 = n13817 ^ n13816;
  assign n13819 = n13817 ^ n687;
  assign n13820 = n13818 & ~n13819;
  assign n13821 = n13820 ^ n687;
  assign n13823 = n13822 ^ n13821;
  assign n13824 = n13822 ^ n693;
  assign n13825 = n13823 & ~n13824;
  assign n13826 = n13825 ^ n693;
  assign n13827 = n13826 ^ n13768;
  assign n13828 = n13769 & ~n13827;
  assign n13829 = n13828 ^ n705;
  assign n13830 = n13829 ^ n13766;
  assign n13831 = ~n13767 & n13830;
  assign n13832 = n13831 ^ n767;
  assign n13834 = n13833 ^ n13832;
  assign n13835 = n13833 ^ n873;
  assign n13836 = n13834 & ~n13835;
  assign n13837 = n13836 ^ n873;
  assign n13838 = n13837 ^ n13764;
  assign n13839 = n13765 & ~n13838;
  assign n13840 = n13839 ^ n891;
  assign n13842 = n13841 ^ n13840;
  assign n13843 = n13841 ^ n1026;
  assign n13844 = n13842 & ~n13843;
  assign n13845 = n13844 ^ n1026;
  assign n13846 = n13845 ^ n13762;
  assign n13847 = n13763 & ~n13846;
  assign n13848 = n13847 ^ n1272;
  assign n13849 = n13848 ^ n13760;
  assign n13850 = ~n13761 & n13849;
  assign n13851 = n13850 ^ n1202;
  assign n13852 = n13851 ^ n13758;
  assign n13853 = ~n13759 & n13852;
  assign n13854 = n13853 ^ n2376;
  assign n13856 = n13855 ^ n13854;
  assign n13857 = n13855 ^ n2383;
  assign n13858 = n13856 & ~n13857;
  assign n13859 = n13858 ^ n2383;
  assign n13736 = n13700 & ~n13735;
  assign n13681 = n13680 ^ n13588;
  assign n13682 = n13589 & ~n13681;
  assign n13683 = n13682 ^ n10574;
  assign n13585 = n13121 ^ n1019;
  assign n13581 = n11876 ^ n11295;
  assign n13582 = n12605 & ~n13581;
  assign n13583 = n13582 ^ n11295;
  assign n13578 = n13577 ^ n13446;
  assign n13579 = ~n13447 & ~n13578;
  assign n13580 = n13579 ^ n13445;
  assign n13584 = n13583 ^ n13580;
  assign n13586 = n13585 ^ n13584;
  assign n13587 = n13586 ^ n10607;
  assign n13699 = n13683 ^ n13587;
  assign n13756 = n13736 ^ n13699;
  assign n13757 = n13756 ^ n2395;
  assign n13903 = n13859 ^ n13757;
  assign n13900 = n12180 ^ n12059;
  assign n13901 = n13295 & ~n13900;
  assign n13902 = n13901 ^ n12180;
  assign n14001 = n13903 ^ n13902;
  assign n14064 = n14001 ^ n10676;
  assign n14109 = n1490 & n14064;
  assign n14110 = n14109 ^ n1476;
  assign n13904 = n13902 & ~n13903;
  assign n13895 = n12174 ^ n12057;
  assign n13896 = ~n13310 & ~n13895;
  assign n13897 = n13896 ^ n12174;
  assign n14004 = n13904 ^ n13897;
  assign n13737 = ~n13699 & ~n13736;
  assign n13695 = n13124 ^ n13076;
  assign n13691 = n11920 ^ n11323;
  assign n13692 = n12600 & ~n13691;
  assign n13693 = n13692 ^ n11323;
  assign n13687 = n13585 ^ n13583;
  assign n13688 = n13585 ^ n13580;
  assign n13689 = n13687 & n13688;
  assign n13690 = n13689 ^ n13583;
  assign n13694 = n13693 ^ n13690;
  assign n13696 = n13695 ^ n13694;
  assign n13697 = n13696 ^ n10665;
  assign n13684 = n13683 ^ n13586;
  assign n13685 = n13587 & ~n13684;
  assign n13686 = n13685 ^ n10607;
  assign n13698 = n13697 ^ n13686;
  assign n13863 = n13737 ^ n13698;
  assign n13860 = n13859 ^ n13756;
  assign n13861 = ~n13757 & n13860;
  assign n13862 = n13861 ^ n2395;
  assign n13864 = n13863 ^ n13862;
  assign n13898 = n13864 ^ n2476;
  assign n14005 = n14004 ^ n13898;
  assign n14002 = n10676 & ~n14001;
  assign n14003 = n14002 ^ n10670;
  assign n14065 = n14005 ^ n14003;
  assign n14111 = n14065 ^ n14064;
  assign n14112 = n14111 ^ n14109;
  assign n14113 = n14110 & n14112;
  assign n14114 = n14113 ^ n1476;
  assign n14006 = n14005 ^ n14002;
  assign n14007 = ~n14003 & n14006;
  assign n14008 = n14007 ^ n10670;
  assign n13899 = n13898 ^ n13897;
  assign n13905 = n13904 ^ n13898;
  assign n13906 = n13899 & n13905;
  assign n13907 = n13906 ^ n13904;
  assign n13865 = n13863 ^ n2476;
  assign n13866 = ~n13864 & n13865;
  assign n13867 = n13866 ^ n2476;
  assign n13749 = n13127 ^ n13074;
  assign n13745 = n13695 ^ n13693;
  assign n13746 = n13695 ^ n13690;
  assign n13747 = ~n13745 & ~n13746;
  assign n13748 = n13747 ^ n13693;
  assign n13750 = n13749 ^ n13748;
  assign n13742 = n11968 ^ n11292;
  assign n13743 = n12617 & n13742;
  assign n13744 = n13743 ^ n11292;
  assign n13751 = n13750 ^ n13744;
  assign n13752 = n13751 ^ n10840;
  assign n13739 = n13696 ^ n13686;
  assign n13740 = n13697 & ~n13739;
  assign n13741 = n13740 ^ n10665;
  assign n13753 = n13752 ^ n13741;
  assign n13738 = ~n13698 & n13737;
  assign n13754 = n13753 ^ n13738;
  assign n13755 = n13754 ^ n2471;
  assign n13893 = n13867 ^ n13755;
  assign n13890 = n12168 ^ n12050;
  assign n13891 = n13322 & ~n13890;
  assign n13892 = n13891 ^ n12168;
  assign n13894 = n13893 ^ n13892;
  assign n13999 = n13907 ^ n13894;
  assign n14000 = n13999 ^ n11345;
  assign n14067 = n14008 ^ n14000;
  assign n14066 = ~n14064 & n14065;
  assign n14107 = n14067 ^ n14066;
  assign n14108 = n14107 ^ n1453;
  assign n14556 = n14114 ^ n14108;
  assign n13418 = n13348 ^ n13339;
  assign n15708 = n14556 ^ n13418;
  assign n14401 = n13837 ^ n13765;
  assign n13930 = n13135 ^ n2314;
  assign n14397 = n12600 ^ n11881;
  assign n14398 = n13930 & n14397;
  assign n14399 = n14398 ^ n11881;
  assign n14334 = n13834 ^ n873;
  assign n13881 = n13130 ^ n13072;
  assign n14330 = n12605 ^ n11887;
  assign n14331 = ~n13881 & ~n14330;
  assign n14332 = n14331 ^ n11887;
  assign n14393 = n14334 ^ n14332;
  assign n14289 = n13264 ^ n12584;
  assign n14290 = ~n13749 & ~n14289;
  assign n14291 = n14290 ^ n12584;
  assign n14288 = n13829 ^ n13767;
  assign n14292 = n14291 ^ n14288;
  assign n14247 = n13143 ^ n12074;
  assign n14248 = ~n13446 & ~n14247;
  assign n14249 = n14248 ^ n12074;
  assign n14246 = n13818 ^ n687;
  assign n14250 = n14249 ^ n14246;
  assign n14254 = n13813 ^ n13774;
  assign n14251 = n13065 ^ n12075;
  assign n14252 = n13451 & n14251;
  assign n14253 = n14252 ^ n12075;
  assign n14255 = n14254 ^ n14253;
  assign n14257 = n13023 ^ n12081;
  assign n14258 = ~n13456 & n14257;
  assign n14259 = n14258 ^ n12081;
  assign n14256 = n13810 ^ n13807;
  assign n14260 = n14259 ^ n14256;
  assign n14227 = n13802 ^ n13776;
  assign n14223 = n12947 ^ n12087;
  assign n14224 = n13461 & n14223;
  assign n14225 = n14224 ^ n12087;
  assign n14261 = n14227 ^ n14225;
  assign n14203 = n12856 ^ n12093;
  assign n14204 = n13466 & n14203;
  assign n14205 = n14204 ^ n12093;
  assign n14202 = n13799 ^ n13796;
  assign n14206 = n14205 ^ n14202;
  assign n14183 = n13791 ^ n13778;
  assign n14180 = n12861 ^ n12098;
  assign n14181 = ~n13471 & n14180;
  assign n14182 = n14181 ^ n12098;
  assign n14184 = n14183 ^ n14182;
  assign n14052 = n12866 ^ n12104;
  assign n14053 = n13476 & ~n14052;
  assign n14054 = n14053 ^ n12104;
  assign n14051 = n13788 ^ n2165;
  assign n14055 = n14054 ^ n14051;
  assign n13968 = n12871 ^ n12109;
  assign n13969 = n13481 & ~n13968;
  assign n13970 = n13969 ^ n12109;
  assign n13967 = n13783 ^ n13780;
  assign n13971 = n13970 ^ n13967;
  assign n13386 = n13385 ^ n1980;
  assign n12847 = n12846 ^ n12115;
  assign n12848 = n12845 & ~n12847;
  assign n12849 = n12848 ^ n12115;
  assign n13387 = n13386 ^ n12849;
  assign n13392 = n13365 ^ n13331;
  assign n13389 = n12877 ^ n12120;
  assign n13390 = n13388 & ~n13389;
  assign n13391 = n13390 ^ n12120;
  assign n13393 = n13392 ^ n13391;
  assign n13398 = n13362 ^ n13333;
  assign n13395 = n12882 ^ n12129;
  assign n13396 = n13394 & n13395;
  assign n13397 = n13396 ^ n12129;
  assign n13399 = n13398 ^ n13397;
  assign n13404 = n13359 ^ n13335;
  assign n13401 = n12890 ^ n12134;
  assign n13402 = n13400 & ~n13401;
  assign n13403 = n13402 ^ n12134;
  assign n13405 = n13404 ^ n13403;
  assign n13410 = n13356 ^ n13337;
  assign n13407 = n12895 ^ n11495;
  assign n13408 = ~n13406 & n13407;
  assign n13409 = n13408 ^ n11495;
  assign n13411 = n13410 ^ n13409;
  assign n13416 = n13353 ^ n1717;
  assign n13413 = n12900 ^ n12040;
  assign n13414 = n13412 & ~n13413;
  assign n13415 = n13414 ^ n12040;
  assign n13417 = n13416 ^ n13415;
  assign n13420 = n12905 ^ n12046;
  assign n13421 = n13419 & n13420;
  assign n13422 = n13421 ^ n12046;
  assign n13423 = n13422 ^ n13418;
  assign n13426 = n12835 ^ n12053;
  assign n13427 = n13425 & ~n13426;
  assign n13428 = n13427 ^ n12053;
  assign n13424 = n13345 ^ n13344;
  assign n13429 = n13428 ^ n13424;
  assign n13432 = n12812 ^ n12061;
  assign n13433 = n13431 & n13432;
  assign n13434 = n13433 ^ n12061;
  assign n13430 = n13241 ^ n1412;
  assign n13435 = n13434 ^ n13430;
  assign n13885 = ~n13738 & ~n13753;
  assign n13878 = n13749 ^ n13744;
  assign n13879 = n13750 & n13878;
  assign n13880 = n13879 ^ n13744;
  assign n13882 = n13881 ^ n13880;
  assign n13875 = n11990 ^ n10684;
  assign n13876 = n12598 & ~n13875;
  assign n13877 = n13876 ^ n10684;
  assign n13883 = n13882 ^ n13877;
  assign n13871 = n13751 ^ n13741;
  assign n13872 = ~n13752 & ~n13871;
  assign n13873 = n13872 ^ n10840;
  assign n13874 = n13873 ^ n10817;
  assign n13884 = n13883 ^ n13874;
  assign n13886 = n13885 ^ n13884;
  assign n13868 = n13867 ^ n13754;
  assign n13869 = n13755 & ~n13868;
  assign n13870 = n13869 ^ n2471;
  assign n13887 = n13886 ^ n13870;
  assign n13888 = n13887 ^ n1497;
  assign n13440 = n12068 ^ n12044;
  assign n13441 = ~n13380 & n13440;
  assign n13442 = n13441 ^ n12068;
  assign n13889 = n13888 ^ n13442;
  assign n13908 = n13907 ^ n13893;
  assign n13909 = ~n13894 & ~n13908;
  assign n13910 = n13909 ^ n13892;
  assign n13911 = n13910 ^ n13888;
  assign n13912 = ~n13889 & ~n13911;
  assign n13913 = n13912 ^ n13442;
  assign n13437 = n12159 ^ n12038;
  assign n13438 = ~n13436 & n13437;
  assign n13439 = n13438 ^ n12159;
  assign n13914 = n13913 ^ n13439;
  assign n13927 = n12030 ^ n10678;
  assign n13928 = ~n12590 & ~n13927;
  assign n13929 = n13928 ^ n10678;
  assign n13931 = n13930 ^ n13929;
  assign n13932 = n13931 ^ n10809;
  assign n13924 = n13881 ^ n13877;
  assign n13925 = ~n13882 & n13924;
  assign n13926 = n13925 ^ n13877;
  assign n13933 = n13932 ^ n13926;
  assign n13923 = ~n13884 & ~n13885;
  assign n13934 = n13933 ^ n13923;
  assign n13919 = n13883 ^ n10817;
  assign n13920 = n13883 ^ n13873;
  assign n13921 = ~n13919 & ~n13920;
  assign n13922 = n13921 ^ n10817;
  assign n13935 = n13934 ^ n13922;
  assign n13915 = n13886 ^ n1497;
  assign n13916 = n13887 & ~n13915;
  assign n13917 = n13916 ^ n1497;
  assign n13918 = n13917 ^ n1463;
  assign n13936 = n13935 ^ n13918;
  assign n13937 = n13936 ^ n13913;
  assign n13938 = n13914 & n13937;
  assign n13939 = n13938 ^ n13439;
  assign n13940 = n13939 ^ n13430;
  assign n13941 = ~n13435 & n13940;
  assign n13942 = n13941 ^ n13434;
  assign n13943 = n13942 ^ n13424;
  assign n13944 = n13429 & ~n13943;
  assign n13945 = n13944 ^ n13428;
  assign n13946 = n13945 ^ n13418;
  assign n13947 = n13423 & n13946;
  assign n13948 = n13947 ^ n13422;
  assign n13949 = n13948 ^ n13416;
  assign n13950 = n13417 & n13949;
  assign n13951 = n13950 ^ n13415;
  assign n13952 = n13951 ^ n13410;
  assign n13953 = ~n13411 & n13952;
  assign n13954 = n13953 ^ n13409;
  assign n13955 = n13954 ^ n13404;
  assign n13956 = ~n13405 & n13955;
  assign n13957 = n13956 ^ n13403;
  assign n13958 = n13957 ^ n13398;
  assign n13959 = ~n13399 & n13958;
  assign n13960 = n13959 ^ n13397;
  assign n13961 = n13960 ^ n13392;
  assign n13962 = n13393 & ~n13961;
  assign n13963 = n13962 ^ n13391;
  assign n13964 = n13963 ^ n13386;
  assign n13965 = ~n13387 & ~n13964;
  assign n13966 = n13965 ^ n12849;
  assign n14048 = n13967 ^ n13966;
  assign n14049 = ~n13971 & ~n14048;
  assign n14050 = n14049 ^ n13970;
  assign n14177 = n14051 ^ n14050;
  assign n14178 = n14055 & n14177;
  assign n14179 = n14178 ^ n14054;
  assign n14199 = n14183 ^ n14179;
  assign n14200 = ~n14184 & n14199;
  assign n14201 = n14200 ^ n14182;
  assign n14220 = n14202 ^ n14201;
  assign n14221 = ~n14206 & n14220;
  assign n14222 = n14221 ^ n14205;
  assign n14262 = n14227 ^ n14222;
  assign n14263 = n14261 & n14262;
  assign n14264 = n14263 ^ n14225;
  assign n14265 = n14264 ^ n14256;
  assign n14266 = n14260 & n14265;
  assign n14267 = n14266 ^ n14259;
  assign n14268 = n14267 ^ n14254;
  assign n14269 = ~n14255 & ~n14268;
  assign n14270 = n14269 ^ n14253;
  assign n14271 = n14270 ^ n14246;
  assign n14272 = ~n14250 & n14271;
  assign n14273 = n14272 ^ n14249;
  assign n14245 = n13823 ^ n693;
  assign n14274 = n14273 ^ n14245;
  assign n14275 = n13179 ^ n12377;
  assign n14276 = ~n13585 & n14275;
  assign n14277 = n14276 ^ n12377;
  assign n14278 = n14277 ^ n14245;
  assign n14279 = n14274 & n14278;
  assign n14280 = n14279 ^ n14277;
  assign n14234 = n13826 ^ n13769;
  assign n14281 = n14280 ^ n14234;
  assign n14282 = n13222 ^ n12562;
  assign n14283 = ~n13695 & n14282;
  assign n14284 = n14283 ^ n12562;
  assign n14285 = n14284 ^ n14280;
  assign n14286 = ~n14281 & n14285;
  assign n14287 = n14286 ^ n14234;
  assign n14327 = n14288 ^ n14287;
  assign n14328 = n14292 & n14327;
  assign n14329 = n14328 ^ n14291;
  assign n14394 = n14334 ^ n14329;
  assign n14395 = n14393 & ~n14394;
  assign n14396 = n14395 ^ n14332;
  assign n14400 = n14399 ^ n14396;
  assign n14402 = n14401 ^ n14400;
  assign n14403 = n14402 ^ n11301;
  assign n14333 = n14332 ^ n14329;
  assign n14335 = n14334 ^ n14333;
  assign n14293 = n14292 ^ n14287;
  assign n14294 = n14293 ^ n11959;
  assign n14295 = n14284 ^ n14234;
  assign n14296 = n14295 ^ n14280;
  assign n14297 = n14296 ^ n11912;
  assign n14298 = n14277 ^ n14274;
  assign n14299 = n14298 ^ n11870;
  assign n14300 = n14270 ^ n14250;
  assign n14301 = n14300 ^ n11765;
  assign n14302 = n14267 ^ n14255;
  assign n14303 = n14302 ^ n11749;
  assign n14304 = n14264 ^ n14260;
  assign n14305 = n14304 ^ n11705;
  assign n14226 = n14225 ^ n14222;
  assign n14228 = n14227 ^ n14226;
  assign n14229 = n14228 ^ n11619;
  assign n14207 = n14206 ^ n14201;
  assign n14208 = n14207 ^ n11508;
  assign n14185 = n14184 ^ n14179;
  assign n14186 = n14185 ^ n11513;
  assign n14056 = n14055 ^ n14050;
  assign n14057 = n14056 ^ n11519;
  assign n13972 = n13971 ^ n13966;
  assign n13973 = n13972 ^ n11524;
  assign n13974 = n13963 ^ n12849;
  assign n13975 = n13974 ^ n13386;
  assign n13976 = n13975 ^ n11527;
  assign n13977 = n13960 ^ n13393;
  assign n13978 = n13977 ^ n11532;
  assign n13979 = n13957 ^ n13397;
  assign n13980 = n13979 ^ n13398;
  assign n13981 = n13980 ^ n11497;
  assign n13982 = n13954 ^ n13405;
  assign n13983 = n13982 ^ n11541;
  assign n13984 = n13951 ^ n13411;
  assign n13985 = n13984 ^ n11550;
  assign n13986 = n13948 ^ n13417;
  assign n13987 = n13986 ^ n11555;
  assign n13988 = n13945 ^ n13423;
  assign n13989 = n13988 ^ n11557;
  assign n13990 = n13942 ^ n13429;
  assign n13991 = n13990 ^ n11566;
  assign n13992 = n13939 ^ n13435;
  assign n13993 = n13992 ^ n11572;
  assign n13994 = n13936 ^ n13439;
  assign n13995 = n13994 ^ n13913;
  assign n13996 = n13995 ^ n11488;
  assign n13997 = n13910 ^ n13889;
  assign n13998 = n13997 ^ n11403;
  assign n14009 = n14008 ^ n13999;
  assign n14010 = n14000 & ~n14009;
  assign n14011 = n14010 ^ n11345;
  assign n14012 = n14011 ^ n13997;
  assign n14013 = n13998 & n14012;
  assign n14014 = n14013 ^ n11403;
  assign n14015 = n14014 ^ n13995;
  assign n14016 = ~n13996 & n14015;
  assign n14017 = n14016 ^ n11488;
  assign n14018 = n14017 ^ n13992;
  assign n14019 = ~n13993 & n14018;
  assign n14020 = n14019 ^ n11572;
  assign n14021 = n14020 ^ n13990;
  assign n14022 = ~n13991 & ~n14021;
  assign n14023 = n14022 ^ n11566;
  assign n14024 = n14023 ^ n13988;
  assign n14025 = ~n13989 & n14024;
  assign n14026 = n14025 ^ n11557;
  assign n14027 = n14026 ^ n13986;
  assign n14028 = n13987 & ~n14027;
  assign n14029 = n14028 ^ n11555;
  assign n14030 = n14029 ^ n13984;
  assign n14031 = ~n13985 & ~n14030;
  assign n14032 = n14031 ^ n11550;
  assign n14033 = n14032 ^ n13982;
  assign n14034 = ~n13983 & n14033;
  assign n14035 = n14034 ^ n11541;
  assign n14036 = n14035 ^ n13980;
  assign n14037 = n13981 & n14036;
  assign n14038 = n14037 ^ n11497;
  assign n14039 = n14038 ^ n13977;
  assign n14040 = n13978 & n14039;
  assign n14041 = n14040 ^ n11532;
  assign n14042 = n14041 ^ n13975;
  assign n14043 = n13976 & n14042;
  assign n14044 = n14043 ^ n11527;
  assign n14045 = n14044 ^ n13972;
  assign n14046 = n13973 & n14045;
  assign n14047 = n14046 ^ n11524;
  assign n14174 = n14056 ^ n14047;
  assign n14175 = ~n14057 & ~n14174;
  assign n14176 = n14175 ^ n11519;
  assign n14196 = n14185 ^ n14176;
  assign n14197 = ~n14186 & n14196;
  assign n14198 = n14197 ^ n11513;
  assign n14217 = n14207 ^ n14198;
  assign n14218 = n14208 & n14217;
  assign n14219 = n14218 ^ n11508;
  assign n14306 = n14228 ^ n14219;
  assign n14307 = n14229 & n14306;
  assign n14308 = n14307 ^ n11619;
  assign n14309 = n14308 ^ n14304;
  assign n14310 = ~n14305 & n14309;
  assign n14311 = n14310 ^ n11705;
  assign n14312 = n14311 ^ n14302;
  assign n14313 = n14303 & n14312;
  assign n14314 = n14313 ^ n11749;
  assign n14315 = n14314 ^ n14300;
  assign n14316 = ~n14301 & n14315;
  assign n14317 = n14316 ^ n11765;
  assign n14318 = n14317 ^ n14298;
  assign n14319 = ~n14299 & ~n14318;
  assign n14320 = n14319 ^ n11870;
  assign n14321 = n14320 ^ n14296;
  assign n14322 = ~n14297 & ~n14321;
  assign n14323 = n14322 ^ n11912;
  assign n14324 = n14323 ^ n14293;
  assign n14325 = n14294 & ~n14324;
  assign n14326 = n14325 ^ n11959;
  assign n14336 = n14335 ^ n14326;
  assign n14390 = n14335 ^ n11307;
  assign n14391 = n14336 & n14390;
  assign n14392 = n14391 ^ n11307;
  assign n14404 = n14403 ^ n14392;
  assign n14337 = n14336 ^ n11307;
  assign n14338 = n14314 ^ n14301;
  assign n14339 = n14311 ^ n14303;
  assign n14340 = n14308 ^ n14305;
  assign n14209 = n14208 ^ n14198;
  assign n14058 = n14057 ^ n14047;
  assign n14059 = n14044 ^ n13973;
  assign n14060 = n14041 ^ n13976;
  assign n14061 = n14038 ^ n13978;
  assign n14062 = n14023 ^ n13989;
  assign n14063 = n14011 ^ n13998;
  assign n14068 = n14066 & ~n14067;
  assign n14069 = n14063 & ~n14068;
  assign n14070 = n14014 ^ n13996;
  assign n14071 = n14069 & n14070;
  assign n14072 = n14017 ^ n13993;
  assign n14073 = ~n14071 & ~n14072;
  assign n14074 = n14020 ^ n13991;
  assign n14075 = n14073 & ~n14074;
  assign n14076 = ~n14062 & ~n14075;
  assign n14077 = n14026 ^ n13987;
  assign n14078 = n14076 & n14077;
  assign n14079 = n14029 ^ n13985;
  assign n14080 = ~n14078 & n14079;
  assign n14081 = n14032 ^ n13983;
  assign n14082 = n14080 & ~n14081;
  assign n14083 = n14035 ^ n13981;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = n14061 & n14084;
  assign n14086 = ~n14060 & n14085;
  assign n14087 = n14059 & n14086;
  assign n14173 = ~n14058 & ~n14087;
  assign n14187 = n14186 ^ n14176;
  assign n14210 = n14173 & n14187;
  assign n14216 = n14209 & ~n14210;
  assign n14230 = n14229 ^ n14219;
  assign n14341 = ~n14216 & n14230;
  assign n14342 = n14340 & n14341;
  assign n14343 = ~n14339 & n14342;
  assign n14344 = ~n14338 & n14343;
  assign n14345 = n14317 ^ n11870;
  assign n14346 = n14345 ^ n14298;
  assign n14347 = n14344 & ~n14346;
  assign n14348 = n14320 ^ n14297;
  assign n14349 = ~n14347 & ~n14348;
  assign n14350 = n14323 ^ n14294;
  assign n14351 = ~n14349 & n14350;
  assign n14405 = ~n14337 & ~n14351;
  assign n14426 = n14404 & ~n14405;
  assign n14422 = n13842 ^ n1026;
  assign n14418 = n12617 ^ n11876;
  assign n14419 = ~n13162 & n14418;
  assign n14420 = n14419 ^ n11876;
  assign n14414 = n14401 ^ n14399;
  assign n14415 = n14401 ^ n14396;
  assign n14416 = n14414 & n14415;
  assign n14417 = n14416 ^ n14399;
  assign n14421 = n14420 ^ n14417;
  assign n14423 = n14422 ^ n14421;
  assign n14424 = n14423 ^ n11295;
  assign n14411 = n14402 ^ n14392;
  assign n14412 = ~n14403 & ~n14411;
  assign n14413 = n14412 ^ n11301;
  assign n14425 = n14424 ^ n14413;
  assign n14427 = n14426 ^ n14425;
  assign n14406 = n14405 ^ n14404;
  assign n14352 = n14351 ^ n14337;
  assign n14353 = n14352 ^ n1315;
  assign n14354 = n14350 ^ n14349;
  assign n14355 = n14354 ^ n1309;
  assign n14356 = n14348 ^ n14347;
  assign n14357 = n14356 ^ n1124;
  assign n14376 = n14346 ^ n14344;
  assign n14358 = n14343 ^ n14338;
  assign n14359 = n14358 ^ n963;
  assign n14368 = n14342 ^ n14339;
  assign n14360 = n14341 ^ n14340;
  assign n14361 = n14360 ^ n847;
  assign n14231 = n14230 ^ n14216;
  assign n14232 = n14231 ^ n841;
  assign n14211 = n14210 ^ n14209;
  assign n14188 = n14187 ^ n14173;
  assign n14088 = n14087 ^ n14058;
  assign n14089 = n14088 ^ n528;
  assign n14165 = n14086 ^ n14059;
  assign n14090 = n14085 ^ n14060;
  assign n14091 = n14090 ^ n610;
  assign n14154 = n14084 ^ n14061;
  assign n14092 = n14083 ^ n14082;
  assign n14096 = n14095 ^ n14092;
  assign n14143 = n14081 ^ n14080;
  assign n14097 = n14079 ^ n14078;
  assign n14098 = n14097 ^ n2101;
  assign n14135 = n14077 ^ n14076;
  assign n14099 = n14075 ^ n14062;
  assign n14100 = n14099 ^ n1955;
  assign n14101 = n14074 ^ n14073;
  assign n14102 = n14101 ^ n1757;
  assign n14103 = n14072 ^ n14071;
  assign n14104 = n14103 ^ n1939;
  assign n14105 = n14070 ^ n14069;
  assign n14106 = n14105 ^ n1640;
  assign n14118 = n14068 ^ n14063;
  assign n14115 = n14114 ^ n14107;
  assign n14116 = ~n14108 & n14115;
  assign n14117 = n14116 ^ n1453;
  assign n14119 = n14118 ^ n14117;
  assign n14120 = n14118 ^ n1459;
  assign n14121 = ~n14119 & n14120;
  assign n14122 = n14121 ^ n1459;
  assign n14123 = n14122 ^ n14105;
  assign n14124 = ~n14106 & n14123;
  assign n14125 = n14124 ^ n1640;
  assign n14126 = n14125 ^ n14103;
  assign n14127 = n14104 & ~n14126;
  assign n14128 = n14127 ^ n1939;
  assign n14129 = n14128 ^ n14101;
  assign n14130 = ~n14102 & n14129;
  assign n14131 = n14130 ^ n1757;
  assign n14132 = n14131 ^ n14099;
  assign n14133 = ~n14100 & n14132;
  assign n14134 = n14133 ^ n1955;
  assign n14136 = n14135 ^ n14134;
  assign n14137 = n14135 ^ n1973;
  assign n14138 = n14136 & ~n14137;
  assign n14139 = n14138 ^ n1973;
  assign n14140 = n14139 ^ n14097;
  assign n14141 = ~n14098 & n14140;
  assign n14142 = n14141 ^ n2101;
  assign n14144 = n14143 ^ n14142;
  assign n14148 = n14147 ^ n14143;
  assign n14149 = n14144 & ~n14148;
  assign n14150 = n14149 ^ n14147;
  assign n14151 = n14150 ^ n14092;
  assign n14152 = ~n14096 & n14151;
  assign n14153 = n14152 ^ n14095;
  assign n14155 = n14154 ^ n14153;
  assign n14159 = n14158 ^ n14154;
  assign n14160 = n14155 & ~n14159;
  assign n14161 = n14160 ^ n14158;
  assign n14162 = n14161 ^ n14090;
  assign n14163 = n14091 & ~n14162;
  assign n14164 = n14163 ^ n610;
  assign n14166 = n14165 ^ n14164;
  assign n14167 = n14165 ^ n575;
  assign n14168 = n14166 & ~n14167;
  assign n14169 = n14168 ^ n575;
  assign n14170 = n14169 ^ n14088;
  assign n14171 = n14089 & ~n14170;
  assign n14172 = n14171 ^ n528;
  assign n14189 = n14188 ^ n14172;
  assign n14193 = n14192 ^ n14188;
  assign n14194 = ~n14189 & n14193;
  assign n14195 = n14194 ^ n14192;
  assign n14212 = n14211 ^ n14195;
  assign n14213 = n14211 ^ n542;
  assign n14214 = ~n14212 & n14213;
  assign n14215 = n14214 ^ n542;
  assign n14362 = n14231 ^ n14215;
  assign n14363 = ~n14232 & n14362;
  assign n14364 = n14363 ^ n841;
  assign n14365 = n14364 ^ n14360;
  assign n14366 = n14361 & ~n14365;
  assign n14367 = n14366 ^ n847;
  assign n14369 = n14368 ^ n14367;
  assign n14370 = n14368 ^ n859;
  assign n14371 = n14369 & ~n14370;
  assign n14372 = n14371 ^ n859;
  assign n14373 = n14372 ^ n14358;
  assign n14374 = ~n14359 & n14373;
  assign n14375 = n14374 ^ n963;
  assign n14377 = n14376 ^ n14375;
  assign n14378 = n14376 ^ n975;
  assign n14379 = n14377 & ~n14378;
  assign n14380 = n14379 ^ n975;
  assign n14381 = n14380 ^ n14356;
  assign n14382 = ~n14357 & n14381;
  assign n14383 = n14382 ^ n1124;
  assign n14384 = n14383 ^ n14354;
  assign n14385 = ~n14355 & n14384;
  assign n14386 = n14385 ^ n1309;
  assign n14387 = n14386 ^ n14352;
  assign n14388 = ~n14353 & n14387;
  assign n14389 = n14388 ^ n1315;
  assign n14407 = n14406 ^ n14389;
  assign n2307 = n2267 ^ x166;
  assign n2308 = n2307 ^ x358;
  assign n2309 = n2308 ^ x102;
  assign n14408 = n14406 ^ n2309;
  assign n14409 = n14407 & ~n14408;
  assign n14410 = n14409 ^ n2309;
  assign n14428 = n14427 ^ n14410;
  assign n1536 = n1535 ^ x165;
  assign n1537 = n1536 ^ x357;
  assign n1538 = n1537 ^ x101;
  assign n14429 = n14428 ^ n1538;
  assign n14243 = n13430 ^ n12059;
  assign n14244 = n14243 ^ n13322;
  assign n14613 = n14429 ^ n14244;
  assign n14671 = n14613 ^ n12180;
  assign n14835 = n14747 ^ n14671;
  assign n15709 = n15708 ^ n14835;
  assign n15502 = n13903 ^ n13162;
  assign n15026 = n14386 ^ n14353;
  assign n15503 = n15502 ^ n15026;
  assign n14818 = n14150 ^ n14096;
  assign n14816 = n13461 ^ n12861;
  assign n14817 = n14816 ^ n14246;
  assign n14819 = n14818 ^ n14817;
  assign n14711 = n14147 ^ n14144;
  assign n14697 = n14139 ^ n14098;
  assign n14695 = n14256 ^ n12871;
  assign n14696 = n14695 ^ n13471;
  assign n14698 = n14697 ^ n14696;
  assign n14658 = n14136 ^ n1973;
  assign n14589 = n14131 ^ n14100;
  assign n14587 = n13481 ^ n12877;
  assign n14588 = n14587 ^ n14202;
  assign n14590 = n14589 ^ n14588;
  assign n14580 = n14128 ^ n14102;
  assign n14237 = n13388 ^ n12890;
  assign n14238 = n14237 ^ n14051;
  assign n14236 = n14125 ^ n14104;
  assign n14239 = n14238 ^ n14236;
  assign n14570 = n14122 ^ n14106;
  assign n14563 = n14119 ^ n1459;
  assign n14549 = n14111 ^ n14110;
  assign n14531 = n13856 ^ n2383;
  assign n14528 = n12630 ^ n12030;
  assign n14529 = ~n13273 & ~n14528;
  assign n14530 = n14529 ^ n12030;
  assign n14532 = n14531 ^ n14530;
  assign n14498 = n13851 ^ n13759;
  assign n14446 = n13845 ^ n13763;
  assign n14442 = n12598 ^ n11920;
  assign n14443 = n13160 & ~n14442;
  assign n14444 = n14443 ^ n11920;
  assign n14468 = n14446 ^ n14444;
  assign n14438 = n14422 ^ n14420;
  assign n14439 = n14422 ^ n14417;
  assign n14440 = ~n14438 & n14439;
  assign n14441 = n14440 ^ n14420;
  assign n14469 = n14446 ^ n14441;
  assign n14470 = ~n14468 & ~n14469;
  assign n14471 = n14470 ^ n14444;
  assign n14467 = n13848 ^ n13761;
  assign n14472 = n14471 ^ n14467;
  assign n14464 = n12590 ^ n11968;
  assign n14465 = n13194 & n14464;
  assign n14466 = n14465 ^ n11968;
  assign n14495 = n14467 ^ n14466;
  assign n14496 = ~n14472 & n14495;
  assign n14497 = n14496 ^ n14466;
  assign n14499 = n14498 ^ n14497;
  assign n14492 = n12066 ^ n11990;
  assign n14493 = ~n13235 & ~n14492;
  assign n14494 = n14493 ^ n11990;
  assign n14524 = n14498 ^ n14494;
  assign n14525 = ~n14499 & ~n14524;
  assign n14526 = n14525 ^ n14494;
  assign n14527 = n14526 ^ n10678;
  assign n14533 = n14532 ^ n14527;
  assign n14500 = n14499 ^ n14494;
  assign n14473 = n14472 ^ n14466;
  assign n14474 = n14473 ^ n11292;
  assign n14445 = n14444 ^ n14441;
  assign n14447 = n14446 ^ n14445;
  assign n14448 = n14447 ^ n11323;
  assign n14435 = n14423 ^ n14413;
  assign n14436 = n14424 & n14435;
  assign n14437 = n14436 ^ n11295;
  assign n14461 = n14447 ^ n14437;
  assign n14462 = ~n14448 & ~n14461;
  assign n14463 = n14462 ^ n11323;
  assign n14488 = n14473 ^ n14463;
  assign n14489 = n14474 & n14488;
  assign n14490 = n14489 ^ n11292;
  assign n14491 = n14490 ^ n10684;
  assign n14501 = n14500 ^ n14491;
  assign n14449 = n14448 ^ n14437;
  assign n14450 = ~n14425 & ~n14426;
  assign n14460 = ~n14449 & n14450;
  assign n14475 = n14474 ^ n14463;
  assign n14502 = ~n14460 & n14475;
  assign n14523 = ~n14501 & ~n14502;
  assign n14534 = n14533 ^ n14523;
  assign n14519 = n14500 ^ n10684;
  assign n14520 = n14500 ^ n14490;
  assign n14521 = ~n14519 & n14520;
  assign n14522 = n14521 ^ n10684;
  assign n14535 = n14534 ^ n14522;
  assign n14503 = n14502 ^ n14501;
  assign n14476 = n14475 ^ n14460;
  assign n14477 = n14476 ^ n2589;
  assign n14451 = n14450 ^ n14449;
  assign n14432 = n14427 ^ n1538;
  assign n14433 = n14428 & ~n14432;
  assign n14434 = n14433 ^ n1538;
  assign n14452 = n14451 ^ n14434;
  assign n14457 = n14451 ^ n2426;
  assign n14458 = ~n14452 & n14457;
  assign n14459 = n14458 ^ n2426;
  assign n14485 = n14476 ^ n14459;
  assign n14486 = ~n14477 & n14485;
  assign n14487 = n14486 ^ n2589;
  assign n14504 = n14503 ^ n14487;
  assign n14512 = n14503 ^ n2616;
  assign n14513 = n14504 & ~n14512;
  assign n14514 = n14513 ^ n2616;
  assign n14518 = n14517 ^ n14514;
  assign n14536 = n14535 ^ n14518;
  assign n14505 = n14504 ^ n2616;
  assign n14478 = n14477 ^ n14459;
  assign n14430 = n14244 & ~n14429;
  assign n14241 = n13380 ^ n12057;
  assign n14242 = n14241 ^ n13424;
  assign n14431 = n14430 ^ n14242;
  assign n14453 = n14452 ^ n2426;
  assign n14454 = n14453 ^ n14242;
  assign n14455 = ~n14431 & n14454;
  assign n14456 = n14455 ^ n14430;
  assign n14479 = n14478 ^ n14456;
  assign n14480 = n13436 ^ n12050;
  assign n14481 = n14480 ^ n13418;
  assign n14482 = n14481 ^ n14478;
  assign n14483 = n14479 & ~n14482;
  assign n14484 = n14483 ^ n14481;
  assign n14506 = n14505 ^ n14484;
  assign n14507 = n13431 ^ n12044;
  assign n14508 = n14507 ^ n13416;
  assign n14509 = n14508 ^ n14505;
  assign n14510 = n14506 & ~n14509;
  assign n14511 = n14510 ^ n14508;
  assign n14537 = n14536 ^ n14511;
  assign n14538 = n13425 ^ n12038;
  assign n14539 = n14538 ^ n13410;
  assign n14540 = n14539 ^ n14536;
  assign n14541 = ~n14537 & ~n14540;
  assign n14542 = n14541 ^ n14539;
  assign n14240 = n14064 ^ n1490;
  assign n14543 = n14542 ^ n14240;
  assign n14544 = n13419 ^ n12812;
  assign n14545 = n14544 ^ n13404;
  assign n14546 = n14545 ^ n14240;
  assign n14547 = n14543 & ~n14546;
  assign n14548 = n14547 ^ n14545;
  assign n14550 = n14549 ^ n14548;
  assign n14551 = n13412 ^ n12835;
  assign n14552 = n14551 ^ n13398;
  assign n14553 = n14552 ^ n14549;
  assign n14554 = ~n14550 & ~n14553;
  assign n14555 = n14554 ^ n14552;
  assign n14557 = n14556 ^ n14555;
  assign n14558 = n13406 ^ n12905;
  assign n14559 = n14558 ^ n13392;
  assign n14560 = n14559 ^ n14556;
  assign n14561 = n14557 & ~n14560;
  assign n14562 = n14561 ^ n14559;
  assign n14564 = n14563 ^ n14562;
  assign n14565 = n13400 ^ n12900;
  assign n14566 = n14565 ^ n13386;
  assign n14567 = n14566 ^ n14563;
  assign n14568 = ~n14564 & ~n14567;
  assign n14569 = n14568 ^ n14566;
  assign n14571 = n14570 ^ n14569;
  assign n14572 = n13394 ^ n12895;
  assign n14573 = n14572 ^ n13967;
  assign n14574 = n14573 ^ n14570;
  assign n14575 = ~n14571 & n14574;
  assign n14576 = n14575 ^ n14573;
  assign n14577 = n14576 ^ n14236;
  assign n14578 = n14239 & n14577;
  assign n14579 = n14578 ^ n14238;
  assign n14581 = n14580 ^ n14579;
  assign n14582 = n12882 ^ n12845;
  assign n14583 = n14582 ^ n14183;
  assign n14584 = n14583 ^ n14580;
  assign n14585 = n14581 & ~n14584;
  assign n14586 = n14585 ^ n14583;
  assign n14655 = n14589 ^ n14586;
  assign n14656 = n14590 & n14655;
  assign n14657 = n14656 ^ n14588;
  assign n14659 = n14658 ^ n14657;
  assign n14653 = n13476 ^ n12846;
  assign n14654 = n14653 ^ n14227;
  assign n14692 = n14658 ^ n14654;
  assign n14693 = ~n14659 & ~n14692;
  assign n14694 = n14693 ^ n14654;
  assign n14708 = n14697 ^ n14694;
  assign n14709 = n14698 & n14708;
  assign n14710 = n14709 ^ n14696;
  assign n14712 = n14711 ^ n14710;
  assign n14706 = n13466 ^ n12866;
  assign n14707 = n14706 ^ n14254;
  assign n14813 = n14711 ^ n14707;
  assign n14814 = ~n14712 & n14813;
  assign n14815 = n14814 ^ n14707;
  assign n14820 = n14819 ^ n14815;
  assign n14821 = n14820 ^ n12098;
  assign n14713 = n14712 ^ n14707;
  assign n14714 = n14713 ^ n12104;
  assign n14699 = n14698 ^ n14694;
  assign n14700 = n14699 ^ n12109;
  assign n14660 = n14659 ^ n14654;
  assign n14661 = n14660 ^ n12115;
  assign n14591 = n14590 ^ n14586;
  assign n14592 = n14591 ^ n12120;
  assign n14593 = n14583 ^ n14581;
  assign n14594 = n14593 ^ n12129;
  assign n14595 = n14576 ^ n14239;
  assign n14596 = n14595 ^ n12134;
  assign n14597 = n14573 ^ n14571;
  assign n14598 = n14597 ^ n11495;
  assign n14599 = n14566 ^ n14564;
  assign n14600 = n14599 ^ n12040;
  assign n14601 = n14559 ^ n14557;
  assign n14602 = n14601 ^ n12046;
  assign n14603 = n14552 ^ n14550;
  assign n14604 = n14603 ^ n12053;
  assign n14605 = n14545 ^ n14543;
  assign n14606 = n14605 ^ n12061;
  assign n14607 = n14539 ^ n14537;
  assign n14608 = n14607 ^ n12159;
  assign n14609 = n14508 ^ n14506;
  assign n14610 = n14609 ^ n12068;
  assign n14611 = n14481 ^ n14479;
  assign n14612 = n14611 ^ n12168;
  assign n14614 = n12180 & ~n14613;
  assign n14615 = n14614 ^ n12174;
  assign n14616 = n14453 ^ n14431;
  assign n14617 = n14616 ^ n14614;
  assign n14618 = ~n14615 & n14617;
  assign n14619 = n14618 ^ n12174;
  assign n14620 = n14619 ^ n14611;
  assign n14621 = n14612 & ~n14620;
  assign n14622 = n14621 ^ n12168;
  assign n14623 = n14622 ^ n14609;
  assign n14624 = ~n14610 & ~n14623;
  assign n14625 = n14624 ^ n12068;
  assign n14626 = n14625 ^ n14607;
  assign n14627 = ~n14608 & n14626;
  assign n14628 = n14627 ^ n12159;
  assign n14629 = n14628 ^ n14605;
  assign n14630 = n14606 & ~n14629;
  assign n14631 = n14630 ^ n12061;
  assign n14632 = n14631 ^ n14603;
  assign n14633 = n14604 & ~n14632;
  assign n14634 = n14633 ^ n12053;
  assign n14635 = n14634 ^ n14601;
  assign n14636 = n14602 & n14635;
  assign n14637 = n14636 ^ n12046;
  assign n14638 = n14637 ^ n14599;
  assign n14639 = ~n14600 & ~n14638;
  assign n14640 = n14639 ^ n12040;
  assign n14641 = n14640 ^ n14597;
  assign n14642 = ~n14598 & n14641;
  assign n14643 = n14642 ^ n11495;
  assign n14644 = n14643 ^ n14595;
  assign n14645 = ~n14596 & n14644;
  assign n14646 = n14645 ^ n12134;
  assign n14647 = n14646 ^ n14593;
  assign n14648 = ~n14594 & n14647;
  assign n14649 = n14648 ^ n12129;
  assign n14650 = n14649 ^ n14591;
  assign n14651 = n14592 & ~n14650;
  assign n14652 = n14651 ^ n12120;
  assign n14689 = n14660 ^ n14652;
  assign n14690 = ~n14661 & ~n14689;
  assign n14691 = n14690 ^ n12115;
  assign n14703 = n14699 ^ n14691;
  assign n14704 = n14700 & n14703;
  assign n14705 = n14704 ^ n12109;
  assign n14810 = n14713 ^ n14705;
  assign n14811 = n14714 & n14810;
  assign n14812 = n14811 ^ n12104;
  assign n14944 = n14820 ^ n14812;
  assign n14945 = ~n14821 & n14944;
  assign n14946 = n14945 ^ n12098;
  assign n14860 = n14818 ^ n14815;
  assign n14861 = ~n14819 & ~n14860;
  assign n14862 = n14861 ^ n14817;
  assign n14858 = n14158 ^ n14155;
  assign n14856 = n13456 ^ n12856;
  assign n14857 = n14856 ^ n14245;
  assign n14859 = n14858 ^ n14857;
  assign n14942 = n14862 ^ n14859;
  assign n14943 = n14942 ^ n12093;
  assign n14996 = n14946 ^ n14943;
  assign n14822 = n14821 ^ n14812;
  assign n14662 = n14661 ^ n14652;
  assign n14663 = n14649 ^ n14592;
  assign n14664 = n14646 ^ n14594;
  assign n14665 = n14640 ^ n14598;
  assign n14666 = n14637 ^ n14600;
  assign n14667 = n14631 ^ n14604;
  assign n14668 = n14625 ^ n14608;
  assign n14669 = n14622 ^ n14610;
  assign n14670 = n14619 ^ n14612;
  assign n14672 = n14616 ^ n14615;
  assign n14673 = ~n14671 & n14672;
  assign n14674 = ~n14670 & n14673;
  assign n14675 = n14669 & n14674;
  assign n14676 = ~n14668 & n14675;
  assign n14677 = n14628 ^ n14606;
  assign n14678 = ~n14676 & ~n14677;
  assign n14679 = n14667 & ~n14678;
  assign n14680 = n14634 ^ n14602;
  assign n14681 = ~n14679 & ~n14680;
  assign n14682 = ~n14666 & n14681;
  assign n14683 = n14665 & n14682;
  assign n14684 = n14643 ^ n14596;
  assign n14685 = ~n14683 & ~n14684;
  assign n14686 = n14664 & ~n14685;
  assign n14687 = n14663 & ~n14686;
  assign n14688 = n14662 & ~n14687;
  assign n14701 = n14700 ^ n14691;
  assign n14702 = n14688 & n14701;
  assign n14715 = n14714 ^ n14705;
  assign n14823 = n14702 & ~n14715;
  assign n14997 = ~n14822 & n14823;
  assign n14998 = n14996 & ~n14997;
  assign n14947 = n14946 ^ n14942;
  assign n14948 = ~n14943 & n14947;
  assign n14949 = n14948 ^ n12093;
  assign n14868 = n13451 ^ n12947;
  assign n14869 = n14868 ^ n14234;
  assign n14866 = n14161 ^ n14091;
  assign n14863 = n14862 ^ n14858;
  assign n14864 = n14859 & n14863;
  assign n14865 = n14864 ^ n14857;
  assign n14867 = n14866 ^ n14865;
  assign n14940 = n14869 ^ n14867;
  assign n14941 = n14940 ^ n12087;
  assign n14999 = n14949 ^ n14941;
  assign n15000 = n14998 & n14999;
  assign n14950 = n14949 ^ n14940;
  assign n14951 = ~n14941 & ~n14950;
  assign n14952 = n14951 ^ n12087;
  assign n14870 = n14869 ^ n14866;
  assign n14871 = n14867 & n14870;
  assign n14872 = n14871 ^ n14869;
  assign n14853 = n13446 ^ n13023;
  assign n14854 = n14853 ^ n14288;
  assign n14852 = n14166 ^ n575;
  assign n14855 = n14854 ^ n14852;
  assign n14938 = n14872 ^ n14855;
  assign n14939 = n14938 ^ n12081;
  assign n14995 = n14952 ^ n14939;
  assign n15055 = n15000 ^ n14995;
  assign n15042 = n14999 ^ n14998;
  assign n15043 = n15042 ^ n568;
  assign n15044 = n14997 ^ n14996;
  assign n15045 = n15044 ^ n562;
  assign n14824 = n14823 ^ n14822;
  assign n14825 = n14824 ^ n656;
  assign n14716 = n14715 ^ n14702;
  assign n14717 = n14716 ^ n650;
  assign n14799 = n14701 ^ n14688;
  assign n14718 = n14687 ^ n14662;
  assign n14722 = n14721 ^ n14718;
  assign n14723 = n14686 ^ n14663;
  assign n14727 = n14726 ^ n14723;
  assign n14728 = n14685 ^ n14664;
  assign n14732 = n14731 ^ n14728;
  assign n14785 = n14684 ^ n14683;
  assign n14733 = n14682 ^ n14665;
  assign n14734 = n14733 ^ n2235;
  assign n14777 = n14681 ^ n14666;
  assign n14735 = n14680 ^ n14679;
  assign n14736 = n14735 ^ n1814;
  assign n14737 = n14678 ^ n14667;
  assign n14738 = n14737 ^ n1817;
  assign n14766 = n14677 ^ n14676;
  assign n14739 = n14675 ^ n14668;
  assign n14740 = n14739 ^ n1635;
  assign n14741 = n14674 ^ n14669;
  assign n14742 = n14741 ^ n1613;
  assign n14743 = n14673 ^ n14670;
  assign n14744 = n14743 ^ n1607;
  assign n14748 = n14671 & n14747;
  assign n14752 = n14751 ^ n14748;
  assign n14753 = n14672 ^ n14671;
  assign n14754 = n14753 ^ n14748;
  assign n14755 = n14752 & n14754;
  assign n14756 = n14755 ^ n14751;
  assign n14757 = n14756 ^ n14743;
  assign n14758 = ~n14744 & n14757;
  assign n14759 = n14758 ^ n1607;
  assign n14760 = n14759 ^ n14741;
  assign n14761 = n14742 & ~n14760;
  assign n14762 = n14761 ^ n1613;
  assign n14763 = n14762 ^ n14739;
  assign n14764 = ~n14740 & n14763;
  assign n14765 = n14764 ^ n1635;
  assign n14767 = n14766 ^ n14765;
  assign n14768 = n14766 ^ n1703;
  assign n14769 = n14767 & ~n14768;
  assign n14770 = n14769 ^ n1703;
  assign n14771 = n14770 ^ n14737;
  assign n14772 = ~n14738 & n14771;
  assign n14773 = n14772 ^ n1817;
  assign n14774 = n14773 ^ n14735;
  assign n14775 = ~n14736 & n14774;
  assign n14776 = n14775 ^ n1814;
  assign n14778 = n14777 ^ n14776;
  assign n14779 = n14777 ^ n1986;
  assign n14780 = ~n14778 & n14779;
  assign n14781 = n14780 ^ n1986;
  assign n14782 = n14781 ^ n14733;
  assign n14783 = ~n14734 & n14782;
  assign n14784 = n14783 ^ n2235;
  assign n14786 = n14785 ^ n14784;
  assign n14787 = n14785 ^ n581;
  assign n14788 = ~n14786 & n14787;
  assign n14789 = n14788 ^ n581;
  assign n14790 = n14789 ^ n14728;
  assign n14791 = n14732 & ~n14790;
  assign n14792 = n14791 ^ n14731;
  assign n14793 = n14792 ^ n14723;
  assign n14794 = ~n14727 & n14793;
  assign n14795 = n14794 ^ n14726;
  assign n14796 = n14795 ^ n14718;
  assign n14797 = n14722 & ~n14796;
  assign n14798 = n14797 ^ n14721;
  assign n14800 = n14799 ^ n14798;
  assign n14804 = n14803 ^ n14799;
  assign n14805 = n14800 & ~n14804;
  assign n14806 = n14805 ^ n14803;
  assign n14807 = n14806 ^ n14716;
  assign n14808 = n14717 & ~n14807;
  assign n14809 = n14808 ^ n650;
  assign n15046 = n14824 ^ n14809;
  assign n15047 = n14825 & ~n15046;
  assign n15048 = n15047 ^ n656;
  assign n15049 = n15048 ^ n15044;
  assign n15050 = ~n15045 & n15049;
  assign n15051 = n15050 ^ n562;
  assign n15052 = n15051 ^ n15042;
  assign n15053 = n15043 & ~n15052;
  assign n15054 = n15053 ^ n568;
  assign n15056 = n15055 ^ n15054;
  assign n15057 = n15055 ^ n756;
  assign n15058 = ~n15056 & n15057;
  assign n15059 = n15058 ^ n756;
  assign n14953 = n14952 ^ n14938;
  assign n14954 = ~n14939 & ~n14953;
  assign n14955 = n14954 ^ n12081;
  assign n14873 = n14872 ^ n14852;
  assign n14874 = n14855 & n14873;
  assign n14875 = n14874 ^ n14854;
  assign n14848 = n13585 ^ n13065;
  assign n14849 = n14848 ^ n14334;
  assign n14935 = n14875 ^ n14849;
  assign n14850 = n14169 ^ n14089;
  assign n14936 = n14935 ^ n14850;
  assign n14937 = n14936 ^ n12075;
  assign n15002 = n14955 ^ n14937;
  assign n15001 = n14995 & ~n15000;
  assign n15040 = n15002 ^ n15001;
  assign n15041 = n15040 ^ n1083;
  assign n15501 = n15059 ^ n15041;
  assign n15504 = n15503 ^ n15501;
  assign n15423 = n15056 ^ n756;
  assign n15421 = n14531 ^ n13930;
  assign n14988 = n14383 ^ n14355;
  assign n15422 = n15421 ^ n14988;
  assign n15424 = n15423 ^ n15422;
  assign n15414 = n15051 ^ n15043;
  assign n15331 = n14467 ^ n13749;
  assign n14838 = n14377 ^ n975;
  assign n15332 = n15331 ^ n14838;
  assign n15330 = n15048 ^ n15045;
  assign n15333 = n15332 ^ n15330;
  assign n15334 = n14446 ^ n13695;
  assign n14904 = n14372 ^ n14359;
  assign n15335 = n15334 ^ n14904;
  assign n14826 = n14825 ^ n14809;
  assign n15336 = n15335 ^ n14826;
  assign n15401 = n14806 ^ n14717;
  assign n15338 = n14401 ^ n13446;
  assign n14839 = n14364 ^ n14361;
  assign n15339 = n15338 ^ n14839;
  assign n15337 = n14803 ^ n14800;
  assign n15340 = n15339 ^ n15337;
  assign n15391 = n14795 ^ n14722;
  assign n15342 = n14288 ^ n13456;
  assign n14842 = n14212 ^ n542;
  assign n15343 = n15342 ^ n14842;
  assign n15341 = n14792 ^ n14727;
  assign n15344 = n15343 ^ n15341;
  assign n15347 = n14789 ^ n14732;
  assign n15345 = n14234 ^ n13461;
  assign n14846 = n14192 ^ n14189;
  assign n15346 = n15345 ^ n14846;
  assign n15348 = n15347 ^ n15346;
  assign n15378 = n14786 ^ n581;
  assign n15350 = n14246 ^ n13471;
  assign n15351 = n15350 ^ n14852;
  assign n15349 = n14781 ^ n14734;
  assign n15352 = n15351 ^ n15349;
  assign n15354 = n14256 ^ n13481;
  assign n15355 = n15354 ^ n14858;
  assign n15353 = n14773 ^ n14736;
  assign n15356 = n15355 ^ n15353;
  assign n15300 = n14767 ^ n1703;
  assign n15298 = n14202 ^ n13388;
  assign n15299 = n15298 ^ n14711;
  assign n15301 = n15300 ^ n15299;
  assign n15236 = n14762 ^ n1635;
  assign n15237 = n15236 ^ n14739;
  assign n15206 = n14051 ^ n13400;
  assign n15207 = n15206 ^ n14658;
  assign n15205 = n14759 ^ n14742;
  assign n15208 = n15207 ^ n15205;
  assign n14832 = n13412 ^ n13386;
  assign n14833 = n14832 ^ n14580;
  assign n14831 = n14753 ^ n14752;
  assign n14834 = n14833 ^ n14831;
  assign n15123 = n13425 ^ n13398;
  assign n15124 = n15123 ^ n14570;
  assign n14917 = n14380 ^ n14357;
  assign n14897 = n14369 ^ n859;
  assign n14840 = n13749 ^ n13179;
  assign n14841 = n14840 ^ n14422;
  assign n14843 = n14842 ^ n14841;
  assign n14844 = n13695 ^ n13143;
  assign n14845 = n14844 ^ n14401;
  assign n14847 = n14846 ^ n14845;
  assign n14851 = n14850 ^ n14849;
  assign n14876 = n14875 ^ n14850;
  assign n14877 = n14851 & n14876;
  assign n14878 = n14877 ^ n14849;
  assign n14879 = n14878 ^ n14846;
  assign n14880 = n14847 & ~n14879;
  assign n14881 = n14880 ^ n14845;
  assign n14882 = n14881 ^ n14841;
  assign n14883 = ~n14843 & n14882;
  assign n14884 = n14883 ^ n14842;
  assign n14233 = n14232 ^ n14215;
  assign n14885 = n14884 ^ n14233;
  assign n14886 = n13881 ^ n13222;
  assign n14887 = n14886 ^ n14446;
  assign n14888 = n14887 ^ n14233;
  assign n14889 = n14885 & n14888;
  assign n14890 = n14889 ^ n14887;
  assign n14891 = n14890 ^ n14839;
  assign n14892 = n13930 ^ n13264;
  assign n14893 = n14892 ^ n14467;
  assign n14894 = n14893 ^ n14839;
  assign n14895 = n14891 & ~n14894;
  assign n14896 = n14895 ^ n14893;
  assign n14898 = n14897 ^ n14896;
  assign n14899 = n13162 ^ n12605;
  assign n14900 = n14899 ^ n14498;
  assign n14901 = n14900 ^ n14897;
  assign n14902 = ~n14898 & ~n14901;
  assign n14903 = n14902 ^ n14900;
  assign n14905 = n14904 ^ n14903;
  assign n14906 = n13160 ^ n12600;
  assign n14907 = n14906 ^ n14531;
  assign n14908 = n14907 ^ n14904;
  assign n14909 = n14905 & n14908;
  assign n14910 = n14909 ^ n14907;
  assign n14911 = n14910 ^ n14838;
  assign n14912 = n13194 ^ n12617;
  assign n14913 = n14912 ^ n13903;
  assign n14914 = n14913 ^ n14838;
  assign n14915 = ~n14911 & n14914;
  assign n14916 = n14915 ^ n14913;
  assign n14918 = n14917 ^ n14916;
  assign n14836 = n13235 ^ n12598;
  assign n14837 = n14836 ^ n13898;
  assign n14985 = n14917 ^ n14837;
  assign n14986 = ~n14918 & n14985;
  assign n14987 = n14986 ^ n14837;
  assign n14989 = n14988 ^ n14987;
  assign n14983 = n13273 ^ n12590;
  assign n14984 = n14983 ^ n13893;
  assign n14990 = n14989 ^ n14984;
  assign n14991 = n14990 ^ n11968;
  assign n14919 = n14918 ^ n14837;
  assign n14920 = n14919 ^ n11920;
  assign n14921 = n14913 ^ n14911;
  assign n14922 = n14921 ^ n11876;
  assign n14923 = n14907 ^ n14905;
  assign n14924 = n14923 ^ n11881;
  assign n14925 = n14900 ^ n14898;
  assign n14926 = n14925 ^ n11887;
  assign n14927 = n14893 ^ n14891;
  assign n14928 = n14927 ^ n12584;
  assign n14929 = n14887 ^ n14885;
  assign n14930 = n14929 ^ n12562;
  assign n14931 = n14881 ^ n14843;
  assign n14932 = n14931 ^ n12377;
  assign n14933 = n14878 ^ n14847;
  assign n14934 = n14933 ^ n12074;
  assign n14956 = n14955 ^ n14936;
  assign n14957 = ~n14937 & ~n14956;
  assign n14958 = n14957 ^ n12075;
  assign n14959 = n14958 ^ n14933;
  assign n14960 = n14934 & ~n14959;
  assign n14961 = n14960 ^ n12074;
  assign n14962 = n14961 ^ n14931;
  assign n14963 = n14932 & n14962;
  assign n14964 = n14963 ^ n12377;
  assign n14965 = n14964 ^ n14929;
  assign n14966 = n14930 & n14965;
  assign n14967 = n14966 ^ n12562;
  assign n14968 = n14967 ^ n14927;
  assign n14969 = ~n14928 & ~n14968;
  assign n14970 = n14969 ^ n12584;
  assign n14971 = n14970 ^ n14925;
  assign n14972 = ~n14926 & n14971;
  assign n14973 = n14972 ^ n11887;
  assign n14974 = n14973 ^ n14923;
  assign n14975 = n14924 & n14974;
  assign n14976 = n14975 ^ n11881;
  assign n14977 = n14976 ^ n14921;
  assign n14978 = ~n14922 & n14977;
  assign n14979 = n14978 ^ n11876;
  assign n14980 = n14979 ^ n14919;
  assign n14981 = n14920 & n14980;
  assign n14982 = n14981 ^ n11920;
  assign n14992 = n14991 ^ n14982;
  assign n14993 = n14976 ^ n14922;
  assign n14994 = n14958 ^ n14934;
  assign n15003 = n15001 & ~n15002;
  assign n15004 = n14994 & ~n15003;
  assign n15005 = n14961 ^ n14932;
  assign n15006 = ~n15004 & ~n15005;
  assign n15007 = n14964 ^ n14930;
  assign n15008 = n15006 & n15007;
  assign n15009 = n14967 ^ n14928;
  assign n15010 = ~n15008 & ~n15009;
  assign n15011 = n14970 ^ n14926;
  assign n15012 = ~n15010 & ~n15011;
  assign n15013 = n14973 ^ n14924;
  assign n15014 = n15012 & n15013;
  assign n15015 = n14993 & n15014;
  assign n15016 = n14979 ^ n14920;
  assign n15017 = ~n15015 & n15016;
  assign n15018 = ~n14992 & ~n15017;
  assign n15028 = n13295 ^ n12066;
  assign n15029 = n15028 ^ n13888;
  assign n15023 = n14988 ^ n14984;
  assign n15024 = ~n14989 & ~n15023;
  assign n15025 = n15024 ^ n14984;
  assign n15027 = n15026 ^ n15025;
  assign n15030 = n15029 ^ n15027;
  assign n15019 = n14990 ^ n14982;
  assign n15020 = ~n14991 & n15019;
  assign n15021 = n15020 ^ n11968;
  assign n15022 = n15021 ^ n11990;
  assign n15031 = n15030 ^ n15022;
  assign n15120 = n15018 & ~n15031;
  assign n15115 = n13310 ^ n12630;
  assign n15116 = n15115 ^ n13936;
  assign n15112 = n15029 ^ n15026;
  assign n15113 = n15027 & ~n15112;
  assign n15114 = n15113 ^ n15029;
  assign n15117 = n15116 ^ n15114;
  assign n15111 = n14407 ^ n2309;
  assign n15118 = n15117 ^ n15111;
  assign n15106 = n15030 ^ n11990;
  assign n15107 = n15030 ^ n15021;
  assign n15108 = ~n15106 & ~n15107;
  assign n15109 = n15108 ^ n11990;
  assign n15110 = n15109 ^ n12030;
  assign n15119 = n15118 ^ n15110;
  assign n15121 = n15120 ^ n15119;
  assign n15032 = n15031 ^ n15018;
  assign n15033 = n15032 ^ n2639;
  assign n15097 = n15017 ^ n14992;
  assign n15092 = n15016 ^ n15015;
  assign n15087 = n15014 ^ n14993;
  assign n15082 = n15013 ^ n15012;
  assign n15034 = n15011 ^ n15010;
  assign n15035 = n15034 ^ n2286;
  assign n15036 = n15009 ^ n15008;
  assign n1241 = n1144 ^ x200;
  assign n1242 = n1241 ^ x392;
  assign n1243 = n1242 ^ x136;
  assign n15037 = n15036 ^ n1243;
  assign n15071 = n15007 ^ n15006;
  assign n15038 = n15005 ^ n15004;
  assign n15039 = n15038 ^ n1075;
  assign n15063 = n15003 ^ n14994;
  assign n15060 = n15059 ^ n15040;
  assign n15061 = n15041 & ~n15060;
  assign n15062 = n15061 ^ n1083;
  assign n15064 = n15063 ^ n15062;
  assign n15065 = n15063 ^ n901;
  assign n15066 = n15064 & ~n15065;
  assign n15067 = n15066 ^ n901;
  assign n15068 = n15067 ^ n15038;
  assign n15069 = ~n15039 & n15068;
  assign n15070 = n15069 ^ n1075;
  assign n15072 = n15071 ^ n15070;
  assign n15073 = n15071 ^ n1105;
  assign n15074 = n15072 & ~n15073;
  assign n15075 = n15074 ^ n1105;
  assign n15076 = n15075 ^ n15036;
  assign n15077 = n15037 & ~n15076;
  assign n15078 = n15077 ^ n1243;
  assign n15079 = n15078 ^ n15034;
  assign n15080 = ~n15035 & n15079;
  assign n15081 = n15080 ^ n2286;
  assign n15083 = n15082 ^ n15081;
  assign n15084 = n15082 ^ n2294;
  assign n15085 = n15083 & ~n15084;
  assign n15086 = n15085 ^ n2294;
  assign n15088 = n15087 ^ n15086;
  assign n15089 = n15087 ^ n2356;
  assign n15090 = n15088 & ~n15089;
  assign n15091 = n15090 ^ n2356;
  assign n15093 = n15092 ^ n15091;
  assign n2482 = n2414 ^ x196;
  assign n2483 = n2482 ^ x388;
  assign n2484 = n2483 ^ x132;
  assign n15094 = n15092 ^ n2484;
  assign n15095 = n15093 & ~n15094;
  assign n15096 = n15095 ^ n2484;
  assign n15098 = n15097 ^ n15096;
  assign n15099 = n15097 ^ n1514;
  assign n15100 = n15098 & ~n15099;
  assign n15101 = n15100 ^ n1514;
  assign n15102 = n15101 ^ n15032;
  assign n15103 = n15033 & ~n15102;
  assign n15104 = n15103 ^ n2639;
  assign n15105 = n15104 ^ n1427;
  assign n15122 = n15121 ^ n15105;
  assign n15125 = n15124 ^ n15122;
  assign n15144 = n15101 ^ n2639;
  assign n15145 = n15144 ^ n15032;
  assign n15137 = n15098 ^ n1514;
  assign n15128 = n15088 ^ n2356;
  assign n15129 = n13418 ^ n13322;
  assign n15130 = n15129 ^ n14240;
  assign n15131 = ~n15128 & ~n15130;
  assign n15126 = n13416 ^ n13380;
  assign n15127 = n15126 ^ n14549;
  assign n15132 = n15131 ^ n15127;
  assign n15133 = n15093 ^ n2484;
  assign n15134 = n15133 ^ n15127;
  assign n15135 = n15132 & n15134;
  assign n15136 = n15135 ^ n15131;
  assign n15138 = n15137 ^ n15136;
  assign n15139 = n14556 ^ n13436;
  assign n15140 = n15139 ^ n13410;
  assign n15141 = n15140 ^ n15137;
  assign n15142 = n15138 & n15141;
  assign n15143 = n15142 ^ n15140;
  assign n15146 = n15145 ^ n15143;
  assign n15147 = n13431 ^ n13404;
  assign n15148 = n15147 ^ n14563;
  assign n15149 = n15148 ^ n15145;
  assign n15150 = n15146 & ~n15149;
  assign n15151 = n15150 ^ n15148;
  assign n15152 = n15151 ^ n15122;
  assign n15153 = ~n15125 & ~n15152;
  assign n15154 = n15153 ^ n15124;
  assign n15155 = n15154 ^ n14835;
  assign n15156 = n13419 ^ n13392;
  assign n15157 = n15156 ^ n14236;
  assign n15158 = n15157 ^ n14835;
  assign n15159 = ~n15155 & n15158;
  assign n15160 = n15159 ^ n15157;
  assign n15161 = n15160 ^ n14831;
  assign n15162 = n14834 & n15161;
  assign n15163 = n15162 ^ n14833;
  assign n14830 = n14756 ^ n14744;
  assign n15164 = n15163 ^ n14830;
  assign n14828 = n13967 ^ n13406;
  assign n14829 = n14828 ^ n14589;
  assign n15202 = n14830 ^ n14829;
  assign n15203 = ~n15164 & n15202;
  assign n15204 = n15203 ^ n14829;
  assign n15233 = n15205 ^ n15204;
  assign n15234 = n15208 & n15233;
  assign n15235 = n15234 ^ n15207;
  assign n15238 = n15237 ^ n15235;
  assign n15231 = n14183 ^ n13394;
  assign n15232 = n15231 ^ n14697;
  assign n15295 = n15237 ^ n15232;
  assign n15296 = n15238 & n15295;
  assign n15297 = n15296 ^ n15232;
  assign n15357 = n15300 ^ n15297;
  assign n15358 = n15301 & ~n15357;
  assign n15359 = n15358 ^ n15299;
  assign n15325 = n14770 ^ n14738;
  assign n15360 = n15359 ^ n15325;
  assign n15361 = n14227 ^ n12845;
  assign n15362 = n15361 ^ n14818;
  assign n15363 = n15362 ^ n15325;
  assign n15364 = ~n15360 & n15363;
  assign n15365 = n15364 ^ n15362;
  assign n15366 = n15365 ^ n15353;
  assign n15367 = ~n15356 & ~n15366;
  assign n15368 = n15367 ^ n15355;
  assign n15319 = n14778 ^ n1986;
  assign n15369 = n15368 ^ n15319;
  assign n15370 = n14254 ^ n13476;
  assign n15371 = n15370 ^ n14866;
  assign n15372 = n15371 ^ n15319;
  assign n15373 = ~n15369 & ~n15372;
  assign n15374 = n15373 ^ n15371;
  assign n15375 = n15374 ^ n15349;
  assign n15376 = n15352 & ~n15375;
  assign n15377 = n15376 ^ n15351;
  assign n15379 = n15378 ^ n15377;
  assign n15380 = n14245 ^ n13466;
  assign n15381 = n15380 ^ n14850;
  assign n15382 = n15381 ^ n15378;
  assign n15383 = n15379 & ~n15382;
  assign n15384 = n15383 ^ n15381;
  assign n15385 = n15384 ^ n15347;
  assign n15386 = n15348 & n15385;
  assign n15387 = n15386 ^ n15346;
  assign n15388 = n15387 ^ n15341;
  assign n15389 = ~n15344 & n15388;
  assign n15390 = n15389 ^ n15343;
  assign n15392 = n15391 ^ n15390;
  assign n15393 = n14334 ^ n13451;
  assign n15394 = n15393 ^ n14233;
  assign n15395 = n15394 ^ n15391;
  assign n15396 = ~n15392 & n15395;
  assign n15397 = n15396 ^ n15394;
  assign n15398 = n15397 ^ n15337;
  assign n15399 = n15340 & n15398;
  assign n15400 = n15399 ^ n15339;
  assign n15402 = n15401 ^ n15400;
  assign n15403 = n14422 ^ n13585;
  assign n15404 = n15403 ^ n14897;
  assign n15405 = n15404 ^ n15401;
  assign n15406 = n15402 & ~n15405;
  assign n15407 = n15406 ^ n15404;
  assign n15408 = n15407 ^ n14826;
  assign n15409 = n15336 & n15408;
  assign n15410 = n15409 ^ n15335;
  assign n15411 = n15410 ^ n15330;
  assign n15412 = n15333 & n15411;
  assign n15413 = n15412 ^ n15332;
  assign n15415 = n15414 ^ n15413;
  assign n15416 = n14917 ^ n13881;
  assign n15417 = n15416 ^ n14498;
  assign n15418 = n15417 ^ n15414;
  assign n15419 = n15415 & ~n15418;
  assign n15420 = n15419 ^ n15417;
  assign n15498 = n15423 ^ n15420;
  assign n15499 = n15424 & n15498;
  assign n15500 = n15499 ^ n15422;
  assign n15544 = n15501 ^ n15500;
  assign n15545 = ~n15504 & ~n15544;
  assign n15546 = n15545 ^ n15503;
  assign n15543 = n15064 ^ n901;
  assign n15547 = n15546 ^ n15543;
  assign n15541 = n13898 ^ n13160;
  assign n15542 = n15541 ^ n15111;
  assign n15548 = n15547 ^ n15542;
  assign n15549 = n15548 ^ n12600;
  assign n15505 = n15504 ^ n15500;
  assign n15506 = n15505 ^ n12605;
  assign n15425 = n15424 ^ n15420;
  assign n15426 = n15425 ^ n13264;
  assign n15427 = n15417 ^ n15415;
  assign n15428 = n15427 ^ n13222;
  assign n15429 = n15410 ^ n15333;
  assign n15430 = n15429 ^ n13179;
  assign n15431 = n15407 ^ n15336;
  assign n15432 = n15431 ^ n13143;
  assign n15433 = n15404 ^ n15402;
  assign n15434 = n15433 ^ n13065;
  assign n15435 = n15397 ^ n15340;
  assign n15436 = n15435 ^ n13023;
  assign n15437 = n15394 ^ n15392;
  assign n15438 = n15437 ^ n12947;
  assign n15439 = n15387 ^ n15344;
  assign n15440 = n15439 ^ n12856;
  assign n15441 = n15384 ^ n15348;
  assign n15442 = n15441 ^ n12861;
  assign n15443 = n15381 ^ n15379;
  assign n15444 = n15443 ^ n12866;
  assign n15445 = n15374 ^ n15352;
  assign n15446 = n15445 ^ n12871;
  assign n15447 = n15371 ^ n15369;
  assign n15448 = n15447 ^ n12846;
  assign n15449 = n15365 ^ n15356;
  assign n15450 = n15449 ^ n12877;
  assign n15451 = n15362 ^ n15360;
  assign n15452 = n15451 ^ n12882;
  assign n15302 = n15301 ^ n15297;
  assign n15303 = n15302 ^ n12890;
  assign n15239 = n15238 ^ n15232;
  assign n15240 = n15239 ^ n12895;
  assign n15209 = n15208 ^ n15204;
  assign n15210 = n15209 ^ n12900;
  assign n15165 = n15164 ^ n14829;
  assign n15166 = n15165 ^ n12905;
  assign n15167 = n15160 ^ n14834;
  assign n15168 = n15167 ^ n12835;
  assign n15169 = n15157 ^ n15155;
  assign n15170 = n15169 ^ n12812;
  assign n15171 = n15151 ^ n15125;
  assign n15172 = n15171 ^ n12038;
  assign n15173 = n15148 ^ n15146;
  assign n15174 = n15173 ^ n12044;
  assign n15175 = n15140 ^ n15138;
  assign n15176 = n15175 ^ n12050;
  assign n15177 = n15130 ^ n15128;
  assign n15178 = ~n12059 & n15177;
  assign n15179 = n15178 ^ n12057;
  assign n15180 = n15133 ^ n15132;
  assign n15181 = n15180 ^ n15178;
  assign n15182 = n15179 & n15181;
  assign n15183 = n15182 ^ n12057;
  assign n15184 = n15183 ^ n15175;
  assign n15185 = n15176 & ~n15184;
  assign n15186 = n15185 ^ n12050;
  assign n15187 = n15186 ^ n15173;
  assign n15188 = n15174 & ~n15187;
  assign n15189 = n15188 ^ n12044;
  assign n15190 = n15189 ^ n15171;
  assign n15191 = n15172 & ~n15190;
  assign n15192 = n15191 ^ n12038;
  assign n15193 = n15192 ^ n15169;
  assign n15194 = n15170 & ~n15193;
  assign n15195 = n15194 ^ n12812;
  assign n15196 = n15195 ^ n15167;
  assign n15197 = ~n15168 & ~n15196;
  assign n15198 = n15197 ^ n12835;
  assign n15199 = n15198 ^ n15165;
  assign n15200 = n15166 & ~n15199;
  assign n15201 = n15200 ^ n12905;
  assign n15228 = n15209 ^ n15201;
  assign n15229 = n15210 & ~n15228;
  assign n15230 = n15229 ^ n12900;
  assign n15292 = n15239 ^ n15230;
  assign n15293 = n15240 & n15292;
  assign n15294 = n15293 ^ n12895;
  assign n15453 = n15302 ^ n15294;
  assign n15454 = n15303 & n15453;
  assign n15455 = n15454 ^ n12890;
  assign n15456 = n15455 ^ n15451;
  assign n15457 = ~n15452 & ~n15456;
  assign n15458 = n15457 ^ n12882;
  assign n15459 = n15458 ^ n15449;
  assign n15460 = ~n15450 & ~n15459;
  assign n15461 = n15460 ^ n12877;
  assign n15462 = n15461 ^ n15447;
  assign n15463 = ~n15448 & ~n15462;
  assign n15464 = n15463 ^ n12846;
  assign n15465 = n15464 ^ n15445;
  assign n15466 = n15446 & n15465;
  assign n15467 = n15466 ^ n12871;
  assign n15468 = n15467 ^ n15443;
  assign n15469 = n15444 & n15468;
  assign n15470 = n15469 ^ n12866;
  assign n15471 = n15470 ^ n15441;
  assign n15472 = n15442 & n15471;
  assign n15473 = n15472 ^ n12861;
  assign n15474 = n15473 ^ n15439;
  assign n15475 = n15440 & ~n15474;
  assign n15476 = n15475 ^ n12856;
  assign n15477 = n15476 ^ n15437;
  assign n15478 = n15438 & n15477;
  assign n15479 = n15478 ^ n12947;
  assign n15480 = n15479 ^ n15435;
  assign n15481 = ~n15436 & ~n15480;
  assign n15482 = n15481 ^ n13023;
  assign n15483 = n15482 ^ n15433;
  assign n15484 = n15434 & n15483;
  assign n15485 = n15484 ^ n13065;
  assign n15486 = n15485 ^ n15431;
  assign n15487 = n15432 & n15486;
  assign n15488 = n15487 ^ n13143;
  assign n15489 = n15488 ^ n15429;
  assign n15490 = ~n15430 & n15489;
  assign n15491 = n15490 ^ n13179;
  assign n15492 = n15491 ^ n15427;
  assign n15493 = n15428 & n15492;
  assign n15494 = n15493 ^ n13222;
  assign n15495 = n15494 ^ n15425;
  assign n15496 = ~n15426 & n15495;
  assign n15497 = n15496 ^ n13264;
  assign n15538 = n15505 ^ n15497;
  assign n15539 = ~n15506 & n15538;
  assign n15540 = n15539 ^ n12605;
  assign n15550 = n15549 ^ n15540;
  assign n15507 = n15506 ^ n15497;
  assign n15508 = n15482 ^ n15434;
  assign n15509 = n15476 ^ n15438;
  assign n15510 = n15467 ^ n15444;
  assign n15511 = n15464 ^ n15446;
  assign n15512 = n15455 ^ n15452;
  assign n15211 = n15210 ^ n15201;
  assign n15212 = n15189 ^ n15172;
  assign n15213 = n15186 ^ n15174;
  assign n15214 = n15183 ^ n15176;
  assign n15215 = n15177 ^ n12059;
  assign n15216 = n15180 ^ n15179;
  assign n15217 = ~n15215 & ~n15216;
  assign n15218 = n15214 & n15217;
  assign n15219 = n15213 & n15218;
  assign n15220 = n15212 & n15219;
  assign n15221 = n15192 ^ n15170;
  assign n15222 = ~n15220 & ~n15221;
  assign n15223 = n15195 ^ n15168;
  assign n15224 = ~n15222 & ~n15223;
  assign n15225 = n15198 ^ n15166;
  assign n15226 = ~n15224 & n15225;
  assign n15227 = n15211 & n15226;
  assign n15241 = n15240 ^ n15230;
  assign n15291 = n15227 & n15241;
  assign n15304 = n15303 ^ n15294;
  assign n15513 = ~n15291 & n15304;
  assign n15514 = ~n15512 & ~n15513;
  assign n15515 = n15458 ^ n15450;
  assign n15516 = ~n15514 & ~n15515;
  assign n15517 = n15461 ^ n15448;
  assign n15518 = ~n15516 & ~n15517;
  assign n15519 = ~n15511 & n15518;
  assign n15520 = n15510 & n15519;
  assign n15521 = n15470 ^ n15442;
  assign n15522 = n15520 & ~n15521;
  assign n15523 = n15473 ^ n15440;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = ~n15509 & n15524;
  assign n15526 = n15479 ^ n15436;
  assign n15527 = ~n15525 & n15526;
  assign n15528 = n15508 & n15527;
  assign n15529 = n15485 ^ n15432;
  assign n15530 = ~n15528 & n15529;
  assign n15531 = n15488 ^ n15430;
  assign n15532 = ~n15530 & ~n15531;
  assign n15533 = n15491 ^ n15428;
  assign n15534 = n15532 & n15533;
  assign n15535 = n15494 ^ n15426;
  assign n15536 = ~n15534 & ~n15535;
  assign n15537 = n15507 & ~n15536;
  assign n15657 = n15550 ^ n15537;
  assign n15567 = n15536 ^ n15507;
  assign n1302 = x423 ^ x231;
  assign n1303 = n1302 ^ n1202;
  assign n1304 = n1303 ^ x167;
  assign n15568 = n15567 ^ n1304;
  assign n15569 = n15535 ^ n15534;
  assign n15570 = n15569 ^ n1380;
  assign n15646 = n15533 ^ n15532;
  assign n15571 = n15531 ^ n15530;
  assign n15572 = n15571 ^ n955;
  assign n15638 = n15529 ^ n15528;
  assign n15573 = n15527 ^ n15508;
  assign n15574 = n15573 ^ n827;
  assign n15630 = n15526 ^ n15525;
  assign n15575 = n15524 ^ n15509;
  assign n15576 = n15575 ^ n731;
  assign n15577 = n15523 ^ n15522;
  assign n15578 = n15577 ^ n745;
  assign n15579 = n15521 ^ n15520;
  assign n15583 = n15582 ^ n15579;
  assign n15584 = n15519 ^ n15510;
  assign n15588 = n15587 ^ n15584;
  assign n15613 = n15518 ^ n15511;
  assign n15589 = n15517 ^ n15516;
  assign n15593 = n15592 ^ n15589;
  assign n15594 = n15515 ^ n15514;
  assign n15595 = n15594 ^ n594;
  assign n15596 = n15513 ^ n15512;
  assign n15600 = n15599 ^ n15596;
  assign n15305 = n15304 ^ n15291;
  assign n15242 = n15241 ^ n15227;
  assign n15243 = n15242 ^ n2070;
  assign n15283 = n15226 ^ n15211;
  assign n15244 = n15225 ^ n15224;
  assign n15245 = n15244 ^ n1917;
  assign n15246 = n15223 ^ n15222;
  assign n15247 = n15246 ^ n1801;
  assign n15272 = n15221 ^ n15220;
  assign n15248 = n15219 ^ n15212;
  assign n15249 = n15248 ^ n1783;
  assign n15250 = n15218 ^ n15213;
  assign n15251 = n15250 ^ n1448;
  assign n15252 = n15217 ^ n15214;
  assign n15256 = n15255 ^ n15252;
  assign n15257 = n1466 & n15215;
  assign n15258 = n15257 ^ n1415;
  assign n15259 = n15216 ^ n15215;
  assign n15260 = n15259 ^ n15257;
  assign n15261 = n15258 & ~n15260;
  assign n15262 = n15261 ^ n1415;
  assign n15263 = n15262 ^ n15252;
  assign n15264 = n15256 & ~n15263;
  assign n15265 = n15264 ^ n15255;
  assign n15266 = n15265 ^ n15250;
  assign n15267 = n15251 & ~n15266;
  assign n15268 = n15267 ^ n1448;
  assign n15269 = n15268 ^ n15248;
  assign n15270 = n15249 & ~n15269;
  assign n15271 = n15270 ^ n1783;
  assign n15273 = n15272 ^ n15271;
  assign n15274 = n15272 ^ n1789;
  assign n15275 = n15273 & ~n15274;
  assign n15276 = n15275 ^ n1789;
  assign n15277 = n15276 ^ n15246;
  assign n15278 = n15247 & ~n15277;
  assign n15279 = n15278 ^ n1801;
  assign n15280 = n15279 ^ n15244;
  assign n15281 = n15245 & ~n15280;
  assign n15282 = n15281 ^ n1917;
  assign n15284 = n15283 ^ n15282;
  assign n15285 = n15283 ^ n1927;
  assign n15286 = n15284 & ~n15285;
  assign n15287 = n15286 ^ n1927;
  assign n15288 = n15287 ^ n15242;
  assign n15289 = ~n15243 & n15288;
  assign n15290 = n15289 ^ n2070;
  assign n15306 = n15305 ^ n15290;
  assign n15601 = n15309 ^ n15305;
  assign n15602 = n15306 & ~n15601;
  assign n15603 = n15602 ^ n15309;
  assign n15604 = n15603 ^ n15596;
  assign n15605 = ~n15600 & n15604;
  assign n15606 = n15605 ^ n15599;
  assign n15607 = n15606 ^ n15594;
  assign n15608 = n15595 & ~n15607;
  assign n15609 = n15608 ^ n594;
  assign n15610 = n15609 ^ n15589;
  assign n15611 = ~n15593 & n15610;
  assign n15612 = n15611 ^ n15592;
  assign n15614 = n15613 ^ n15612;
  assign n15615 = n15613 ^ n518;
  assign n15616 = ~n15614 & n15615;
  assign n15617 = n15616 ^ n518;
  assign n15618 = n15617 ^ n15584;
  assign n15619 = ~n15588 & n15618;
  assign n15620 = n15619 ^ n15587;
  assign n15621 = n15620 ^ n15579;
  assign n15622 = n15583 & ~n15621;
  assign n15623 = n15622 ^ n15582;
  assign n15624 = n15623 ^ n15577;
  assign n15625 = n15578 & ~n15624;
  assign n15626 = n15625 ^ n745;
  assign n15627 = n15626 ^ n15575;
  assign n15628 = ~n15576 & n15627;
  assign n15629 = n15628 ^ n731;
  assign n15631 = n15630 ^ n15629;
  assign n15632 = n15630 ^ n737;
  assign n15633 = ~n15631 & n15632;
  assign n15634 = n15633 ^ n737;
  assign n15635 = n15634 ^ n15573;
  assign n15636 = ~n15574 & n15635;
  assign n15637 = n15636 ^ n827;
  assign n15639 = n15638 ^ n15637;
  assign n15640 = n15638 ^ n949;
  assign n15641 = n15639 & ~n15640;
  assign n15642 = n15641 ^ n949;
  assign n15643 = n15642 ^ n15571;
  assign n15644 = ~n15572 & n15643;
  assign n15645 = n15644 ^ n955;
  assign n15647 = n15646 ^ n15645;
  assign n15648 = n15646 ^ n1113;
  assign n15649 = n15647 & ~n15648;
  assign n15650 = n15649 ^ n1113;
  assign n15651 = n15650 ^ n15569;
  assign n15652 = n15570 & ~n15651;
  assign n15653 = n15652 ^ n1380;
  assign n15654 = n15653 ^ n15567;
  assign n15655 = n15568 & ~n15654;
  assign n15656 = n15655 ^ n1304;
  assign n15658 = n15657 ^ n15656;
  assign n2450 = n2376 ^ x230;
  assign n2451 = n2450 ^ x422;
  assign n2452 = n2451 ^ x166;
  assign n15659 = n15657 ^ n2452;
  assign n15660 = n15658 & ~n15659;
  assign n15661 = n15660 ^ n2452;
  assign n15559 = n15543 ^ n15542;
  assign n15560 = ~n15547 & n15559;
  assign n15561 = n15560 ^ n15542;
  assign n15558 = n15067 ^ n15039;
  assign n15562 = n15561 ^ n15558;
  assign n15556 = n13893 ^ n13194;
  assign n15557 = n15556 ^ n14429;
  assign n15563 = n15562 ^ n15557;
  assign n15552 = n15548 ^ n15540;
  assign n15553 = ~n15549 & n15552;
  assign n15554 = n15553 ^ n12600;
  assign n15555 = n15554 ^ n12617;
  assign n15564 = n15563 ^ n15555;
  assign n15551 = n15537 & n15550;
  assign n15565 = n15564 ^ n15551;
  assign n15566 = n15565 ^ n2437;
  assign n15707 = n15661 ^ n15566;
  assign n15864 = n15709 ^ n15707;
  assign n15865 = n13322 & ~n15864;
  assign n15866 = n15865 ^ n13380;
  assign n15673 = n15558 ^ n15557;
  assign n15674 = ~n15562 & n15673;
  assign n15675 = n15674 ^ n15557;
  assign n15672 = n15072 ^ n1105;
  assign n15676 = n15675 ^ n15672;
  assign n15670 = n13888 ^ n13235;
  assign n15671 = n15670 ^ n14453;
  assign n15677 = n15676 ^ n15671;
  assign n15678 = n15677 ^ n12598;
  assign n15666 = n15563 ^ n12617;
  assign n15667 = n15563 ^ n15554;
  assign n15668 = ~n15666 & n15667;
  assign n15669 = n15668 ^ n12617;
  assign n15679 = n15678 ^ n15669;
  assign n15665 = n15551 & n15564;
  assign n15680 = n15679 ^ n15665;
  assign n15662 = n15661 ^ n15565;
  assign n15663 = ~n15566 & n15662;
  assign n15664 = n15663 ^ n2437;
  assign n15681 = n15680 ^ n15664;
  assign n15712 = n15681 ^ n2445;
  assign n15710 = ~n15707 & n15709;
  assign n15705 = n14563 ^ n13416;
  assign n15706 = n15705 ^ n14831;
  assign n15711 = n15710 ^ n15706;
  assign n15867 = n15712 ^ n15711;
  assign n15868 = n15867 ^ n15865;
  assign n15869 = ~n15866 & ~n15868;
  assign n15870 = n15869 ^ n13380;
  assign n15713 = n15712 ^ n15706;
  assign n15714 = ~n15711 & ~n15713;
  assign n15715 = n15714 ^ n15710;
  assign n15702 = n14570 ^ n13410;
  assign n15703 = n15702 ^ n14830;
  assign n15694 = n13936 ^ n13273;
  assign n15695 = n15694 ^ n14478;
  assign n15692 = n15075 ^ n15037;
  assign n15689 = n15672 ^ n15671;
  assign n15690 = ~n15676 & ~n15689;
  assign n15691 = n15690 ^ n15671;
  assign n15693 = n15692 ^ n15691;
  assign n15696 = n15695 ^ n15693;
  assign n15697 = n15696 ^ n12590;
  assign n15686 = n15677 ^ n15669;
  assign n15687 = n15678 & ~n15686;
  assign n15688 = n15687 ^ n12598;
  assign n15698 = n15697 ^ n15688;
  assign n15685 = ~n15665 & n15679;
  assign n15699 = n15698 ^ n15685;
  assign n15700 = n15699 ^ n2551;
  assign n15682 = n15680 ^ n2445;
  assign n15683 = n15681 & ~n15682;
  assign n15684 = n15683 ^ n2445;
  assign n15701 = n15700 ^ n15684;
  assign n15704 = n15703 ^ n15701;
  assign n15862 = n15715 ^ n15704;
  assign n15863 = n15862 ^ n13436;
  assign n15934 = n15870 ^ n15863;
  assign n15935 = n15864 ^ n13322;
  assign n15936 = n15867 ^ n15866;
  assign n15937 = ~n15935 & ~n15936;
  assign n15938 = n15934 & n15937;
  assign n15871 = n15870 ^ n15862;
  assign n15872 = ~n15863 & n15871;
  assign n15873 = n15872 ^ n13436;
  assign n15740 = n15205 ^ n14236;
  assign n15741 = n15740 ^ n13404;
  assign n15735 = ~n15685 & ~n15698;
  assign n15731 = n13430 ^ n13295;
  assign n15732 = n15731 ^ n14505;
  assign n15727 = n15695 ^ n15692;
  assign n15728 = ~n15693 & ~n15727;
  assign n15729 = n15728 ^ n15695;
  assign n15726 = n15078 ^ n15035;
  assign n15730 = n15729 ^ n15726;
  assign n15733 = n15732 ^ n15730;
  assign n15722 = n15696 ^ n15688;
  assign n15723 = n15697 & n15722;
  assign n15724 = n15723 ^ n12590;
  assign n15725 = n15724 ^ n12066;
  assign n15734 = n15733 ^ n15725;
  assign n15736 = n15735 ^ n15734;
  assign n15719 = n15699 ^ n15684;
  assign n15720 = ~n15700 & n15719;
  assign n15721 = n15720 ^ n2551;
  assign n15737 = n15736 ^ n15721;
  assign n15738 = n15737 ^ n2546;
  assign n15716 = n15715 ^ n15701;
  assign n15717 = n15704 & n15716;
  assign n15718 = n15717 ^ n15703;
  assign n15739 = n15738 ^ n15718;
  assign n15860 = n15741 ^ n15739;
  assign n15861 = n15860 ^ n13431;
  assign n15933 = n15873 ^ n15861;
  assign n15989 = n15938 ^ n15933;
  assign n15990 = n15989 ^ n1599;
  assign n15991 = n15937 ^ n15934;
  assign n15992 = n15991 ^ n1482;
  assign n15996 = n15935 & n15995;
  assign n15997 = n15996 ^ n1493;
  assign n15998 = n15936 ^ n15935;
  assign n15999 = n15998 ^ n15996;
  assign n16000 = n15997 & ~n15999;
  assign n16001 = n16000 ^ n1493;
  assign n16002 = n16001 ^ n15991;
  assign n16003 = n15992 & ~n16002;
  assign n16004 = n16003 ^ n1482;
  assign n16005 = n16004 ^ n15989;
  assign n16006 = ~n15990 & n16005;
  assign n16007 = n16006 ^ n1599;
  assign n15939 = ~n15933 & n15938;
  assign n15874 = n15873 ^ n15860;
  assign n15875 = n15861 & n15874;
  assign n15876 = n15875 ^ n13431;
  assign n15764 = ~n15734 & n15735;
  assign n15761 = n15083 ^ n2294;
  assign n15758 = n13424 ^ n13310;
  assign n15759 = n15758 ^ n14536;
  assign n15755 = n15732 ^ n15726;
  assign n15756 = ~n15730 & ~n15755;
  assign n15757 = n15756 ^ n15732;
  assign n15760 = n15759 ^ n15757;
  assign n15762 = n15761 ^ n15760;
  assign n15750 = n15733 ^ n12066;
  assign n15751 = n15733 ^ n15724;
  assign n15752 = ~n15750 & n15751;
  assign n15753 = n15752 ^ n12066;
  assign n15754 = n15753 ^ n12630;
  assign n15763 = n15762 ^ n15754;
  assign n15765 = n15764 ^ n15763;
  assign n15746 = n15736 ^ n2546;
  assign n15747 = ~n15737 & n15746;
  assign n15748 = n15747 ^ n2546;
  assign n15749 = n15748 ^ n1499;
  assign n15766 = n15765 ^ n15749;
  assign n15328 = n14580 ^ n13398;
  assign n15329 = n15328 ^ n15237;
  assign n15857 = n15766 ^ n15329;
  assign n15742 = n15741 ^ n15718;
  assign n15743 = n15739 & n15742;
  assign n15744 = n15743 ^ n15741;
  assign n15858 = n15857 ^ n15744;
  assign n15859 = n15858 ^ n13425;
  assign n15932 = n15876 ^ n15859;
  assign n15987 = n15939 ^ n15932;
  assign n15988 = n15987 ^ n1628;
  assign n16158 = n16007 ^ n15988;
  assign n15316 = n15268 ^ n15249;
  assign n17613 = n16158 ^ n15316;
  assign n15770 = n15215 ^ n1466;
  assign n16419 = n15770 ^ n14830;
  assign n16420 = n16419 ^ n14556;
  assign n16089 = n15614 ^ n518;
  assign n16069 = n15609 ^ n15593;
  assign n16067 = n14897 ^ n14334;
  assign n16068 = n16067 ^ n15414;
  assign n16070 = n16069 ^ n16068;
  assign n15831 = n15603 ^ n15600;
  assign n15318 = n14711 ^ n14051;
  assign n15320 = n15319 ^ n15318;
  assign n15317 = n15265 ^ n15251;
  assign n15321 = n15320 ^ n15317;
  assign n15324 = n14658 ^ n13386;
  assign n15326 = n15325 ^ n15324;
  assign n15323 = n15259 ^ n15258;
  assign n15327 = n15326 ^ n15323;
  assign n15745 = n15744 ^ n15329;
  assign n15767 = n15766 ^ n15744;
  assign n15768 = n15745 & n15767;
  assign n15769 = n15768 ^ n15329;
  assign n15771 = n15770 ^ n15769;
  assign n15772 = n14589 ^ n13392;
  assign n15773 = n15772 ^ n15300;
  assign n15774 = n15773 ^ n15770;
  assign n15775 = n15771 & n15774;
  assign n15776 = n15775 ^ n15773;
  assign n15777 = n15776 ^ n15323;
  assign n15778 = n15327 & ~n15777;
  assign n15779 = n15778 ^ n15326;
  assign n15322 = n15262 ^ n15256;
  assign n15780 = n15779 ^ n15322;
  assign n15781 = n14697 ^ n13967;
  assign n15782 = n15781 ^ n15353;
  assign n15783 = n15782 ^ n15322;
  assign n15784 = ~n15780 & ~n15783;
  assign n15785 = n15784 ^ n15782;
  assign n15786 = n15785 ^ n15317;
  assign n15787 = n15321 & n15786;
  assign n15788 = n15787 ^ n15320;
  assign n15789 = n15788 ^ n15316;
  assign n15790 = n14818 ^ n14183;
  assign n15791 = n15790 ^ n15349;
  assign n15792 = n15791 ^ n15316;
  assign n15793 = ~n15789 & n15792;
  assign n15794 = n15793 ^ n15791;
  assign n15315 = n15273 ^ n1789;
  assign n15795 = n15794 ^ n15315;
  assign n15796 = n14858 ^ n14202;
  assign n15797 = n15796 ^ n15378;
  assign n15798 = n15797 ^ n15315;
  assign n15799 = n15795 & n15798;
  assign n15800 = n15799 ^ n15797;
  assign n15314 = n15276 ^ n15247;
  assign n15801 = n15800 ^ n15314;
  assign n15802 = n14866 ^ n14227;
  assign n15803 = n15802 ^ n15347;
  assign n15804 = n15803 ^ n15314;
  assign n15805 = n15801 & n15804;
  assign n15806 = n15805 ^ n15803;
  assign n15313 = n15279 ^ n15245;
  assign n15807 = n15806 ^ n15313;
  assign n15808 = n14852 ^ n14256;
  assign n15809 = n15808 ^ n15341;
  assign n15810 = n15809 ^ n15313;
  assign n15811 = ~n15807 & ~n15810;
  assign n15812 = n15811 ^ n15809;
  assign n15312 = n15284 ^ n1927;
  assign n15813 = n15812 ^ n15312;
  assign n15814 = n14850 ^ n14254;
  assign n15815 = n15814 ^ n15391;
  assign n15816 = n15815 ^ n15312;
  assign n15817 = ~n15813 & n15816;
  assign n15818 = n15817 ^ n15815;
  assign n15311 = n15287 ^ n15243;
  assign n15819 = n15818 ^ n15311;
  assign n15820 = n14846 ^ n14246;
  assign n15821 = n15820 ^ n15337;
  assign n15822 = n15821 ^ n15311;
  assign n15823 = ~n15819 & ~n15822;
  assign n15824 = n15823 ^ n15821;
  assign n15310 = n15309 ^ n15306;
  assign n15825 = n15824 ^ n15310;
  assign n15826 = n15401 ^ n14842;
  assign n15827 = n15826 ^ n14245;
  assign n15828 = n15827 ^ n15310;
  assign n15829 = n15825 & n15828;
  assign n15830 = n15829 ^ n15827;
  assign n15832 = n15831 ^ n15830;
  assign n14235 = n14234 ^ n14233;
  assign n14827 = n14826 ^ n14235;
  assign n15919 = n15831 ^ n14827;
  assign n15920 = ~n15832 & n15919;
  assign n15921 = n15920 ^ n14827;
  assign n15918 = n15606 ^ n15595;
  assign n15922 = n15921 ^ n15918;
  assign n15916 = n14839 ^ n14288;
  assign n15917 = n15916 ^ n15330;
  assign n16064 = n15918 ^ n15917;
  assign n16065 = n15922 & n16064;
  assign n16066 = n16065 ^ n15917;
  assign n16086 = n16069 ^ n16066;
  assign n16087 = ~n16070 & n16086;
  assign n16088 = n16087 ^ n16068;
  assign n16090 = n16089 ^ n16088;
  assign n16084 = n14904 ^ n14401;
  assign n16085 = n16084 ^ n15423;
  assign n16091 = n16090 ^ n16085;
  assign n16071 = n16070 ^ n16066;
  assign n15923 = n15922 ^ n15917;
  assign n15924 = n15923 ^ n13456;
  assign n15833 = n15832 ^ n14827;
  assign n15834 = n15833 ^ n13461;
  assign n15835 = n15827 ^ n15825;
  assign n15836 = n15835 ^ n13466;
  assign n15837 = n15821 ^ n15819;
  assign n15838 = n15837 ^ n13471;
  assign n15839 = n15815 ^ n15813;
  assign n15840 = n15839 ^ n13476;
  assign n15841 = n15809 ^ n15807;
  assign n15842 = n15841 ^ n13481;
  assign n15843 = n15803 ^ n15801;
  assign n15844 = n15843 ^ n12845;
  assign n15845 = n15797 ^ n15795;
  assign n15846 = n15845 ^ n13388;
  assign n15847 = n15791 ^ n15789;
  assign n15848 = n15847 ^ n13394;
  assign n15849 = n15785 ^ n15321;
  assign n15850 = n15849 ^ n13400;
  assign n15851 = n15782 ^ n15780;
  assign n15852 = n15851 ^ n13406;
  assign n15853 = n15776 ^ n15327;
  assign n15854 = n15853 ^ n13412;
  assign n15855 = n15773 ^ n15771;
  assign n15856 = n15855 ^ n13419;
  assign n15877 = n15876 ^ n15858;
  assign n15878 = n15859 & ~n15877;
  assign n15879 = n15878 ^ n13425;
  assign n15880 = n15879 ^ n15855;
  assign n15881 = ~n15856 & n15880;
  assign n15882 = n15881 ^ n13419;
  assign n15883 = n15882 ^ n15853;
  assign n15884 = n15854 & ~n15883;
  assign n15885 = n15884 ^ n13412;
  assign n15886 = n15885 ^ n15851;
  assign n15887 = n15852 & n15886;
  assign n15888 = n15887 ^ n13406;
  assign n15889 = n15888 ^ n15849;
  assign n15890 = ~n15850 & ~n15889;
  assign n15891 = n15890 ^ n13400;
  assign n15892 = n15891 ^ n15847;
  assign n15893 = n15848 & ~n15892;
  assign n15894 = n15893 ^ n13394;
  assign n15895 = n15894 ^ n15845;
  assign n15896 = n15846 & ~n15895;
  assign n15897 = n15896 ^ n13388;
  assign n15898 = n15897 ^ n15843;
  assign n15899 = ~n15844 & n15898;
  assign n15900 = n15899 ^ n12845;
  assign n15901 = n15900 ^ n15841;
  assign n15902 = ~n15842 & n15901;
  assign n15903 = n15902 ^ n13481;
  assign n15904 = n15903 ^ n15839;
  assign n15905 = ~n15840 & n15904;
  assign n15906 = n15905 ^ n13476;
  assign n15907 = n15906 ^ n15837;
  assign n15908 = ~n15838 & ~n15907;
  assign n15909 = n15908 ^ n13471;
  assign n15910 = n15909 ^ n15835;
  assign n15911 = n15836 & n15910;
  assign n15912 = n15911 ^ n13466;
  assign n15913 = n15912 ^ n15833;
  assign n15914 = ~n15834 & n15913;
  assign n15915 = n15914 ^ n13461;
  assign n16061 = n15923 ^ n15915;
  assign n16062 = n15924 & n16061;
  assign n16063 = n16062 ^ n13456;
  assign n16072 = n16071 ^ n16063;
  assign n16081 = n16071 ^ n13451;
  assign n16082 = ~n16072 & ~n16081;
  assign n16083 = n16082 ^ n13451;
  assign n16092 = n16091 ^ n16083;
  assign n16269 = n16091 ^ n13446;
  assign n16270 = n16092 & n16269;
  assign n16271 = n16270 ^ n13446;
  assign n16213 = n14838 ^ n14422;
  assign n16214 = n16213 ^ n15501;
  assign n16209 = n16089 ^ n16085;
  assign n16210 = ~n16090 & ~n16209;
  assign n16211 = n16210 ^ n16085;
  assign n16138 = n15617 ^ n15588;
  assign n16212 = n16211 ^ n16138;
  assign n16267 = n16214 ^ n16212;
  assign n16268 = n16267 ^ n13585;
  assign n16317 = n16271 ^ n16268;
  assign n16073 = n16072 ^ n13451;
  assign n15925 = n15924 ^ n15915;
  assign n15926 = n15909 ^ n13466;
  assign n15927 = n15926 ^ n15835;
  assign n15928 = n15903 ^ n15840;
  assign n15929 = n15891 ^ n15848;
  assign n15930 = n15888 ^ n15850;
  assign n15931 = n15885 ^ n15852;
  assign n15940 = n15932 & n15939;
  assign n15941 = n15879 ^ n15856;
  assign n15942 = ~n15940 & n15941;
  assign n15943 = n15882 ^ n15854;
  assign n15944 = ~n15942 & n15943;
  assign n15945 = ~n15931 & ~n15944;
  assign n15946 = ~n15930 & n15945;
  assign n15947 = ~n15929 & n15946;
  assign n15948 = n15894 ^ n15846;
  assign n15949 = ~n15947 & n15948;
  assign n15950 = n15897 ^ n15844;
  assign n15951 = ~n15949 & n15950;
  assign n15952 = n15900 ^ n15842;
  assign n15953 = ~n15951 & ~n15952;
  assign n15954 = n15928 & ~n15953;
  assign n15955 = n15906 ^ n15838;
  assign n15956 = n15954 & n15955;
  assign n15957 = n15927 & n15956;
  assign n15958 = n15912 ^ n15834;
  assign n15959 = n15957 & n15958;
  assign n16074 = n15925 & ~n15959;
  assign n16080 = n16073 & n16074;
  assign n16093 = n16092 ^ n13446;
  assign n16318 = ~n16080 & ~n16093;
  assign n16319 = ~n16317 & n16318;
  assign n16272 = n16271 ^ n16267;
  assign n16273 = ~n16268 & n16272;
  assign n16274 = n16273 ^ n13585;
  assign n16215 = n16214 ^ n16138;
  assign n16216 = ~n16212 & ~n16215;
  assign n16217 = n16216 ^ n16214;
  assign n16206 = n14917 ^ n14446;
  assign n16207 = n16206 ^ n15543;
  assign n16133 = n15620 ^ n15583;
  assign n16208 = n16207 ^ n16133;
  assign n16265 = n16217 ^ n16208;
  assign n16266 = n16265 ^ n13695;
  assign n16320 = n16274 ^ n16266;
  assign n16321 = ~n16319 & n16320;
  assign n16275 = n16274 ^ n16265;
  assign n16276 = ~n16266 & n16275;
  assign n16277 = n16276 ^ n13695;
  assign n16218 = n16217 ^ n16207;
  assign n16219 = n16208 & ~n16218;
  assign n16220 = n16219 ^ n16133;
  assign n16203 = n14988 ^ n14467;
  assign n16204 = n16203 ^ n15558;
  assign n16129 = n15623 ^ n15578;
  assign n16205 = n16204 ^ n16129;
  assign n16263 = n16220 ^ n16205;
  assign n16264 = n16263 ^ n13749;
  assign n16322 = n16277 ^ n16264;
  assign n16323 = ~n16321 & n16322;
  assign n16278 = n16277 ^ n16263;
  assign n16279 = n16264 & ~n16278;
  assign n16280 = n16279 ^ n13749;
  assign n16221 = n16220 ^ n16204;
  assign n16222 = ~n16205 & n16221;
  assign n16223 = n16222 ^ n16129;
  assign n16200 = n15026 ^ n14498;
  assign n16201 = n16200 ^ n15672;
  assign n16124 = n15626 ^ n15576;
  assign n16202 = n16201 ^ n16124;
  assign n16261 = n16223 ^ n16202;
  assign n16262 = n16261 ^ n13881;
  assign n16324 = n16280 ^ n16262;
  assign n16325 = n16323 & ~n16324;
  assign n16228 = n15111 ^ n14531;
  assign n16229 = n16228 ^ n15692;
  assign n16224 = n16223 ^ n16124;
  assign n16225 = n16202 & n16224;
  assign n16226 = n16225 ^ n16201;
  assign n16119 = n15631 ^ n737;
  assign n16227 = n16226 ^ n16119;
  assign n16284 = n16229 ^ n16227;
  assign n16281 = n16280 ^ n16261;
  assign n16282 = ~n16262 & n16281;
  assign n16283 = n16282 ^ n13881;
  assign n16285 = n16284 ^ n16283;
  assign n16326 = n16285 ^ n13930;
  assign n16327 = ~n16325 & n16326;
  assign n16286 = n16284 ^ n13930;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = n16287 ^ n13930;
  assign n16328 = n16288 ^ n13162;
  assign n16230 = n16229 ^ n16119;
  assign n16231 = n16227 & n16230;
  assign n16232 = n16231 ^ n16229;
  assign n16197 = n14429 ^ n13903;
  assign n16198 = n16197 ^ n15726;
  assign n16114 = n15634 ^ n15574;
  assign n16199 = n16198 ^ n16114;
  assign n16259 = n16232 ^ n16199;
  assign n16329 = n16328 ^ n16259;
  assign n16330 = ~n16327 & n16329;
  assign n16233 = n16232 ^ n16114;
  assign n16234 = n16199 & n16233;
  assign n16235 = n16234 ^ n16198;
  assign n16194 = n14453 ^ n13898;
  assign n16195 = n16194 ^ n15761;
  assign n16292 = n16235 ^ n16195;
  assign n16109 = n15639 ^ n949;
  assign n16293 = n16292 ^ n16109;
  assign n16260 = n16259 ^ n13162;
  assign n16289 = n16288 ^ n16259;
  assign n16290 = ~n16260 & ~n16289;
  assign n16291 = n16290 ^ n13162;
  assign n16294 = n16293 ^ n16291;
  assign n16316 = n16294 ^ n13160;
  assign n16347 = n16330 ^ n16316;
  assign n16348 = n16347 ^ n2281;
  assign n16349 = n16329 ^ n16327;
  assign n2269 = n1309 ^ x263;
  assign n2270 = n2269 ^ x455;
  assign n2271 = n2270 ^ x199;
  assign n16350 = n16349 ^ n2271;
  assign n16351 = n16326 ^ n16325;
  assign n16352 = n16351 ^ n1223;
  assign n16353 = n16324 ^ n16323;
  assign n1053 = n975 ^ x265;
  assign n1054 = n1053 ^ x457;
  assign n1055 = n1054 ^ x201;
  assign n16354 = n16353 ^ n1055;
  assign n16356 = n16320 ^ n16319;
  assign n16357 = n16356 ^ n918;
  assign n16358 = n16318 ^ n16317;
  assign n16359 = n16358 ^ n912;
  assign n16094 = n16093 ^ n16080;
  assign n16095 = n16094 ^ n926;
  assign n16075 = n16074 ^ n16073;
  assign n15960 = n15959 ^ n15925;
  assign n15964 = n15963 ^ n15960;
  assign n15965 = n15958 ^ n15957;
  assign n15966 = n15965 ^ n537;
  assign n15967 = n15956 ^ n15927;
  assign n15968 = n15967 ^ n625;
  assign n15969 = n15955 ^ n15954;
  assign n15970 = n15969 ^ n619;
  assign n15971 = n15953 ^ n15928;
  assign n15975 = n15974 ^ n15971;
  assign n16038 = n15952 ^ n15951;
  assign n15976 = n15950 ^ n15949;
  assign n15980 = n15979 ^ n15976;
  assign n16030 = n15948 ^ n15947;
  assign n15981 = n15946 ^ n15929;
  assign n15982 = n15981 ^ n2063;
  assign n16022 = n15945 ^ n15930;
  assign n15983 = n15944 ^ n15931;
  assign n15984 = n15983 ^ n1823;
  assign n15985 = n15943 ^ n15942;
  assign n15986 = n15985 ^ n2029;
  assign n16011 = n15941 ^ n15940;
  assign n16008 = n16007 ^ n15987;
  assign n16009 = n15988 & ~n16008;
  assign n16010 = n16009 ^ n1628;
  assign n16012 = n16011 ^ n16010;
  assign n16013 = n16011 ^ n1688;
  assign n16014 = ~n16012 & n16013;
  assign n16015 = n16014 ^ n1688;
  assign n16016 = n16015 ^ n15985;
  assign n16017 = ~n15986 & n16016;
  assign n16018 = n16017 ^ n2029;
  assign n16019 = n16018 ^ n15983;
  assign n16020 = ~n15984 & n16019;
  assign n16021 = n16020 ^ n1823;
  assign n16023 = n16022 ^ n16021;
  assign n16024 = n16022 ^ n2045;
  assign n16025 = ~n16023 & n16024;
  assign n16026 = n16025 ^ n2045;
  assign n16027 = n16026 ^ n15981;
  assign n16028 = n15982 & ~n16027;
  assign n16029 = n16028 ^ n2063;
  assign n16031 = n16030 ^ n16029;
  assign n16032 = n16030 ^ n2206;
  assign n16033 = n16031 & ~n16032;
  assign n16034 = n16033 ^ n2206;
  assign n16035 = n16034 ^ n15976;
  assign n16036 = n15980 & ~n16035;
  assign n16037 = n16036 ^ n15979;
  assign n16039 = n16038 ^ n16037;
  assign n16043 = n16042 ^ n16038;
  assign n16044 = ~n16039 & n16043;
  assign n16045 = n16044 ^ n16042;
  assign n16046 = n16045 ^ n15971;
  assign n16047 = n15975 & ~n16046;
  assign n16048 = n16047 ^ n15974;
  assign n16049 = n16048 ^ n15969;
  assign n16050 = ~n15970 & n16049;
  assign n16051 = n16050 ^ n619;
  assign n16052 = n16051 ^ n15967;
  assign n16053 = ~n15968 & n16052;
  assign n16054 = n16053 ^ n625;
  assign n16055 = n16054 ^ n537;
  assign n16056 = ~n15966 & ~n16055;
  assign n16057 = n16056 ^ n15965;
  assign n16058 = n16057 ^ n15963;
  assign n16059 = ~n15964 & n16058;
  assign n16060 = n16059 ^ n15960;
  assign n16076 = n16075 ^ n16060;
  assign n16077 = n16075 ^ n557;
  assign n16078 = n16076 & n16077;
  assign n16079 = n16078 ^ n557;
  assign n16360 = n16094 ^ n16079;
  assign n16361 = ~n16095 & n16360;
  assign n16362 = n16361 ^ n926;
  assign n16363 = n16362 ^ n16358;
  assign n16364 = n16359 & ~n16363;
  assign n16365 = n16364 ^ n912;
  assign n16366 = n16365 ^ n16356;
  assign n16367 = ~n16357 & n16366;
  assign n16368 = n16367 ^ n918;
  assign n16355 = n16322 ^ n16321;
  assign n16369 = n16368 ^ n16355;
  assign n16370 = n16355 ^ n1049;
  assign n16371 = ~n16369 & n16370;
  assign n16372 = n16371 ^ n1049;
  assign n16373 = n16372 ^ n16353;
  assign n16374 = n16354 & ~n16373;
  assign n16375 = n16374 ^ n1055;
  assign n16376 = n16375 ^ n16351;
  assign n16377 = ~n16352 & n16376;
  assign n16378 = n16377 ^ n1223;
  assign n16379 = n16378 ^ n16349;
  assign n16380 = n16350 & ~n16379;
  assign n16381 = n16380 ^ n2271;
  assign n16382 = n16381 ^ n16347;
  assign n16383 = n16348 & ~n16382;
  assign n16384 = n16383 ^ n2281;
  assign n2349 = n2309 ^ x261;
  assign n2350 = n2349 ^ x453;
  assign n2351 = n2350 ^ x197;
  assign n16417 = n16384 ^ n2351;
  assign n16331 = ~n16316 & n16330;
  assign n16295 = n16293 ^ n13160;
  assign n16296 = ~n16294 & ~n16295;
  assign n16297 = n16296 ^ n13160;
  assign n16314 = n16297 ^ n13194;
  assign n16196 = n16195 ^ n16109;
  assign n16236 = n16235 ^ n16109;
  assign n16237 = n16196 & ~n16236;
  assign n16238 = n16237 ^ n16195;
  assign n16191 = n14478 ^ n13893;
  assign n16192 = n16191 ^ n15128;
  assign n16256 = n16238 ^ n16192;
  assign n16104 = n15642 ^ n15572;
  assign n16257 = n16256 ^ n16104;
  assign n16315 = n16314 ^ n16257;
  assign n16345 = n16331 ^ n16315;
  assign n16418 = n16417 ^ n16345;
  assign n16563 = n16420 ^ n16418;
  assign n16692 = n16563 ^ n13418;
  assign n16346 = n16345 ^ n2351;
  assign n16385 = n16384 ^ n16345;
  assign n16386 = n16346 & ~n16385;
  assign n16387 = n16386 ^ n2351;
  assign n16332 = ~n16315 & n16331;
  assign n16258 = n16257 ^ n13194;
  assign n16298 = n16297 ^ n16257;
  assign n16299 = n16258 & ~n16298;
  assign n16300 = n16299 ^ n13194;
  assign n16193 = n16192 ^ n16104;
  assign n16239 = n16238 ^ n16104;
  assign n16240 = ~n16193 & ~n16239;
  assign n16241 = n16240 ^ n16192;
  assign n16188 = n14505 ^ n13888;
  assign n16189 = n16188 ^ n15133;
  assign n16253 = n16241 ^ n16189;
  assign n16099 = n15647 ^ n1113;
  assign n16254 = n16253 ^ n16099;
  assign n16255 = n16254 ^ n13235;
  assign n16313 = n16300 ^ n16255;
  assign n16343 = n16332 ^ n16313;
  assign n1539 = n1538 ^ x260;
  assign n1540 = n1539 ^ x452;
  assign n1541 = n1540 ^ x196;
  assign n16344 = n16343 ^ n1541;
  assign n16423 = n16387 ^ n16344;
  assign n16421 = n16418 & n16420;
  assign n16415 = n15205 ^ n14563;
  assign n16416 = n16415 ^ n15323;
  assign n16422 = n16421 ^ n16416;
  assign n16566 = n16423 ^ n16422;
  assign n16564 = ~n13418 & n16563;
  assign n16565 = n16564 ^ n13416;
  assign n16693 = n16566 ^ n16565;
  assign n16694 = ~n16692 & n16693;
  assign n16567 = n16566 ^ n16564;
  assign n16568 = n16565 & ~n16567;
  assign n16569 = n16568 ^ n13416;
  assign n16388 = n16387 ^ n1541;
  assign n16389 = n16344 & ~n16388;
  assign n16390 = n16389 ^ n16343;
  assign n16333 = ~n16313 & ~n16332;
  assign n16190 = n16189 ^ n16099;
  assign n16242 = n16241 ^ n16099;
  assign n16243 = n16190 & n16242;
  assign n16244 = n16243 ^ n16189;
  assign n16185 = n14536 ^ n13936;
  assign n16186 = n16185 ^ n15137;
  assign n16184 = n15650 ^ n15570;
  assign n16187 = n16186 ^ n16184;
  assign n16304 = n16244 ^ n16187;
  assign n16301 = n16300 ^ n16254;
  assign n16302 = ~n16255 & ~n16301;
  assign n16303 = n16302 ^ n13235;
  assign n16305 = n16304 ^ n16303;
  assign n16312 = n16305 ^ n13273;
  assign n16341 = n16333 ^ n16312;
  assign n16342 = n16341 ^ n2489;
  assign n16430 = n16390 ^ n16342;
  assign n16427 = n15322 ^ n15237;
  assign n16428 = n16427 ^ n14570;
  assign n16560 = n16430 ^ n16428;
  assign n16424 = n16423 ^ n16416;
  assign n16425 = n16422 & ~n16424;
  assign n16426 = n16425 ^ n16421;
  assign n16561 = n16560 ^ n16426;
  assign n16562 = n16561 ^ n13410;
  assign n16691 = n16569 ^ n16562;
  assign n16799 = n16694 ^ n16691;
  assign n16786 = n1430 & n16692;
  assign n16790 = n16789 ^ n16786;
  assign n16791 = n16693 ^ n16692;
  assign n16792 = n16791 ^ n16786;
  assign n16793 = n16790 & n16792;
  assign n16794 = n16793 ^ n16789;
  assign n16798 = n16797 ^ n16794;
  assign n17021 = n16799 ^ n16798;
  assign n17614 = n17613 ^ n17021;
  assign n16654 = n16365 ^ n918;
  assign n16655 = n16654 ^ n16356;
  assign n16970 = n16655 ^ n15672;
  assign n16971 = n16970 ^ n16099;
  assign n16152 = n16018 ^ n15984;
  assign n16150 = n15337 ^ n14852;
  assign n16151 = n16150 ^ n15918;
  assign n16153 = n16152 ^ n16151;
  assign n16458 = n16015 ^ n15986;
  assign n16155 = n15341 ^ n14858;
  assign n16156 = n16155 ^ n15310;
  assign n16154 = n16012 ^ n1688;
  assign n16157 = n16156 ^ n16154;
  assign n16159 = n15347 ^ n14818;
  assign n16160 = n16159 ^ n15311;
  assign n16161 = n16160 ^ n16158;
  assign n16163 = n15378 ^ n14711;
  assign n16164 = n16163 ^ n15312;
  assign n16162 = n16004 ^ n15990;
  assign n16165 = n16164 ^ n16162;
  assign n16167 = n15349 ^ n14697;
  assign n16168 = n16167 ^ n15313;
  assign n16166 = n16001 ^ n15992;
  assign n16169 = n16168 ^ n16166;
  assign n16171 = n15319 ^ n14658;
  assign n16172 = n16171 ^ n15314;
  assign n16170 = n15998 ^ n15997;
  assign n16173 = n16172 ^ n16170;
  assign n16175 = n15353 ^ n14589;
  assign n16176 = n16175 ^ n15315;
  assign n16174 = n15995 ^ n15935;
  assign n16177 = n16176 ^ n16174;
  assign n16334 = n16312 & ~n16333;
  assign n16306 = n16304 ^ n13273;
  assign n16307 = ~n16305 & n16306;
  assign n16308 = n16307 ^ n13273;
  assign n16245 = n16244 ^ n16184;
  assign n16246 = n16187 & n16245;
  assign n16247 = n16246 ^ n16186;
  assign n16181 = n15145 ^ n13430;
  assign n16182 = n16181 ^ n14240;
  assign n16180 = n15653 ^ n15568;
  assign n16183 = n16182 ^ n16180;
  assign n16251 = n16247 ^ n16183;
  assign n16252 = n16251 ^ n13295;
  assign n16335 = n16308 ^ n16252;
  assign n16398 = n16334 & ~n16335;
  assign n16402 = n16401 ^ n16398;
  assign n16403 = n16402 ^ n15758;
  assign n16404 = n16403 ^ n15122;
  assign n16405 = n16404 ^ n14549;
  assign n16397 = n15658 ^ n2452;
  assign n16406 = n16405 ^ n16397;
  assign n16336 = n16335 ^ n16334;
  assign n16340 = n16339 ^ n16336;
  assign n16391 = n16390 ^ n16341;
  assign n16392 = n16342 & ~n16391;
  assign n16393 = n16392 ^ n2489;
  assign n16394 = n16393 ^ n16336;
  assign n16395 = n16340 & ~n16394;
  assign n16396 = n16395 ^ n16339;
  assign n16407 = n16406 ^ n16396;
  assign n16309 = n16308 ^ n16251;
  assign n16310 = ~n16252 & ~n16309;
  assign n16311 = n16310 ^ n13295;
  assign n16408 = n16407 ^ n16311;
  assign n16248 = n16247 ^ n16180;
  assign n16249 = ~n16183 & ~n16248;
  assign n16250 = n16249 ^ n16182;
  assign n16409 = n16408 ^ n16250;
  assign n16178 = n15325 ^ n14580;
  assign n16179 = n16178 ^ n15316;
  assign n16410 = n16409 ^ n16179;
  assign n16413 = n16393 ^ n16340;
  assign n16411 = n15300 ^ n14236;
  assign n16412 = n16411 ^ n15317;
  assign n16414 = n16413 ^ n16412;
  assign n16429 = n16428 ^ n16426;
  assign n16431 = n16430 ^ n16426;
  assign n16432 = n16429 & ~n16431;
  assign n16433 = n16432 ^ n16428;
  assign n16434 = n16433 ^ n16413;
  assign n16435 = ~n16414 & ~n16434;
  assign n16436 = n16435 ^ n16412;
  assign n16437 = n16436 ^ n16179;
  assign n16438 = n16410 & n16437;
  assign n16439 = n16438 ^ n16409;
  assign n16440 = n16439 ^ n16174;
  assign n16441 = ~n16177 & ~n16440;
  assign n16442 = n16441 ^ n16176;
  assign n16443 = n16442 ^ n16170;
  assign n16444 = ~n16173 & n16443;
  assign n16445 = n16444 ^ n16172;
  assign n16446 = n16445 ^ n16166;
  assign n16447 = n16169 & n16446;
  assign n16448 = n16447 ^ n16168;
  assign n16449 = n16448 ^ n16162;
  assign n16450 = ~n16165 & n16449;
  assign n16451 = n16450 ^ n16164;
  assign n16452 = n16451 ^ n16158;
  assign n16453 = n16161 & ~n16452;
  assign n16454 = n16453 ^ n16160;
  assign n16455 = n16454 ^ n16154;
  assign n16456 = ~n16157 & ~n16455;
  assign n16457 = n16456 ^ n16156;
  assign n16459 = n16458 ^ n16457;
  assign n16460 = n15391 ^ n14866;
  assign n16461 = n16460 ^ n15831;
  assign n16462 = n16461 ^ n16458;
  assign n16463 = ~n16459 & n16462;
  assign n16464 = n16463 ^ n16461;
  assign n16465 = n16464 ^ n16152;
  assign n16466 = ~n16153 & ~n16465;
  assign n16467 = n16466 ^ n16151;
  assign n16148 = n16023 ^ n2045;
  assign n16146 = n15401 ^ n14850;
  assign n16147 = n16146 ^ n16069;
  assign n16149 = n16148 ^ n16147;
  assign n16539 = n16467 ^ n16149;
  assign n16540 = n16539 ^ n14254;
  assign n16541 = n16464 ^ n16153;
  assign n16542 = n16541 ^ n14256;
  assign n16543 = n16461 ^ n16459;
  assign n16544 = n16543 ^ n14227;
  assign n16596 = n16454 ^ n16156;
  assign n16597 = n16596 ^ n16154;
  assign n16545 = n16451 ^ n16161;
  assign n16546 = n16545 ^ n14183;
  assign n16547 = n16448 ^ n16165;
  assign n16548 = n16547 ^ n14051;
  assign n16549 = n16445 ^ n16168;
  assign n16550 = n16549 ^ n16166;
  assign n16551 = n16550 ^ n13967;
  assign n16552 = n16442 ^ n16172;
  assign n16553 = n16552 ^ n16170;
  assign n16554 = n16553 ^ n13386;
  assign n16555 = n16439 ^ n16177;
  assign n16556 = n16555 ^ n13392;
  assign n16576 = n16436 ^ n16410;
  assign n16557 = n16433 ^ n16412;
  assign n16558 = n16557 ^ n16413;
  assign n16559 = n16558 ^ n13404;
  assign n16570 = n16569 ^ n16561;
  assign n16571 = ~n16562 & ~n16570;
  assign n16572 = n16571 ^ n13410;
  assign n16573 = n16572 ^ n16558;
  assign n16574 = n16559 & ~n16573;
  assign n16575 = n16574 ^ n13404;
  assign n16577 = n16576 ^ n16575;
  assign n16578 = n16576 ^ n13398;
  assign n16579 = ~n16577 & n16578;
  assign n16580 = n16579 ^ n13398;
  assign n16581 = n16580 ^ n16555;
  assign n16582 = ~n16556 & ~n16581;
  assign n16583 = n16582 ^ n13392;
  assign n16584 = n16583 ^ n16553;
  assign n16585 = n16554 & ~n16584;
  assign n16586 = n16585 ^ n13386;
  assign n16587 = n16586 ^ n16550;
  assign n16588 = n16551 & n16587;
  assign n16589 = n16588 ^ n13967;
  assign n16590 = n16589 ^ n16547;
  assign n16591 = n16548 & ~n16590;
  assign n16592 = n16591 ^ n14051;
  assign n16593 = n16592 ^ n16545;
  assign n16594 = n16546 & n16593;
  assign n16595 = n16594 ^ n14183;
  assign n16598 = n16597 ^ n16595;
  assign n16599 = n16597 ^ n14202;
  assign n16600 = n16598 & ~n16599;
  assign n16601 = n16600 ^ n14202;
  assign n16602 = n16601 ^ n16543;
  assign n16603 = ~n16544 & n16602;
  assign n16604 = n16603 ^ n14227;
  assign n16605 = n16604 ^ n16541;
  assign n16606 = ~n16542 & ~n16605;
  assign n16607 = n16606 ^ n14256;
  assign n16608 = n16607 ^ n16539;
  assign n16609 = n16540 & ~n16608;
  assign n16610 = n16609 ^ n14254;
  assign n16468 = n16467 ^ n16148;
  assign n16469 = ~n16149 & ~n16468;
  assign n16470 = n16469 ^ n16147;
  assign n16144 = n16026 ^ n15982;
  assign n16142 = n14846 ^ n14826;
  assign n16143 = n16142 ^ n16089;
  assign n16145 = n16144 ^ n16143;
  assign n16537 = n16470 ^ n16145;
  assign n16538 = n16537 ^ n14246;
  assign n16684 = n16610 ^ n16538;
  assign n16685 = n16598 ^ n14202;
  assign n16686 = n16586 ^ n16551;
  assign n16687 = n16580 ^ n13392;
  assign n16688 = n16687 ^ n16555;
  assign n16689 = n16577 ^ n13398;
  assign n16690 = n16572 ^ n16559;
  assign n16695 = ~n16691 & n16694;
  assign n16696 = ~n16690 & n16695;
  assign n16697 = ~n16689 & n16696;
  assign n16698 = ~n16688 & ~n16697;
  assign n16699 = n16583 ^ n13386;
  assign n16700 = n16699 ^ n16553;
  assign n16701 = ~n16698 & n16700;
  assign n16702 = ~n16686 & ~n16701;
  assign n16703 = n16589 ^ n16548;
  assign n16704 = n16702 & n16703;
  assign n16705 = n16592 ^ n16546;
  assign n16706 = n16704 & n16705;
  assign n16707 = ~n16685 & ~n16706;
  assign n16708 = n16601 ^ n16544;
  assign n16709 = ~n16707 & n16708;
  assign n16710 = n16604 ^ n16542;
  assign n16711 = ~n16709 & ~n16710;
  assign n16712 = n16607 ^ n16540;
  assign n16713 = ~n16711 & n16712;
  assign n16714 = n16684 & n16713;
  assign n16611 = n16610 ^ n16537;
  assign n16612 = n16538 & ~n16611;
  assign n16613 = n16612 ^ n14246;
  assign n16682 = n16613 ^ n14245;
  assign n16471 = n16470 ^ n16144;
  assign n16472 = n16145 & n16471;
  assign n16473 = n16472 ^ n16143;
  assign n16137 = n15330 ^ n14842;
  assign n16139 = n16138 ^ n16137;
  assign n16534 = n16473 ^ n16139;
  assign n16140 = n16031 ^ n2206;
  assign n16535 = n16534 ^ n16140;
  assign n16683 = n16682 ^ n16535;
  assign n16846 = n16714 ^ n16683;
  assign n16757 = n16713 ^ n16684;
  assign n16761 = n16760 ^ n16757;
  assign n16762 = n16712 ^ n16711;
  assign n16766 = n16765 ^ n16762;
  assign n16767 = n16710 ^ n16709;
  assign n16771 = n16770 ^ n16767;
  assign n16772 = n16708 ^ n16707;
  assign n16773 = n16772 ^ n584;
  assign n16826 = n16706 ^ n16685;
  assign n16821 = n16705 ^ n16704;
  assign n16774 = n16703 ^ n16702;
  assign n16775 = n16774 ^ n1895;
  assign n16776 = n16701 ^ n16686;
  assign n16777 = n16776 ^ n1906;
  assign n16778 = n16700 ^ n16698;
  assign n16779 = n16778 ^ n1769;
  assign n16780 = n16697 ^ n16688;
  assign n16781 = n16780 ^ n1683;
  assign n16782 = n16696 ^ n16689;
  assign n16783 = n16782 ^ n1671;
  assign n16784 = n16695 ^ n16690;
  assign n16785 = n16784 ^ n1665;
  assign n16800 = n16799 ^ n16794;
  assign n16801 = n16798 & n16800;
  assign n16802 = n16801 ^ n16797;
  assign n16803 = n16802 ^ n16784;
  assign n16804 = ~n16785 & n16803;
  assign n16805 = n16804 ^ n1665;
  assign n16806 = n16805 ^ n16782;
  assign n16807 = ~n16783 & n16806;
  assign n16808 = n16807 ^ n1671;
  assign n16809 = n16808 ^ n16780;
  assign n16810 = ~n16781 & n16809;
  assign n16811 = n16810 ^ n1683;
  assign n16812 = n16811 ^ n16778;
  assign n16813 = ~n16779 & n16812;
  assign n16814 = n16813 ^ n1769;
  assign n16815 = n16814 ^ n16776;
  assign n16816 = ~n16777 & n16815;
  assign n16817 = n16816 ^ n1906;
  assign n16818 = n16817 ^ n16774;
  assign n16819 = ~n16775 & n16818;
  assign n16820 = n16819 ^ n1895;
  assign n16822 = n16821 ^ n16820;
  assign n16823 = n16821 ^ n2076;
  assign n16824 = n16822 & ~n16823;
  assign n16825 = n16824 ^ n2076;
  assign n16827 = n16826 ^ n16825;
  assign n16831 = n16830 ^ n16826;
  assign n16832 = ~n16827 & n16831;
  assign n16833 = n16832 ^ n16830;
  assign n16834 = n16833 ^ n16772;
  assign n16835 = n16773 & ~n16834;
  assign n16836 = n16835 ^ n584;
  assign n16837 = n16836 ^ n16767;
  assign n16838 = n16771 & ~n16837;
  assign n16839 = n16838 ^ n16770;
  assign n16840 = n16839 ^ n16762;
  assign n16841 = n16766 & ~n16840;
  assign n16842 = n16841 ^ n16765;
  assign n16843 = n16842 ^ n16757;
  assign n16844 = ~n16761 & n16843;
  assign n16845 = n16844 ^ n16760;
  assign n16847 = n16846 ^ n16845;
  assign n16851 = n16850 ^ n16846;
  assign n16852 = n16847 & ~n16851;
  assign n16853 = n16852 ^ n16850;
  assign n16536 = n16535 ^ n14245;
  assign n16614 = n16613 ^ n16535;
  assign n16615 = n16536 & ~n16614;
  assign n16616 = n16615 ^ n14245;
  assign n16716 = n16616 ^ n14234;
  assign n16141 = n16140 ^ n16139;
  assign n16474 = n16473 ^ n16140;
  assign n16475 = ~n16141 & n16474;
  assign n16476 = n16475 ^ n16139;
  assign n16132 = n15414 ^ n14233;
  assign n16134 = n16133 ^ n16132;
  assign n16531 = n16476 ^ n16134;
  assign n16135 = n16034 ^ n15980;
  assign n16532 = n16531 ^ n16135;
  assign n16717 = n16716 ^ n16532;
  assign n16715 = n16683 & n16714;
  assign n16755 = n16717 ^ n16715;
  assign n16756 = n16755 ^ n668;
  assign n16969 = n16853 ^ n16756;
  assign n16972 = n16971 ^ n16969;
  assign n16975 = n16850 ^ n16847;
  assign n16973 = n16104 ^ n15558;
  assign n16510 = n16362 ^ n912;
  assign n16511 = n16510 ^ n16358;
  assign n16974 = n16973 ^ n16511;
  assign n16976 = n16975 ^ n16974;
  assign n16979 = n16842 ^ n16761;
  assign n16977 = n16109 ^ n15543;
  assign n16096 = n16095 ^ n16079;
  assign n16978 = n16977 ^ n16096;
  assign n16980 = n16979 ^ n16978;
  assign n16097 = n16076 ^ n557;
  assign n16983 = n16114 ^ n16097;
  assign n16984 = n16983 ^ n15501;
  assign n16981 = n16839 ^ n16765;
  assign n16982 = n16981 ^ n16762;
  assign n16985 = n16984 ^ n16982;
  assign n16102 = n16057 ^ n15964;
  assign n16987 = n16119 ^ n16102;
  assign n16988 = n16987 ^ n15423;
  assign n16986 = n16836 ^ n16771;
  assign n16989 = n16988 ^ n16986;
  assign n16992 = n16833 ^ n16773;
  assign n16107 = n16054 ^ n15966;
  assign n16990 = n16107 ^ n15414;
  assign n16991 = n16990 ^ n16124;
  assign n16993 = n16992 ^ n16991;
  assign n16995 = n16129 ^ n15330;
  assign n16112 = n16051 ^ n15968;
  assign n16996 = n16995 ^ n16112;
  assign n16994 = n16830 ^ n16827;
  assign n16997 = n16996 ^ n16994;
  assign n16117 = n16048 ^ n15970;
  assign n16999 = n16133 ^ n16117;
  assign n17000 = n16999 ^ n14826;
  assign n16998 = n16822 ^ n2076;
  assign n17001 = n17000 ^ n16998;
  assign n17003 = n16138 ^ n15401;
  assign n16122 = n16045 ^ n15975;
  assign n17004 = n17003 ^ n16122;
  assign n17002 = n16817 ^ n16775;
  assign n17005 = n17004 ^ n17002;
  assign n17008 = n16069 ^ n15391;
  assign n17009 = n17008 ^ n16135;
  assign n16926 = n16811 ^ n1769;
  assign n16927 = n16926 ^ n16778;
  assign n17010 = n17009 ^ n16927;
  assign n17011 = n15918 ^ n15341;
  assign n17012 = n17011 ^ n16140;
  assign n16932 = n16808 ^ n16781;
  assign n17013 = n17012 ^ n16932;
  assign n17014 = n15831 ^ n15347;
  assign n17015 = n17014 ^ n16144;
  assign n16937 = n16805 ^ n16783;
  assign n17016 = n17015 ^ n16937;
  assign n17018 = n15378 ^ n15310;
  assign n17019 = n17018 ^ n16148;
  assign n17017 = n16802 ^ n16785;
  assign n17020 = n17019 ^ n17017;
  assign n17022 = n15349 ^ n15311;
  assign n17023 = n17022 ^ n16152;
  assign n17024 = n17023 ^ n17021;
  assign n17026 = n15319 ^ n15312;
  assign n17027 = n17026 ^ n16458;
  assign n17025 = n16791 ^ n16790;
  assign n17028 = n17027 ^ n17025;
  assign n17031 = n16692 ^ n1430;
  assign n17029 = n15353 ^ n15313;
  assign n17030 = n17029 ^ n16154;
  assign n17032 = n17031 ^ n17030;
  assign n17090 = n15325 ^ n15314;
  assign n17091 = n17090 ^ n16158;
  assign n17053 = n14835 ^ n14240;
  assign n17054 = n17053 ^ n15738;
  assign n17036 = n15122 ^ n14536;
  assign n17037 = n17036 ^ n15701;
  assign n16954 = n16375 ^ n1223;
  assign n16955 = n16954 ^ n16351;
  assign n17048 = n17037 ^ n16955;
  assign n16901 = n16372 ^ n16354;
  assign n16899 = n15145 ^ n14505;
  assign n16900 = n16899 ^ n15712;
  assign n16902 = n16901 ^ n16900;
  assign n16669 = n16368 ^ n1049;
  assign n16670 = n16669 ^ n16355;
  assign n16656 = n15133 ^ n14453;
  assign n16657 = n16656 ^ n16397;
  assign n16658 = n16657 ^ n16655;
  assign n16507 = n16180 ^ n15128;
  assign n16508 = n16507 ^ n14429;
  assign n16650 = n16511 ^ n16508;
  assign n16098 = n15726 ^ n15026;
  assign n16100 = n16099 ^ n16098;
  assign n16101 = n16100 ^ n16097;
  assign n16103 = n15692 ^ n14988;
  assign n16105 = n16104 ^ n16103;
  assign n16106 = n16105 ^ n16102;
  assign n16108 = n15672 ^ n14917;
  assign n16110 = n16109 ^ n16108;
  assign n16111 = n16110 ^ n16107;
  assign n16113 = n15558 ^ n14838;
  assign n16115 = n16114 ^ n16113;
  assign n16116 = n16115 ^ n16112;
  assign n16118 = n15543 ^ n14904;
  assign n16120 = n16119 ^ n16118;
  assign n16121 = n16120 ^ n16117;
  assign n16123 = n15501 ^ n14897;
  assign n16125 = n16124 ^ n16123;
  assign n16126 = n16125 ^ n16122;
  assign n16128 = n15423 ^ n14839;
  assign n16130 = n16129 ^ n16128;
  assign n16127 = n16042 ^ n16039;
  assign n16131 = n16130 ^ n16127;
  assign n16136 = n16135 ^ n16134;
  assign n16477 = n16476 ^ n16135;
  assign n16478 = ~n16136 & ~n16477;
  assign n16479 = n16478 ^ n16134;
  assign n16480 = n16479 ^ n16127;
  assign n16481 = n16131 & n16480;
  assign n16482 = n16481 ^ n16130;
  assign n16483 = n16482 ^ n16122;
  assign n16484 = n16126 & ~n16483;
  assign n16485 = n16484 ^ n16125;
  assign n16486 = n16485 ^ n16117;
  assign n16487 = ~n16121 & n16486;
  assign n16488 = n16487 ^ n16120;
  assign n16489 = n16488 ^ n16112;
  assign n16490 = n16116 & n16489;
  assign n16491 = n16490 ^ n16115;
  assign n16492 = n16491 ^ n16107;
  assign n16493 = n16111 & ~n16492;
  assign n16494 = n16493 ^ n16110;
  assign n16495 = n16494 ^ n16102;
  assign n16496 = n16106 & n16495;
  assign n16497 = n16496 ^ n16105;
  assign n16498 = n16497 ^ n16097;
  assign n16499 = n16101 & n16498;
  assign n16500 = n16499 ^ n16100;
  assign n16501 = n16500 ^ n16096;
  assign n16502 = n15761 ^ n15111;
  assign n16503 = n16502 ^ n16184;
  assign n16504 = n16503 ^ n16096;
  assign n16505 = ~n16501 & ~n16504;
  assign n16506 = n16505 ^ n16503;
  assign n16651 = n16511 ^ n16506;
  assign n16652 = n16650 & ~n16651;
  assign n16653 = n16652 ^ n16508;
  assign n16666 = n16657 ^ n16653;
  assign n16667 = ~n16658 & ~n16666;
  assign n16668 = n16667 ^ n16655;
  assign n16671 = n16670 ^ n16668;
  assign n16664 = n15137 ^ n14478;
  assign n16665 = n16664 ^ n15707;
  assign n16896 = n16670 ^ n16665;
  assign n16897 = n16671 & ~n16896;
  assign n16898 = n16897 ^ n16665;
  assign n17033 = n16901 ^ n16898;
  assign n17034 = n16902 & n17033;
  assign n17035 = n17034 ^ n16900;
  assign n17049 = n17035 ^ n16955;
  assign n17050 = ~n17048 & n17049;
  assign n17051 = n17050 ^ n17037;
  assign n16949 = n16378 ^ n16350;
  assign n17052 = n17051 ^ n16949;
  assign n17055 = n17054 ^ n17052;
  assign n17056 = n17055 ^ n13430;
  assign n17038 = n17037 ^ n17035;
  assign n17039 = n17038 ^ n16955;
  assign n17040 = n17039 ^ n13936;
  assign n16903 = n16902 ^ n16898;
  assign n17041 = n16903 ^ n13888;
  assign n16672 = n16671 ^ n16665;
  assign n16659 = n16658 ^ n16653;
  assign n16509 = n16508 ^ n16506;
  assign n16512 = n16511 ^ n16509;
  assign n16513 = n16512 ^ n13903;
  assign n16514 = n16503 ^ n16501;
  assign n16515 = n16514 ^ n14531;
  assign n16516 = n16497 ^ n16101;
  assign n16517 = n16516 ^ n14498;
  assign n16518 = n16494 ^ n16106;
  assign n16519 = n16518 ^ n14467;
  assign n16520 = n16491 ^ n16110;
  assign n16521 = n16520 ^ n16107;
  assign n16522 = n16521 ^ n14446;
  assign n16523 = n16488 ^ n16115;
  assign n16524 = n16523 ^ n16112;
  assign n16525 = n16524 ^ n14422;
  assign n16626 = n16485 ^ n16120;
  assign n16627 = n16626 ^ n16117;
  assign n16526 = n16482 ^ n16126;
  assign n16527 = n16526 ^ n14334;
  assign n16528 = n16479 ^ n16130;
  assign n16529 = n16528 ^ n16127;
  assign n16530 = n16529 ^ n14288;
  assign n16533 = n16532 ^ n14234;
  assign n16617 = n16616 ^ n16532;
  assign n16618 = ~n16533 & ~n16617;
  assign n16619 = n16618 ^ n14234;
  assign n16620 = n16619 ^ n16529;
  assign n16621 = n16530 & n16620;
  assign n16622 = n16621 ^ n14288;
  assign n16623 = n16622 ^ n16526;
  assign n16624 = ~n16527 & n16623;
  assign n16625 = n16624 ^ n14334;
  assign n16628 = n16627 ^ n16625;
  assign n16629 = n16627 ^ n14401;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631 = n16630 ^ n14401;
  assign n16632 = n16631 ^ n16524;
  assign n16633 = ~n16525 & ~n16632;
  assign n16634 = n16633 ^ n14422;
  assign n16635 = n16634 ^ n16521;
  assign n16636 = ~n16522 & ~n16635;
  assign n16637 = n16636 ^ n14446;
  assign n16638 = n16637 ^ n16518;
  assign n16639 = n16519 & n16638;
  assign n16640 = n16639 ^ n14467;
  assign n16641 = n16640 ^ n16516;
  assign n16642 = ~n16517 & n16641;
  assign n16643 = n16642 ^ n14498;
  assign n16644 = n16643 ^ n16514;
  assign n16645 = ~n16515 & n16644;
  assign n16646 = n16645 ^ n14531;
  assign n16647 = n16646 ^ n16512;
  assign n16648 = ~n16513 & n16647;
  assign n16649 = n16648 ^ n13903;
  assign n16660 = n16659 ^ n16649;
  assign n16661 = n16659 ^ n13898;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = n16662 ^ n13898;
  assign n16673 = n16672 ^ n16663;
  assign n16892 = n16672 ^ n13893;
  assign n16893 = ~n16673 & n16892;
  assign n16894 = n16893 ^ n13893;
  assign n17042 = n16903 ^ n16894;
  assign n17043 = n17041 & n17042;
  assign n17044 = n17043 ^ n13888;
  assign n17045 = n17044 ^ n17039;
  assign n17046 = n17040 & ~n17045;
  assign n17047 = n17046 ^ n13936;
  assign n17057 = n17056 ^ n17047;
  assign n16895 = n16894 ^ n13888;
  assign n16904 = n16903 ^ n16895;
  assign n16674 = n16673 ^ n13893;
  assign n16675 = n16660 ^ n13898;
  assign n16676 = n16640 ^ n14498;
  assign n16677 = n16676 ^ n16516;
  assign n16678 = n16637 ^ n14467;
  assign n16679 = n16678 ^ n16518;
  assign n16680 = n16631 ^ n16525;
  assign n16681 = n16619 ^ n16530;
  assign n16718 = n16715 & ~n16717;
  assign n16719 = n16681 & ~n16718;
  assign n16720 = n16622 ^ n14334;
  assign n16721 = n16720 ^ n16526;
  assign n16722 = n16719 & n16721;
  assign n16723 = n16628 ^ n14401;
  assign n16724 = ~n16722 & ~n16723;
  assign n16725 = n16680 & n16724;
  assign n16726 = n16634 ^ n16522;
  assign n16727 = ~n16725 & n16726;
  assign n16728 = ~n16679 & ~n16727;
  assign n16729 = ~n16677 & n16728;
  assign n16730 = n16643 ^ n16515;
  assign n16731 = ~n16729 & n16730;
  assign n16732 = n16646 ^ n16513;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = ~n16675 & n16733;
  assign n16905 = ~n16674 & n16734;
  assign n17058 = n16904 & ~n16905;
  assign n17059 = n17044 ^ n17040;
  assign n17060 = ~n17058 & n17059;
  assign n17087 = ~n17057 & n17060;
  assign n17082 = n14831 ^ n14549;
  assign n17083 = n17082 ^ n15766;
  assign n17079 = n17054 ^ n16949;
  assign n17080 = ~n17052 & n17079;
  assign n17081 = n17080 ^ n17054;
  assign n17084 = n17083 ^ n17081;
  assign n16943 = n16381 ^ n16348;
  assign n17085 = n17084 ^ n16943;
  assign n17075 = n17055 ^ n17047;
  assign n17076 = ~n17056 & n17075;
  assign n17077 = n17076 ^ n13430;
  assign n17078 = n17077 ^ n13424;
  assign n17086 = n17085 ^ n17078;
  assign n17088 = n17087 ^ n17086;
  assign n17061 = n17060 ^ n17057;
  assign n17062 = n17061 ^ n1517;
  assign n17063 = n17059 ^ n17058;
  assign n2564 = n2484 ^ x291;
  assign n2565 = n2564 ^ x483;
  assign n2566 = n2565 ^ x227;
  assign n17064 = n17063 ^ n2566;
  assign n16906 = n16905 ^ n16904;
  assign n16907 = n16906 ^ n2409;
  assign n16735 = n16734 ^ n16674;
  assign n16736 = n16735 ^ n2343;
  assign n16737 = n16733 ^ n16675;
  assign n16738 = n16737 ^ n2331;
  assign n16739 = n16732 ^ n16731;
  assign n1349 = n1243 ^ x295;
  assign n1350 = n1349 ^ x487;
  assign n1351 = n1350 ^ x231;
  assign n16740 = n16739 ^ n1351;
  assign n16741 = n16730 ^ n16729;
  assign n16742 = n16741 ^ n1196;
  assign n16743 = n16728 ^ n16677;
  assign n16744 = n16743 ^ n1178;
  assign n16745 = n16727 ^ n16679;
  assign n16746 = n16745 ^ n944;
  assign n16747 = n16726 ^ n16725;
  assign n16748 = n16747 ^ n1162;
  assign n16866 = n16724 ^ n16680;
  assign n16749 = n16723 ^ n16722;
  assign n16750 = n16749 ^ n724;
  assign n16751 = n16721 ^ n16719;
  assign n16752 = n16751 ^ n717;
  assign n16753 = n16718 ^ n16681;
  assign n16754 = n16753 ^ n674;
  assign n16854 = n16853 ^ n16755;
  assign n16855 = n16756 & ~n16854;
  assign n16856 = n16855 ^ n668;
  assign n16857 = n16856 ^ n16753;
  assign n16858 = ~n16754 & n16857;
  assign n16859 = n16858 ^ n674;
  assign n16860 = n16859 ^ n16751;
  assign n16861 = n16752 & ~n16860;
  assign n16862 = n16861 ^ n717;
  assign n16863 = n16862 ^ n16749;
  assign n16864 = ~n16750 & n16863;
  assign n16865 = n16864 ^ n724;
  assign n16867 = n16866 ^ n16865;
  assign n16868 = n16866 ^ n816;
  assign n16869 = n16867 & ~n16868;
  assign n16870 = n16869 ^ n816;
  assign n16871 = n16870 ^ n16747;
  assign n16872 = ~n16748 & n16871;
  assign n16873 = n16872 ^ n1162;
  assign n16874 = n16873 ^ n16745;
  assign n16875 = ~n16746 & n16874;
  assign n16876 = n16875 ^ n944;
  assign n16877 = n16876 ^ n16743;
  assign n16878 = n16744 & ~n16877;
  assign n16879 = n16878 ^ n1178;
  assign n16880 = n16879 ^ n16741;
  assign n16881 = ~n16742 & n16880;
  assign n16882 = n16881 ^ n1196;
  assign n16883 = n16882 ^ n16739;
  assign n16884 = ~n16740 & n16883;
  assign n16885 = n16884 ^ n1351;
  assign n16886 = n16885 ^ n16737;
  assign n16887 = n16738 & ~n16886;
  assign n16888 = n16887 ^ n2331;
  assign n16889 = n16888 ^ n16735;
  assign n16890 = n16736 & ~n16889;
  assign n16891 = n16890 ^ n2343;
  assign n17065 = n16906 ^ n16891;
  assign n17066 = ~n16907 & n17065;
  assign n17067 = n17066 ^ n2409;
  assign n17068 = n17067 ^ n17063;
  assign n17069 = n17064 & ~n17068;
  assign n17070 = n17069 ^ n2566;
  assign n17071 = n17070 ^ n17061;
  assign n17072 = n17062 & ~n17071;
  assign n17073 = n17072 ^ n1517;
  assign n17074 = n17073 ^ n2642;
  assign n17089 = n17088 ^ n17074;
  assign n17092 = n17091 ^ n17089;
  assign n17094 = n15315 ^ n15300;
  assign n17095 = n17094 ^ n16162;
  assign n17093 = n17070 ^ n17062;
  assign n17096 = n17095 ^ n17093;
  assign n17100 = n17067 ^ n17064;
  assign n16911 = n15322 ^ n14830;
  assign n16912 = n16911 ^ n16174;
  assign n16913 = n16888 ^ n16736;
  assign n16914 = ~n16912 & n16913;
  assign n16909 = n15317 ^ n15205;
  assign n16910 = n16909 ^ n16170;
  assign n16915 = n16914 ^ n16910;
  assign n16908 = n16907 ^ n16891;
  assign n17097 = n16910 ^ n16908;
  assign n17098 = n16915 & n17097;
  assign n17099 = n17098 ^ n16914;
  assign n17101 = n17100 ^ n17099;
  assign n17102 = n15316 ^ n15237;
  assign n17103 = n17102 ^ n16166;
  assign n17104 = n17103 ^ n17100;
  assign n17105 = ~n17101 & ~n17104;
  assign n17106 = n17105 ^ n17103;
  assign n17107 = n17106 ^ n17093;
  assign n17108 = ~n17096 & n17107;
  assign n17109 = n17108 ^ n17095;
  assign n17110 = n17109 ^ n17089;
  assign n17111 = ~n17092 & n17110;
  assign n17112 = n17111 ^ n17091;
  assign n17113 = n17112 ^ n17031;
  assign n17114 = ~n17032 & n17113;
  assign n17115 = n17114 ^ n17030;
  assign n17116 = n17115 ^ n17025;
  assign n17117 = ~n17028 & ~n17116;
  assign n17118 = n17117 ^ n17027;
  assign n17119 = n17118 ^ n17021;
  assign n17120 = n17024 & n17119;
  assign n17121 = n17120 ^ n17023;
  assign n17122 = n17121 ^ n17017;
  assign n17123 = n17020 & ~n17122;
  assign n17124 = n17123 ^ n17019;
  assign n17125 = n17124 ^ n16937;
  assign n17126 = n17016 & ~n17125;
  assign n17127 = n17126 ^ n17015;
  assign n17128 = n17127 ^ n16932;
  assign n17129 = ~n17013 & ~n17128;
  assign n17130 = n17129 ^ n17012;
  assign n17131 = n17130 ^ n16927;
  assign n17132 = n17010 & n17131;
  assign n17133 = n17132 ^ n17009;
  assign n17006 = n16089 ^ n15337;
  assign n17007 = n17006 ^ n16127;
  assign n17134 = n17133 ^ n17007;
  assign n17135 = n16814 ^ n16777;
  assign n17136 = n17135 ^ n17133;
  assign n17137 = n17134 & ~n17136;
  assign n17138 = n17137 ^ n17007;
  assign n17139 = n17138 ^ n17002;
  assign n17140 = n17005 & ~n17139;
  assign n17141 = n17140 ^ n17004;
  assign n17142 = n17141 ^ n16998;
  assign n17143 = n17001 & ~n17142;
  assign n17144 = n17143 ^ n17000;
  assign n17145 = n17144 ^ n16994;
  assign n17146 = n16997 & n17145;
  assign n17147 = n17146 ^ n16996;
  assign n17148 = n17147 ^ n16991;
  assign n17149 = ~n16993 & n17148;
  assign n17150 = n17149 ^ n17147;
  assign n17151 = n17150 ^ n16988;
  assign n17152 = ~n16989 & n17151;
  assign n17153 = n17152 ^ n17150;
  assign n17154 = n17153 ^ n16984;
  assign n17155 = ~n16985 & n17154;
  assign n17156 = n17155 ^ n17153;
  assign n17157 = n17156 ^ n16979;
  assign n17158 = n16980 & n17157;
  assign n17159 = n17158 ^ n16978;
  assign n17160 = n17159 ^ n16974;
  assign n17161 = ~n16976 & n17160;
  assign n17162 = n17161 ^ n16975;
  assign n17163 = n17162 ^ n16969;
  assign n17164 = ~n16972 & n17163;
  assign n17165 = n17164 ^ n16971;
  assign n16964 = n16670 ^ n15692;
  assign n16965 = n16964 ^ n16184;
  assign n17201 = n17165 ^ n16965;
  assign n16966 = n16856 ^ n674;
  assign n16967 = n16966 ^ n16753;
  assign n17202 = n17201 ^ n16967;
  assign n17203 = n17202 ^ n14988;
  assign n17204 = n17162 ^ n16971;
  assign n17205 = n17204 ^ n16969;
  assign n17206 = n17205 ^ n14917;
  assign n17306 = n17159 ^ n16976;
  assign n17207 = n17156 ^ n16980;
  assign n17208 = n17207 ^ n14904;
  assign n17209 = n17153 ^ n16985;
  assign n17210 = n17209 ^ n14897;
  assign n17211 = n17150 ^ n16989;
  assign n17212 = n17211 ^ n14839;
  assign n17213 = n17147 ^ n16993;
  assign n17214 = n17213 ^ n14233;
  assign n17215 = n17144 ^ n16996;
  assign n17216 = n17215 ^ n16994;
  assign n17217 = n17216 ^ n14842;
  assign n17218 = n17141 ^ n17000;
  assign n17219 = n17218 ^ n16998;
  assign n17220 = n17219 ^ n14846;
  assign n17282 = n17138 ^ n17004;
  assign n17283 = n17282 ^ n17002;
  assign n17221 = n17135 ^ n17007;
  assign n17222 = n17221 ^ n17133;
  assign n17223 = n17222 ^ n14852;
  assign n17224 = n17130 ^ n17010;
  assign n17225 = n17224 ^ n14866;
  assign n17226 = n17127 ^ n17012;
  assign n17227 = n17226 ^ n16932;
  assign n17228 = n17227 ^ n14858;
  assign n17268 = n17124 ^ n17016;
  assign n17229 = n17121 ^ n17020;
  assign n17230 = n17229 ^ n14711;
  assign n17231 = n17118 ^ n17024;
  assign n17232 = n17231 ^ n14697;
  assign n17233 = n17115 ^ n17028;
  assign n17234 = n17233 ^ n14658;
  assign n17235 = n17112 ^ n17030;
  assign n17236 = n17235 ^ n17031;
  assign n17237 = n17236 ^ n14589;
  assign n17251 = n17109 ^ n17092;
  assign n17238 = n17106 ^ n17096;
  assign n17239 = n17238 ^ n14236;
  assign n17240 = n17103 ^ n17101;
  assign n17241 = n17240 ^ n14570;
  assign n16917 = n16913 ^ n16912;
  assign n16918 = ~n14556 & ~n16917;
  assign n16919 = n16918 ^ n14563;
  assign n16916 = n16915 ^ n16908;
  assign n17242 = n16918 ^ n16916;
  assign n17243 = n16919 & n17242;
  assign n17244 = n17243 ^ n14563;
  assign n17245 = n17244 ^ n17240;
  assign n17246 = n17241 & n17245;
  assign n17247 = n17246 ^ n14570;
  assign n17248 = n17247 ^ n17238;
  assign n17249 = n17239 & n17248;
  assign n17250 = n17249 ^ n14236;
  assign n17252 = n17251 ^ n17250;
  assign n17253 = n17251 ^ n14580;
  assign n17254 = ~n17252 & ~n17253;
  assign n17255 = n17254 ^ n14580;
  assign n17256 = n17255 ^ n17236;
  assign n17257 = ~n17237 & n17256;
  assign n17258 = n17257 ^ n14589;
  assign n17259 = n17258 ^ n17233;
  assign n17260 = ~n17234 & n17259;
  assign n17261 = n17260 ^ n14658;
  assign n17262 = n17261 ^ n17231;
  assign n17263 = ~n17232 & n17262;
  assign n17264 = n17263 ^ n14697;
  assign n17265 = n17264 ^ n17229;
  assign n17266 = n17230 & ~n17265;
  assign n17267 = n17266 ^ n14711;
  assign n17269 = n17268 ^ n17267;
  assign n17270 = n17268 ^ n14818;
  assign n17271 = ~n17269 & n17270;
  assign n17272 = n17271 ^ n14818;
  assign n17273 = n17272 ^ n17227;
  assign n17274 = ~n17228 & n17273;
  assign n17275 = n17274 ^ n14858;
  assign n17276 = n17275 ^ n17224;
  assign n17277 = n17225 & n17276;
  assign n17278 = n17277 ^ n14866;
  assign n17279 = n17278 ^ n17222;
  assign n17280 = n17223 & n17279;
  assign n17281 = n17280 ^ n14852;
  assign n17284 = n17283 ^ n17281;
  assign n17285 = n17283 ^ n14850;
  assign n17286 = ~n17284 & ~n17285;
  assign n17287 = n17286 ^ n14850;
  assign n17288 = n17287 ^ n17219;
  assign n17289 = ~n17220 & n17288;
  assign n17290 = n17289 ^ n14846;
  assign n17291 = n17290 ^ n17216;
  assign n17292 = ~n17217 & n17291;
  assign n17293 = n17292 ^ n14842;
  assign n17294 = n17293 ^ n17213;
  assign n17295 = ~n17214 & ~n17294;
  assign n17296 = n17295 ^ n14233;
  assign n17297 = n17296 ^ n17211;
  assign n17298 = n17212 & n17297;
  assign n17299 = n17298 ^ n14839;
  assign n17300 = n17299 ^ n17209;
  assign n17301 = ~n17210 & ~n17300;
  assign n17302 = n17301 ^ n14897;
  assign n17303 = n17302 ^ n17207;
  assign n17304 = ~n17208 & n17303;
  assign n17305 = n17304 ^ n14904;
  assign n17307 = n17306 ^ n17305;
  assign n17308 = n17306 ^ n14838;
  assign n17309 = n17307 & ~n17308;
  assign n17310 = n17309 ^ n14838;
  assign n17311 = n17310 ^ n17205;
  assign n17312 = ~n17206 & n17311;
  assign n17313 = n17312 ^ n14917;
  assign n17314 = n17313 ^ n17202;
  assign n17315 = ~n17203 & n17314;
  assign n17316 = n17315 ^ n14988;
  assign n17359 = n17316 ^ n15026;
  assign n16968 = n16967 ^ n16965;
  assign n17166 = n17165 ^ n16967;
  assign n17167 = ~n16968 & ~n17166;
  assign n17168 = n17167 ^ n16965;
  assign n16962 = n16859 ^ n16752;
  assign n16960 = n16901 ^ n15726;
  assign n16961 = n16960 ^ n16180;
  assign n16963 = n16962 ^ n16961;
  assign n17199 = n17168 ^ n16963;
  assign n17360 = n17359 ^ n17199;
  assign n17361 = n17302 ^ n17208;
  assign n17362 = n17299 ^ n17210;
  assign n17363 = n17296 ^ n14839;
  assign n17364 = n17363 ^ n17211;
  assign n17365 = n17293 ^ n17214;
  assign n17366 = n17287 ^ n14846;
  assign n17367 = n17366 ^ n17219;
  assign n17368 = n17278 ^ n14852;
  assign n17369 = n17368 ^ n17222;
  assign n17370 = n17272 ^ n17228;
  assign n17371 = n17269 ^ n14818;
  assign n16920 = n16919 ^ n16916;
  assign n16921 = n16917 ^ n14556;
  assign n17372 = ~n16920 & n16921;
  assign n17373 = n17244 ^ n17241;
  assign n17374 = n17372 & n17373;
  assign n17375 = n17247 ^ n17239;
  assign n17376 = n17374 & ~n17375;
  assign n17377 = n17252 ^ n14580;
  assign n17378 = n17376 & ~n17377;
  assign n17379 = n17255 ^ n14589;
  assign n17380 = n17379 ^ n17236;
  assign n17381 = ~n17378 & ~n17380;
  assign n17382 = n17258 ^ n17234;
  assign n17383 = ~n17381 & n17382;
  assign n17384 = n17261 ^ n17232;
  assign n17385 = ~n17383 & ~n17384;
  assign n17386 = n17264 ^ n17230;
  assign n17387 = n17385 & n17386;
  assign n17388 = n17371 & n17387;
  assign n17389 = n17370 & ~n17388;
  assign n17390 = n17275 ^ n17225;
  assign n17391 = ~n17389 & n17390;
  assign n17392 = n17369 & ~n17391;
  assign n17393 = n17284 ^ n14850;
  assign n17394 = ~n17392 & ~n17393;
  assign n17395 = n17367 & n17394;
  assign n17396 = n17290 ^ n17217;
  assign n17397 = n17395 & n17396;
  assign n17398 = n17365 & n17397;
  assign n17399 = ~n17364 & ~n17398;
  assign n17400 = ~n17362 & n17399;
  assign n17401 = ~n17361 & ~n17400;
  assign n17402 = n17307 ^ n14838;
  assign n17403 = n17401 & ~n17402;
  assign n17404 = n17310 ^ n17206;
  assign n17405 = ~n17403 & n17404;
  assign n17406 = n17313 ^ n17203;
  assign n17407 = ~n17405 & ~n17406;
  assign n17408 = n17360 & n17407;
  assign n17200 = n17199 ^ n15026;
  assign n17317 = n17316 ^ n17199;
  assign n17318 = n17200 & ~n17317;
  assign n17319 = n17318 ^ n15026;
  assign n17169 = n17168 ^ n16961;
  assign n17170 = ~n16963 & n17169;
  assign n17171 = n17170 ^ n16962;
  assign n16956 = n16955 ^ n15761;
  assign n16957 = n16956 ^ n16397;
  assign n17196 = n17171 ^ n16957;
  assign n16958 = n16862 ^ n16750;
  assign n17197 = n17196 ^ n16958;
  assign n17198 = n17197 ^ n15111;
  assign n17409 = n17319 ^ n17198;
  assign n17410 = ~n17408 & n17409;
  assign n17320 = n17319 ^ n17197;
  assign n17321 = ~n17198 & n17320;
  assign n17322 = n17321 ^ n15111;
  assign n16959 = n16958 ^ n16957;
  assign n17172 = n17171 ^ n16958;
  assign n17173 = n16959 & n17172;
  assign n17174 = n17173 ^ n16957;
  assign n16952 = n16867 ^ n816;
  assign n16950 = n16949 ^ n15128;
  assign n16951 = n16950 ^ n15707;
  assign n16953 = n16952 ^ n16951;
  assign n17194 = n17174 ^ n16953;
  assign n17195 = n17194 ^ n14429;
  assign n17411 = n17322 ^ n17195;
  assign n17412 = ~n17410 & ~n17411;
  assign n17323 = n17322 ^ n17194;
  assign n17324 = ~n17195 & n17323;
  assign n17325 = n17324 ^ n14429;
  assign n17175 = n17174 ^ n16951;
  assign n17176 = ~n16953 & n17175;
  assign n17177 = n17176 ^ n16952;
  assign n16946 = n16870 ^ n1162;
  assign n16947 = n16946 ^ n16747;
  assign n16944 = n16943 ^ n15712;
  assign n16945 = n16944 ^ n15133;
  assign n16948 = n16947 ^ n16945;
  assign n17192 = n17177 ^ n16948;
  assign n17193 = n17192 ^ n14453;
  assign n17413 = n17325 ^ n17193;
  assign n17414 = n17412 & n17413;
  assign n17326 = n17325 ^ n17192;
  assign n17327 = n17193 & n17326;
  assign n17328 = n17327 ^ n14453;
  assign n17178 = n17177 ^ n16945;
  assign n17179 = ~n16948 & n17178;
  assign n17180 = n17179 ^ n16947;
  assign n16941 = n16873 ^ n16746;
  assign n16939 = n16418 ^ n15701;
  assign n16940 = n16939 ^ n15137;
  assign n16942 = n16941 ^ n16940;
  assign n17190 = n17180 ^ n16942;
  assign n17191 = n17190 ^ n14478;
  assign n17415 = n17328 ^ n17191;
  assign n17416 = n17414 & n17415;
  assign n17329 = n17328 ^ n17190;
  assign n17330 = ~n17191 & ~n17329;
  assign n17331 = n17330 ^ n14478;
  assign n17185 = n15738 ^ n15145;
  assign n17186 = n17185 ^ n16423;
  assign n17184 = n16876 ^ n16744;
  assign n17187 = n17186 ^ n17184;
  assign n17181 = n17180 ^ n16941;
  assign n17182 = ~n16942 & ~n17181;
  assign n17183 = n17182 ^ n16940;
  assign n17188 = n17187 ^ n17183;
  assign n17189 = n17188 ^ n14505;
  assign n17358 = n17331 ^ n17189;
  assign n17424 = n17416 ^ n17358;
  assign n17425 = n17424 ^ n2515;
  assign n17575 = n17415 ^ n17414;
  assign n17426 = n17413 ^ n17412;
  assign n2274 = n1304 ^ x326;
  assign n2275 = n2274 ^ n2267;
  assign n2276 = n2275 ^ x262;
  assign n17427 = n17426 ^ n2276;
  assign n17429 = n1380 ^ x327;
  assign n17430 = n17429 ^ n1213;
  assign n17431 = n17430 ^ x263;
  assign n17428 = n17411 ^ n17410;
  assign n17432 = n17431 ^ n17428;
  assign n17559 = n17407 ^ n17360;
  assign n17433 = n17406 ^ n17405;
  assign n17434 = n17433 ^ n1033;
  assign n17435 = n17404 ^ n17403;
  assign n17436 = n17435 ^ n886;
  assign n17548 = n17402 ^ n17401;
  assign n17437 = n17400 ^ n17361;
  assign n17438 = n17437 ^ n792;
  assign n17439 = n17399 ^ n17362;
  assign n17440 = n17439 ^ n783;
  assign n17534 = n17398 ^ n17364;
  assign n17441 = n17397 ^ n17365;
  assign n17445 = n17444 ^ n17441;
  assign n17446 = n17396 ^ n17395;
  assign n17447 = n17446 ^ n524;
  assign n17449 = n15592 ^ x338;
  assign n17450 = n17449 ^ n572;
  assign n17451 = n17450 ^ x274;
  assign n17448 = n17394 ^ n17367;
  assign n17452 = n17451 ^ n17448;
  assign n17520 = n17393 ^ n17392;
  assign n17453 = n17391 ^ n17369;
  assign n17457 = n17456 ^ n17453;
  assign n17458 = n17390 ^ n17389;
  assign n17462 = n17461 ^ n17458;
  assign n17463 = n17388 ^ n17370;
  assign n17464 = n17463 ^ n2172;
  assign n17465 = n17387 ^ n17371;
  assign n17466 = n17465 ^ n2017;
  assign n17467 = n17386 ^ n17385;
  assign n17468 = n17467 ^ n2004;
  assign n17500 = n17384 ^ n17383;
  assign n17469 = n17382 ^ n17381;
  assign n17470 = n17469 ^ n1864;
  assign n17471 = n17380 ^ n17378;
  assign n17472 = n17471 ^ n1858;
  assign n17473 = n17377 ^ n17376;
  assign n17474 = n17473 ^ n1623;
  assign n17475 = n17375 ^ n17374;
  assign n17479 = n17478 ^ n17475;
  assign n16923 = n1502 & ~n16921;
  assign n16924 = n16923 ^ n1472;
  assign n16922 = n16921 ^ n16920;
  assign n17480 = n16923 ^ n16922;
  assign n17481 = n16924 & n17480;
  assign n17482 = n17481 ^ n1472;
  assign n17483 = n17482 ^ n1421;
  assign n17484 = n17373 ^ n17372;
  assign n17485 = n17484 ^ n17482;
  assign n17486 = n17483 & ~n17485;
  assign n17487 = n17486 ^ n1421;
  assign n17488 = n17487 ^ n17475;
  assign n17489 = ~n17479 & n17488;
  assign n17490 = n17489 ^ n17478;
  assign n17491 = n17490 ^ n17473;
  assign n17492 = ~n17474 & n17491;
  assign n17493 = n17492 ^ n1623;
  assign n17494 = n17493 ^ n17471;
  assign n17495 = ~n17472 & n17494;
  assign n17496 = n17495 ^ n1858;
  assign n17497 = n17496 ^ n17469;
  assign n17498 = ~n17470 & n17497;
  assign n17499 = n17498 ^ n1864;
  assign n17501 = n17500 ^ n17499;
  assign n17502 = n17500 ^ n1879;
  assign n17503 = n17501 & ~n17502;
  assign n17504 = n17503 ^ n1879;
  assign n17505 = n17504 ^ n17467;
  assign n17506 = ~n17468 & n17505;
  assign n17507 = n17506 ^ n2004;
  assign n17508 = n17507 ^ n17465;
  assign n17509 = ~n17466 & n17508;
  assign n17510 = n17509 ^ n2017;
  assign n17511 = n17510 ^ n17463;
  assign n17512 = ~n17464 & n17511;
  assign n17513 = n17512 ^ n2172;
  assign n17514 = n17513 ^ n17458;
  assign n17515 = n17462 & ~n17514;
  assign n17516 = n17515 ^ n17461;
  assign n17517 = n17516 ^ n17453;
  assign n17518 = ~n17457 & n17517;
  assign n17519 = n17518 ^ n17456;
  assign n17521 = n17520 ^ n17519;
  assign n17522 = n17520 ^ n603;
  assign n17523 = n17521 & ~n17522;
  assign n17524 = n17523 ^ n603;
  assign n17525 = n17524 ^ n17448;
  assign n17526 = ~n17452 & n17525;
  assign n17527 = n17526 ^ n17451;
  assign n17528 = n17527 ^ n17446;
  assign n17529 = ~n17447 & n17528;
  assign n17530 = n17529 ^ n524;
  assign n17531 = n17530 ^ n17441;
  assign n17532 = ~n17445 & n17531;
  assign n17533 = n17532 ^ n17444;
  assign n17535 = n17534 ^ n17533;
  assign n17539 = n17538 ^ n17534;
  assign n17540 = ~n17535 & n17539;
  assign n17541 = n17540 ^ n17538;
  assign n17542 = n17541 ^ n17439;
  assign n17543 = ~n17440 & n17542;
  assign n17544 = n17543 ^ n783;
  assign n17545 = n17544 ^ n17437;
  assign n17546 = ~n17438 & n17545;
  assign n17547 = n17546 ^ n792;
  assign n17549 = n17548 ^ n17547;
  assign n17550 = n17548 ^ n807;
  assign n17551 = ~n17549 & n17550;
  assign n17552 = n17551 ^ n807;
  assign n17553 = n17552 ^ n17435;
  assign n17554 = ~n17436 & n17553;
  assign n17555 = n17554 ^ n886;
  assign n17556 = n17555 ^ n17433;
  assign n17557 = ~n17434 & n17556;
  assign n17558 = n17557 ^ n1033;
  assign n17560 = n17559 ^ n17558;
  assign n17561 = n17559 ^ n1042;
  assign n17562 = n17560 & ~n17561;
  assign n17563 = n17562 ^ n1042;
  assign n1204 = n1113 ^ x328;
  assign n1208 = n1207 ^ n1204;
  assign n1209 = n1208 ^ x264;
  assign n17564 = n17563 ^ n1209;
  assign n17565 = n17409 ^ n17408;
  assign n17566 = n17565 ^ n17563;
  assign n17567 = n17564 & n17566;
  assign n17568 = n17567 ^ n1209;
  assign n17569 = n17568 ^ n17431;
  assign n17570 = ~n17432 & ~n17569;
  assign n17571 = n17570 ^ n17428;
  assign n17572 = n17571 ^ n17426;
  assign n17573 = ~n17427 & ~n17572;
  assign n17574 = n17573 ^ n2276;
  assign n17576 = n17575 ^ n17574;
  assign n2506 = n2452 ^ x325;
  assign n2507 = n2506 ^ n1535;
  assign n2508 = n2507 ^ x261;
  assign n17577 = n17575 ^ n2508;
  assign n17578 = n17576 & ~n17577;
  assign n17579 = n17578 ^ n2508;
  assign n17580 = n17579 ^ n17424;
  assign n17581 = ~n17425 & n17580;
  assign n17582 = n17581 ^ n2515;
  assign n17611 = n17582 ^ n2530;
  assign n17340 = n16879 ^ n1196;
  assign n17341 = n17340 ^ n16741;
  assign n17338 = n16430 ^ n15122;
  assign n17339 = n17338 ^ n15766;
  assign n17342 = n17341 ^ n17339;
  assign n17335 = n17184 ^ n17183;
  assign n17336 = n17187 & ~n17335;
  assign n17337 = n17336 ^ n17186;
  assign n17343 = n17342 ^ n17337;
  assign n17332 = n17331 ^ n17188;
  assign n17333 = ~n17189 & n17332;
  assign n17334 = n17333 ^ n14505;
  assign n17344 = n17343 ^ n17334;
  assign n17418 = n17344 ^ n14536;
  assign n17417 = n17358 & ~n17416;
  assign n17422 = n17418 ^ n17417;
  assign n17612 = n17611 ^ n17422;
  assign n17615 = n17614 ^ n17612;
  assign n17618 = n17576 ^ n2508;
  assign n17619 = n17031 ^ n16166;
  assign n17620 = n17619 ^ n15322;
  assign n17621 = ~n17618 & n17620;
  assign n17616 = n17025 ^ n16162;
  assign n17617 = n17616 ^ n15317;
  assign n17622 = n17621 ^ n17617;
  assign n17623 = n17579 ^ n17425;
  assign n17624 = n17623 ^ n17617;
  assign n17625 = n17622 & n17624;
  assign n17626 = n17625 ^ n17621;
  assign n17627 = n17626 ^ n17612;
  assign n17628 = ~n17615 & ~n17627;
  assign n17629 = n17628 ^ n17614;
  assign n17607 = n16154 ^ n15315;
  assign n17608 = n17607 ^ n17017;
  assign n17655 = n17629 ^ n17608;
  assign n17423 = n17422 ^ n2530;
  assign n17583 = n17582 ^ n17422;
  assign n17584 = n17423 & ~n17583;
  assign n17585 = n17584 ^ n2530;
  assign n17419 = ~n17417 & n17418;
  assign n17354 = n16413 ^ n15770;
  assign n17355 = n17354 ^ n14835;
  assign n17350 = n17341 ^ n17337;
  assign n17351 = n17342 & n17350;
  assign n17352 = n17351 ^ n17339;
  assign n17349 = n16882 ^ n16740;
  assign n17353 = n17352 ^ n17349;
  assign n17356 = n17355 ^ n17353;
  assign n17345 = n17343 ^ n14536;
  assign n17346 = n17344 & n17345;
  assign n17347 = n17346 ^ n14536;
  assign n17348 = n17347 ^ n14240;
  assign n17357 = n17356 ^ n17348;
  assign n17420 = n17419 ^ n17357;
  assign n17421 = n17420 ^ n2632;
  assign n17609 = n17585 ^ n17421;
  assign n17656 = n17655 ^ n17609;
  assign n17657 = n17656 ^ n15300;
  assign n17658 = n17626 ^ n17614;
  assign n17659 = n17658 ^ n17612;
  assign n17660 = n17659 ^ n15237;
  assign n17661 = n17620 ^ n17618;
  assign n17662 = ~n14830 & ~n17661;
  assign n17663 = n17662 ^ n15205;
  assign n17664 = n17623 ^ n17622;
  assign n17665 = n17664 ^ n17662;
  assign n17666 = n17663 & n17665;
  assign n17667 = n17666 ^ n15205;
  assign n17668 = n17667 ^ n17659;
  assign n17669 = n17660 & n17668;
  assign n17670 = n17669 ^ n15237;
  assign n17671 = n17670 ^ n17656;
  assign n17672 = n17657 & ~n17671;
  assign n17673 = n17672 ^ n15300;
  assign n17610 = n17609 ^ n17608;
  assign n17630 = n17629 ^ n17609;
  assign n17631 = n17610 & n17630;
  assign n17632 = n17631 ^ n17608;
  assign n17603 = ~n17357 & n17419;
  assign n17599 = n16885 ^ n16738;
  assign n17597 = n17082 ^ n15323;
  assign n17598 = n17597 ^ n16409;
  assign n17600 = n17599 ^ n17598;
  assign n17593 = n17356 ^ n14240;
  assign n17594 = n17356 ^ n17347;
  assign n17595 = n17593 & ~n17594;
  assign n17596 = n17595 ^ n14240;
  assign n17601 = n17600 ^ n17596;
  assign n17590 = n17355 ^ n17349;
  assign n17591 = ~n17353 & ~n17590;
  assign n17592 = n17591 ^ n17355;
  assign n17602 = n17601 ^ n17592;
  assign n17604 = n17603 ^ n17602;
  assign n17586 = n17585 ^ n17420;
  assign n17587 = n17421 & ~n17586;
  assign n17588 = n17587 ^ n2632;
  assign n17589 = n17588 ^ n2627;
  assign n17605 = n17604 ^ n17589;
  assign n16936 = n16458 ^ n15314;
  assign n16938 = n16937 ^ n16936;
  assign n17606 = n17605 ^ n16938;
  assign n17653 = n17632 ^ n17606;
  assign n17654 = n17653 ^ n15325;
  assign n17698 = n17673 ^ n17654;
  assign n17699 = n17664 ^ n17663;
  assign n17700 = n17661 ^ n14830;
  assign n17701 = ~n17699 & n17700;
  assign n17702 = n17667 ^ n15237;
  assign n17703 = n17702 ^ n17659;
  assign n17704 = n17701 & n17703;
  assign n17705 = n17670 ^ n17657;
  assign n17706 = n17704 & ~n17705;
  assign n17707 = ~n17698 & n17706;
  assign n17674 = n17673 ^ n17653;
  assign n17675 = n17654 & ~n17674;
  assign n17676 = n17675 ^ n15325;
  assign n17633 = n17632 ^ n17605;
  assign n17634 = ~n17606 & n17633;
  assign n17635 = n17634 ^ n16938;
  assign n16933 = n16932 ^ n16152;
  assign n16934 = n16933 ^ n15313;
  assign n16931 = n16921 ^ n1502;
  assign n16935 = n16934 ^ n16931;
  assign n17651 = n17635 ^ n16935;
  assign n17652 = n17651 ^ n15353;
  assign n17708 = n17676 ^ n17652;
  assign n17709 = ~n17707 & n17708;
  assign n17677 = n17676 ^ n17651;
  assign n17678 = n17652 & ~n17677;
  assign n17679 = n17678 ^ n15353;
  assign n17710 = n17679 ^ n15319;
  assign n17636 = n17635 ^ n16931;
  assign n17637 = ~n16935 & n17636;
  assign n17638 = n17637 ^ n16934;
  assign n16928 = n16927 ^ n16148;
  assign n16929 = n16928 ^ n15312;
  assign n17648 = n17638 ^ n16929;
  assign n16925 = n16924 ^ n16922;
  assign n17649 = n17648 ^ n16925;
  assign n17711 = n17710 ^ n17649;
  assign n17712 = ~n17709 & n17711;
  assign n17650 = n17649 ^ n15319;
  assign n17680 = n17679 ^ n17649;
  assign n17681 = ~n17650 & ~n17680;
  assign n17682 = n17681 ^ n15319;
  assign n17644 = n17484 ^ n17483;
  assign n17642 = n17135 ^ n15311;
  assign n17643 = n17642 ^ n16144;
  assign n17645 = n17644 ^ n17643;
  assign n16930 = n16929 ^ n16925;
  assign n17639 = n17638 ^ n16925;
  assign n17640 = ~n16930 & n17639;
  assign n17641 = n17640 ^ n16929;
  assign n17646 = n17645 ^ n17641;
  assign n17647 = n17646 ^ n15349;
  assign n17697 = n17682 ^ n17647;
  assign n17786 = n17712 ^ n17697;
  assign n17749 = n17711 ^ n17709;
  assign n17750 = n17749 ^ n1754;
  assign n17751 = n17708 ^ n17707;
  assign n17752 = n17751 ^ n1657;
  assign n17753 = n17706 ^ n17698;
  assign n17754 = n17753 ^ n1648;
  assign n17755 = n17705 ^ n17704;
  assign n17756 = n17755 ^ n1583;
  assign n17757 = n17703 ^ n17701;
  assign n17758 = n17757 ^ n1574;
  assign n17765 = ~n17700 & n17764;
  assign n17766 = n17765 ^ n17761;
  assign n17767 = n17700 ^ n17699;
  assign n17768 = n17767 ^ n17765;
  assign n17769 = n17766 & n17768;
  assign n17770 = n17769 ^ n17761;
  assign n17771 = n17770 ^ n17757;
  assign n17772 = n17758 & ~n17771;
  assign n17773 = n17772 ^ n1574;
  assign n17774 = n17773 ^ n17755;
  assign n17775 = ~n17756 & n17774;
  assign n17776 = n17775 ^ n1583;
  assign n17777 = n17776 ^ n17753;
  assign n17778 = ~n17754 & n17777;
  assign n17779 = n17778 ^ n1648;
  assign n17780 = n17779 ^ n17751;
  assign n17781 = n17752 & ~n17780;
  assign n17782 = n17781 ^ n1657;
  assign n17783 = n17782 ^ n17749;
  assign n17784 = ~n17750 & n17783;
  assign n17785 = n17784 ^ n1754;
  assign n17787 = n17786 ^ n17785;
  assign n18435 = n17787 ^ n2118;
  assign n18963 = n18435 ^ n16998;
  assign n17860 = n17507 ^ n17466;
  assign n18964 = n18963 ^ n17860;
  assign n18216 = n17021 ^ n16931;
  assign n18217 = n18216 ^ n16166;
  assign n18147 = n17555 ^ n17434;
  assign n18144 = n16430 ^ n15701;
  assign n18145 = n18144 ^ n16913;
  assign n18008 = n17552 ^ n886;
  assign n18009 = n18008 ^ n17435;
  assign n18006 = n16423 ^ n15712;
  assign n18007 = n18006 ^ n17599;
  assign n18010 = n18009 ^ n18007;
  assign n17996 = n17549 ^ n807;
  assign n17918 = n17544 ^ n792;
  assign n17919 = n17918 ^ n17437;
  assign n17916 = n17341 ^ n16397;
  assign n17917 = n17916 ^ n16943;
  assign n17920 = n17919 ^ n17917;
  assign n17829 = n17184 ^ n16949;
  assign n17830 = n17829 ^ n16180;
  assign n17828 = n17541 ^ n17440;
  assign n17831 = n17830 ^ n17828;
  assign n17833 = n16955 ^ n16941;
  assign n17834 = n17833 ^ n16184;
  assign n17832 = n17538 ^ n17535;
  assign n17835 = n17834 ^ n17832;
  assign n17837 = n16901 ^ n16099;
  assign n17838 = n17837 ^ n16947;
  assign n17836 = n17530 ^ n17445;
  assign n17839 = n17838 ^ n17836;
  assign n17842 = n16670 ^ n16104;
  assign n17843 = n17842 ^ n16952;
  assign n17840 = n17527 ^ n524;
  assign n17841 = n17840 ^ n17446;
  assign n17844 = n17843 ^ n17841;
  assign n17847 = n17524 ^ n17451;
  assign n17848 = n17847 ^ n17448;
  assign n17845 = n16655 ^ n16109;
  assign n17846 = n17845 ^ n16958;
  assign n17849 = n17848 ^ n17846;
  assign n17851 = n16511 ^ n16114;
  assign n17852 = n17851 ^ n16962;
  assign n17850 = n17521 ^ n603;
  assign n17853 = n17852 ^ n17850;
  assign n17891 = n17516 ^ n17457;
  assign n17855 = n16975 ^ n16129;
  assign n17856 = n17855 ^ n16102;
  assign n17854 = n17510 ^ n17464;
  assign n17857 = n17856 ^ n17854;
  assign n17858 = n16979 ^ n16107;
  assign n17859 = n17858 ^ n16133;
  assign n17861 = n17860 ^ n17859;
  assign n17872 = n17504 ^ n17468;
  assign n17808 = n16992 ^ n16069;
  assign n17809 = n17808 ^ n16122;
  assign n17806 = n17496 ^ n1864;
  assign n17807 = n17806 ^ n17469;
  assign n17810 = n17809 ^ n17807;
  assign n17737 = n16994 ^ n16127;
  assign n17738 = n17737 ^ n15918;
  assign n17736 = n17493 ^ n17472;
  assign n17739 = n17738 ^ n17736;
  assign n17723 = n16998 ^ n16135;
  assign n17724 = n17723 ^ n15831;
  assign n17722 = n17490 ^ n17474;
  assign n17725 = n17724 ^ n17722;
  assign n17691 = n17643 ^ n17641;
  assign n17692 = n17645 & ~n17691;
  assign n17693 = n17692 ^ n17644;
  assign n17689 = n17487 ^ n17478;
  assign n17690 = n17689 ^ n17475;
  assign n17694 = n17693 ^ n17690;
  assign n17687 = n17002 ^ n15310;
  assign n17688 = n17687 ^ n16140;
  assign n17719 = n17690 ^ n17688;
  assign n17720 = n17694 & n17719;
  assign n17721 = n17720 ^ n17688;
  assign n17733 = n17722 ^ n17721;
  assign n17734 = ~n17725 & ~n17733;
  assign n17735 = n17734 ^ n17724;
  assign n17803 = n17736 ^ n17735;
  assign n17804 = ~n17739 & n17803;
  assign n17805 = n17804 ^ n17738;
  assign n17863 = n17807 ^ n17805;
  assign n17864 = n17810 & n17863;
  assign n17865 = n17864 ^ n17809;
  assign n17862 = n17501 ^ n1879;
  assign n17866 = n17865 ^ n17862;
  assign n17867 = n16986 ^ n16089;
  assign n17868 = n17867 ^ n16117;
  assign n17869 = n17868 ^ n17862;
  assign n17870 = ~n17866 & n17869;
  assign n17871 = n17870 ^ n17868;
  assign n17873 = n17872 ^ n17871;
  assign n17874 = n16982 ^ n16112;
  assign n17875 = n17874 ^ n16138;
  assign n17876 = n17875 ^ n17872;
  assign n17877 = ~n17873 & ~n17876;
  assign n17878 = n17877 ^ n17875;
  assign n17879 = n17878 ^ n17860;
  assign n17880 = ~n17861 & n17879;
  assign n17881 = n17880 ^ n17859;
  assign n17882 = n17881 ^ n17856;
  assign n17883 = n17857 & n17882;
  assign n17884 = n17883 ^ n17854;
  assign n17821 = n17513 ^ n17461;
  assign n17822 = n17821 ^ n17458;
  assign n17885 = n17884 ^ n17822;
  assign n17886 = n16124 ^ n16097;
  assign n17887 = n17886 ^ n16969;
  assign n17888 = n17887 ^ n17822;
  assign n17889 = n17885 & n17888;
  assign n17890 = n17889 ^ n17887;
  assign n17892 = n17891 ^ n17890;
  assign n17893 = n16967 ^ n16119;
  assign n17894 = n17893 ^ n16096;
  assign n17895 = n17894 ^ n17891;
  assign n17896 = n17892 & ~n17895;
  assign n17897 = n17896 ^ n17894;
  assign n17898 = n17897 ^ n17852;
  assign n17899 = n17853 & n17898;
  assign n17900 = n17899 ^ n17850;
  assign n17901 = n17900 ^ n17846;
  assign n17902 = n17849 & ~n17901;
  assign n17903 = n17902 ^ n17848;
  assign n17904 = n17903 ^ n17841;
  assign n17905 = ~n17844 & ~n17904;
  assign n17906 = n17905 ^ n17843;
  assign n17907 = n17906 ^ n17836;
  assign n17908 = ~n17839 & n17907;
  assign n17909 = n17908 ^ n17838;
  assign n17910 = n17909 ^ n17832;
  assign n17911 = n17835 & ~n17910;
  assign n17912 = n17911 ^ n17834;
  assign n17913 = n17912 ^ n17828;
  assign n17914 = ~n17831 & n17913;
  assign n17915 = n17914 ^ n17830;
  assign n17993 = n17919 ^ n17915;
  assign n17994 = ~n17920 & n17993;
  assign n17995 = n17994 ^ n17917;
  assign n17997 = n17996 ^ n17995;
  assign n17991 = n17349 ^ n16418;
  assign n17992 = n17991 ^ n15707;
  assign n18003 = n17996 ^ n17992;
  assign n18004 = ~n17997 & n18003;
  assign n18005 = n18004 ^ n17992;
  assign n18141 = n18007 ^ n18005;
  assign n18142 = n18010 & n18141;
  assign n18143 = n18142 ^ n18009;
  assign n18146 = n18145 ^ n18143;
  assign n18148 = n18147 ^ n18146;
  assign n18149 = n18148 ^ n15137;
  assign n18011 = n18010 ^ n18005;
  assign n17998 = n17997 ^ n17992;
  assign n17921 = n17920 ^ n17915;
  assign n17922 = n17921 ^ n15761;
  assign n17923 = n17912 ^ n17830;
  assign n17924 = n17923 ^ n17828;
  assign n17925 = n17924 ^ n15726;
  assign n17926 = n17909 ^ n17835;
  assign n17927 = n17926 ^ n15692;
  assign n17928 = n17906 ^ n17839;
  assign n17929 = n17928 ^ n15672;
  assign n17930 = n17903 ^ n17844;
  assign n17931 = n17930 ^ n15558;
  assign n17971 = n17900 ^ n17849;
  assign n17966 = n17897 ^ n17853;
  assign n17932 = n17894 ^ n17892;
  assign n17933 = n17932 ^ n15423;
  assign n17958 = n17887 ^ n17885;
  assign n17934 = n17881 ^ n17857;
  assign n17935 = n17934 ^ n15330;
  assign n17936 = n17878 ^ n17859;
  assign n17937 = n17936 ^ n17860;
  assign n17938 = n17937 ^ n14826;
  assign n17939 = n17875 ^ n17873;
  assign n17940 = n17939 ^ n15401;
  assign n17944 = n17868 ^ n17866;
  assign n17811 = n17810 ^ n17805;
  assign n17812 = n17811 ^ n15391;
  assign n17740 = n17739 ^ n17735;
  assign n17741 = n17740 ^ n15341;
  assign n17726 = n17725 ^ n17721;
  assign n17695 = n17694 ^ n17688;
  assign n17715 = n17695 ^ n15378;
  assign n17683 = n17682 ^ n17646;
  assign n17684 = ~n17647 & ~n17683;
  assign n17685 = n17684 ^ n15349;
  assign n17716 = n17695 ^ n17685;
  assign n17717 = n17715 & n17716;
  assign n17718 = n17717 ^ n15378;
  assign n17727 = n17726 ^ n17718;
  assign n17730 = n17726 ^ n15347;
  assign n17731 = ~n17727 & n17730;
  assign n17732 = n17731 ^ n15347;
  assign n17800 = n17740 ^ n17732;
  assign n17801 = n17741 & n17800;
  assign n17802 = n17801 ^ n15341;
  assign n17941 = n17811 ^ n17802;
  assign n17942 = n17812 & n17941;
  assign n17943 = n17942 ^ n15391;
  assign n17945 = n17944 ^ n17943;
  assign n17946 = n17944 ^ n15337;
  assign n17947 = n17945 & n17946;
  assign n17948 = n17947 ^ n15337;
  assign n17949 = n17948 ^ n17939;
  assign n17950 = n17940 & n17949;
  assign n17951 = n17950 ^ n15401;
  assign n17952 = n17951 ^ n17937;
  assign n17953 = ~n17938 & n17952;
  assign n17954 = n17953 ^ n14826;
  assign n17955 = n17954 ^ n17934;
  assign n17956 = ~n17935 & ~n17955;
  assign n17957 = n17956 ^ n15330;
  assign n17959 = n17958 ^ n17957;
  assign n17960 = n17958 ^ n15414;
  assign n17961 = ~n17959 & ~n17960;
  assign n17962 = n17961 ^ n15414;
  assign n17963 = n17962 ^ n17932;
  assign n17964 = ~n17933 & n17963;
  assign n17965 = n17964 ^ n15423;
  assign n17967 = n17966 ^ n17965;
  assign n17968 = n17966 ^ n15501;
  assign n17969 = ~n17967 & n17968;
  assign n17970 = n17969 ^ n15501;
  assign n17972 = n17971 ^ n17970;
  assign n17973 = n17971 ^ n15543;
  assign n17974 = n17972 & n17973;
  assign n17975 = n17974 ^ n15543;
  assign n17976 = n17975 ^ n17930;
  assign n17977 = ~n17931 & n17976;
  assign n17978 = n17977 ^ n15558;
  assign n17979 = n17978 ^ n17928;
  assign n17980 = n17929 & ~n17979;
  assign n17981 = n17980 ^ n15672;
  assign n17982 = n17981 ^ n17926;
  assign n17983 = n17927 & n17982;
  assign n17984 = n17983 ^ n15692;
  assign n17985 = n17984 ^ n17924;
  assign n17986 = n17925 & n17985;
  assign n17987 = n17986 ^ n15726;
  assign n17988 = n17987 ^ n17921;
  assign n17989 = n17922 & ~n17988;
  assign n17990 = n17989 ^ n15761;
  assign n17999 = n17998 ^ n17990;
  assign n18000 = n17998 ^ n15128;
  assign n18001 = n17999 & ~n18000;
  assign n18002 = n18001 ^ n15128;
  assign n18012 = n18011 ^ n18002;
  assign n18138 = n18011 ^ n15133;
  assign n18139 = n18012 & ~n18138;
  assign n18140 = n18139 ^ n15133;
  assign n18150 = n18149 ^ n18140;
  assign n18013 = n18012 ^ n15133;
  assign n18014 = n17987 ^ n17922;
  assign n18015 = n17984 ^ n17925;
  assign n18016 = n17981 ^ n17927;
  assign n18017 = n17975 ^ n17931;
  assign n18018 = n17967 ^ n15501;
  assign n18019 = n17962 ^ n17933;
  assign n18020 = n17948 ^ n15401;
  assign n18021 = n18020 ^ n17939;
  assign n18022 = n17945 ^ n15337;
  assign n17813 = n17812 ^ n17802;
  assign n17686 = n17685 ^ n15378;
  assign n17696 = n17695 ^ n17686;
  assign n17713 = n17697 & ~n17712;
  assign n17714 = n17696 & n17713;
  assign n17728 = n17727 ^ n15347;
  assign n17729 = n17714 & ~n17728;
  assign n17742 = n17741 ^ n17732;
  assign n17814 = ~n17729 & n17742;
  assign n18023 = n17813 & ~n17814;
  assign n18024 = n18022 & ~n18023;
  assign n18025 = n18021 & ~n18024;
  assign n18026 = n17951 ^ n14826;
  assign n18027 = n18026 ^ n17937;
  assign n18028 = n18025 & n18027;
  assign n18029 = n17954 ^ n15330;
  assign n18030 = n18029 ^ n17934;
  assign n18031 = n18028 & n18030;
  assign n18032 = n17959 ^ n15414;
  assign n18033 = n18031 & ~n18032;
  assign n18034 = ~n18019 & ~n18033;
  assign n18035 = n18018 & n18034;
  assign n18036 = n17972 ^ n15543;
  assign n18037 = ~n18035 & ~n18036;
  assign n18038 = ~n18017 & n18037;
  assign n18039 = n17978 ^ n15672;
  assign n18040 = n18039 ^ n17928;
  assign n18041 = ~n18038 & ~n18040;
  assign n18042 = n18016 & ~n18041;
  assign n18043 = ~n18015 & n18042;
  assign n18044 = ~n18014 & ~n18043;
  assign n18045 = n17999 ^ n15128;
  assign n18046 = ~n18044 & ~n18045;
  assign n18137 = ~n18013 & n18046;
  assign n18151 = n18150 ^ n18137;
  assign n18047 = n18046 ^ n18013;
  assign n2304 = n2271 ^ x358;
  assign n2305 = n2304 ^ n1335;
  assign n2306 = n2305 ^ x294;
  assign n18048 = n18047 ^ n2306;
  assign n18049 = n18045 ^ n18044;
  assign n18050 = n18049 ^ n1328;
  assign n18051 = n18043 ^ n18014;
  assign n1150 = n1055 ^ x360;
  assign n1151 = n1150 ^ n1144;
  assign n1152 = n1151 ^ x296;
  assign n18052 = n18051 ^ n1152;
  assign n18053 = n18042 ^ n18015;
  assign n18054 = n18053 ^ n1137;
  assign n18120 = n18041 ^ n18016;
  assign n18055 = n18040 ^ n18038;
  assign n18056 = n18055 ^ n994;
  assign n18057 = n18037 ^ n18017;
  assign n18058 = n18057 ^ n988;
  assign n18059 = n18036 ^ n18035;
  assign n18060 = n18059 ^ n713;
  assign n18103 = n18034 ^ n18018;
  assign n18061 = n18033 ^ n18019;
  assign n18062 = n18061 ^ n549;
  assign n18063 = n18032 ^ n18031;
  assign n18064 = n18063 ^ n643;
  assign n18065 = n18030 ^ n18028;
  assign n18066 = n18065 ^ n634;
  assign n18067 = n18027 ^ n18025;
  assign n18071 = n18070 ^ n18067;
  assign n18072 = n18024 ^ n18021;
  assign n18076 = n18075 ^ n18072;
  assign n18077 = n18023 ^ n18022;
  assign n18081 = n18080 ^ n18077;
  assign n17815 = n17814 ^ n17813;
  assign n17819 = n17818 ^ n17815;
  assign n17743 = n17742 ^ n17729;
  assign n17744 = n17743 ^ n2156;
  assign n17745 = n17728 ^ n17714;
  assign n17746 = n17745 ^ n2138;
  assign n17747 = n17713 ^ n17696;
  assign n17748 = n17747 ^ n1901;
  assign n17788 = n17786 ^ n2118;
  assign n17789 = ~n17787 & n17788;
  assign n17790 = n17789 ^ n2118;
  assign n17791 = n17790 ^ n17747;
  assign n17792 = ~n17748 & n17791;
  assign n17793 = n17792 ^ n1901;
  assign n17794 = n17793 ^ n17745;
  assign n17795 = n17746 & ~n17794;
  assign n17796 = n17795 ^ n2138;
  assign n17797 = n17796 ^ n17743;
  assign n17798 = ~n17744 & n17797;
  assign n17799 = n17798 ^ n2156;
  assign n18082 = n17815 ^ n17799;
  assign n18083 = n17819 & ~n18082;
  assign n18084 = n18083 ^ n17818;
  assign n18085 = n18084 ^ n18077;
  assign n18086 = ~n18081 & n18085;
  assign n18087 = n18086 ^ n18080;
  assign n18088 = n18087 ^ n18072;
  assign n18089 = n18076 & ~n18088;
  assign n18090 = n18089 ^ n18075;
  assign n18091 = n18090 ^ n18067;
  assign n18092 = ~n18071 & n18091;
  assign n18093 = n18092 ^ n18070;
  assign n18094 = n18093 ^ n18065;
  assign n18095 = ~n18066 & n18094;
  assign n18096 = n18095 ^ n634;
  assign n18097 = n18096 ^ n18063;
  assign n18098 = n18064 & ~n18097;
  assign n18099 = n18098 ^ n643;
  assign n18100 = n18099 ^ n18061;
  assign n18101 = n18062 & ~n18100;
  assign n18102 = n18101 ^ n549;
  assign n18104 = n18103 ^ n18102;
  assign n18108 = n18107 ^ n18103;
  assign n18109 = ~n18104 & n18108;
  assign n18110 = n18109 ^ n18107;
  assign n18111 = n18110 ^ n18059;
  assign n18112 = ~n18060 & n18111;
  assign n18113 = n18112 ^ n713;
  assign n18114 = n18113 ^ n18057;
  assign n18115 = n18058 & ~n18114;
  assign n18116 = n18115 ^ n988;
  assign n18117 = n18116 ^ n18055;
  assign n18118 = n18056 & ~n18117;
  assign n18119 = n18118 ^ n994;
  assign n18121 = n18120 ^ n18119;
  assign n18122 = n18120 ^ n1009;
  assign n18123 = ~n18121 & n18122;
  assign n18124 = n18123 ^ n1009;
  assign n18125 = n18124 ^ n18053;
  assign n18126 = n18054 & ~n18125;
  assign n18127 = n18126 ^ n1137;
  assign n18128 = n18127 ^ n18051;
  assign n18129 = n18052 & ~n18128;
  assign n18130 = n18129 ^ n1152;
  assign n18131 = n18130 ^ n18049;
  assign n18132 = ~n18050 & n18131;
  assign n18133 = n18132 ^ n1328;
  assign n18134 = n18133 ^ n18047;
  assign n18135 = n18048 & ~n18134;
  assign n18136 = n18135 ^ n2306;
  assign n18152 = n18151 ^ n18136;
  assign n18215 = n18152 ^ n2323;
  assign n18264 = n18217 ^ n18215;
  assign n18291 = n18264 ^ n15322;
  assign n18360 = n18291 & n18359;
  assign n18361 = n18360 ^ n1433;
  assign n18170 = n18137 & n18150;
  assign n18165 = n17560 ^ n1042;
  assign n18163 = n16908 ^ n16413;
  assign n18164 = n18163 ^ n15738;
  assign n18166 = n18165 ^ n18164;
  assign n18159 = n18147 ^ n18145;
  assign n18160 = n18147 ^ n18143;
  assign n18161 = n18159 & ~n18160;
  assign n18162 = n18161 ^ n18145;
  assign n18167 = n18166 ^ n18162;
  assign n18168 = n18167 ^ n15145;
  assign n18156 = n18148 ^ n18140;
  assign n18157 = n18149 & ~n18156;
  assign n18158 = n18157 ^ n15137;
  assign n18169 = n18168 ^ n18158;
  assign n18171 = n18170 ^ n18169;
  assign n18153 = n18151 ^ n2323;
  assign n18154 = n18152 & ~n18153;
  assign n18155 = n18154 ^ n2323;
  assign n18172 = n18171 ^ n18155;
  assign n2418 = n2351 ^ x356;
  assign n2419 = n2418 ^ n2414;
  assign n2420 = n2419 ^ x292;
  assign n18220 = n18172 ^ n2420;
  assign n18218 = ~n18215 & n18217;
  assign n18213 = n16925 ^ n16162;
  assign n18214 = n18213 ^ n17017;
  assign n18219 = n18218 ^ n18214;
  assign n18267 = n18220 ^ n18219;
  assign n18265 = n15322 & ~n18264;
  assign n18266 = n18265 ^ n15317;
  assign n18292 = n18267 ^ n18266;
  assign n18362 = n18292 ^ n18291;
  assign n18363 = n18362 ^ n18360;
  assign n18364 = n18361 & n18363;
  assign n18365 = n18364 ^ n1433;
  assign n18961 = n18370 ^ n18365;
  assign n18268 = n18267 ^ n18265;
  assign n18269 = n18266 & ~n18268;
  assign n18270 = n18269 ^ n15317;
  assign n18226 = n16937 ^ n16158;
  assign n18227 = n18226 ^ n17644;
  assign n18185 = n17565 ^ n17564;
  assign n18182 = n18165 ^ n18162;
  assign n18183 = n18166 & ~n18182;
  assign n18184 = n18183 ^ n18164;
  assign n18186 = n18185 ^ n18184;
  assign n18180 = n17100 ^ n16409;
  assign n18181 = n18180 ^ n15766;
  assign n18187 = n18186 ^ n18181;
  assign n18188 = n18187 ^ n15122;
  assign n18177 = n18167 ^ n18158;
  assign n18178 = ~n18168 & ~n18177;
  assign n18179 = n18178 ^ n15145;
  assign n18189 = n18188 ^ n18179;
  assign n18176 = n18169 & ~n18170;
  assign n18190 = n18189 ^ n18176;
  assign n18173 = n18171 ^ n2420;
  assign n18174 = n18172 & ~n18173;
  assign n18175 = n18174 ^ n2420;
  assign n18191 = n18190 ^ n18175;
  assign n1542 = n1541 ^ x355;
  assign n1543 = n1542 ^ n1511;
  assign n1544 = n1543 ^ x291;
  assign n18224 = n18191 ^ n1544;
  assign n18221 = n18220 ^ n18214;
  assign n18222 = ~n18219 & ~n18221;
  assign n18223 = n18222 ^ n18218;
  assign n18225 = n18224 ^ n18223;
  assign n18262 = n18227 ^ n18225;
  assign n18263 = n18262 ^ n15316;
  assign n18294 = n18270 ^ n18263;
  assign n18293 = ~n18291 & n18292;
  assign n18366 = n18294 ^ n18293;
  assign n18962 = n18961 ^ n18366;
  assign n18965 = n18964 ^ n18962;
  assign n18968 = n18362 ^ n18361;
  assign n18439 = n17782 ^ n17750;
  assign n18966 = n18439 ^ n17002;
  assign n18967 = n18966 ^ n17872;
  assign n18969 = n18968 ^ n18967;
  assign n18999 = n18359 ^ n18291;
  assign n18985 = n17605 ^ n17025;
  assign n18986 = n18985 ^ n16170;
  assign n18984 = n18133 ^ n18048;
  assign n18987 = n18986 ^ n18984;
  assign n18883 = n18130 ^ n18050;
  assign n18834 = n18127 ^ n18052;
  assign n18831 = n17089 ^ n16409;
  assign n18832 = n18831 ^ n17612;
  assign n18879 = n18834 ^ n18832;
  assign n18801 = n17623 ^ n16413;
  assign n18802 = n18801 ^ n17093;
  assign n18800 = n18124 ^ n18054;
  assign n18803 = n18802 ^ n18800;
  assign n18775 = n18121 ^ n1009;
  assign n18658 = n18116 ^ n18056;
  assign n18249 = n17571 ^ n17427;
  assign n18656 = n18249 ^ n16423;
  assign n18657 = n18656 ^ n16908;
  assign n18659 = n18658 ^ n18657;
  assign n18643 = n18113 ^ n988;
  assign n18644 = n18643 ^ n18057;
  assign n18629 = n18110 ^ n18060;
  assign n18627 = n18185 ^ n17599;
  assign n18628 = n18627 ^ n16943;
  assign n18630 = n18629 ^ n18628;
  assign n18615 = n18107 ^ n18104;
  assign n18613 = n18165 ^ n16949;
  assign n18614 = n18613 ^ n17349;
  assign n18616 = n18615 ^ n18614;
  assign n18601 = n18099 ^ n18062;
  assign n18586 = n18096 ^ n18064;
  assign n18584 = n18009 ^ n16901;
  assign n18585 = n18584 ^ n17184;
  assign n18587 = n18586 ^ n18585;
  assign n18549 = n18093 ^ n18066;
  assign n18546 = n17996 ^ n16941;
  assign n18547 = n18546 ^ n16670;
  assign n18580 = n18549 ^ n18547;
  assign n18423 = n17832 ^ n16958;
  assign n18424 = n18423 ^ n16096;
  assign n18422 = n18084 ^ n18081;
  assign n18425 = n18424 ^ n18422;
  assign n18426 = n17836 ^ n16097;
  assign n18427 = n18426 ^ n16962;
  assign n17820 = n17819 ^ n17799;
  assign n18428 = n18427 ^ n17820;
  assign n18432 = n17850 ^ n16975;
  assign n18433 = n18432 ^ n16112;
  assign n18431 = n17790 ^ n17748;
  assign n18434 = n18433 ^ n18431;
  assign n18436 = n16979 ^ n16117;
  assign n18437 = n18436 ^ n17891;
  assign n18438 = n18437 ^ n18435;
  assign n18443 = n17779 ^ n1657;
  assign n18444 = n18443 ^ n17751;
  assign n18403 = n17776 ^ n17754;
  assign n18401 = n17860 ^ n16135;
  assign n18402 = n18401 ^ n16992;
  assign n18404 = n18403 ^ n18402;
  assign n18338 = n17773 ^ n1583;
  assign n18339 = n18338 ^ n17755;
  assign n18323 = n17862 ^ n16998;
  assign n18324 = n18323 ^ n16144;
  assign n18321 = n17770 ^ n1574;
  assign n18322 = n18321 ^ n17757;
  assign n18325 = n18324 ^ n18322;
  assign n18286 = n17764 ^ n17700;
  assign n18283 = n17736 ^ n16152;
  assign n18284 = n18283 ^ n17135;
  assign n18306 = n18286 ^ n18284;
  assign n18203 = n17568 ^ n17432;
  assign n18201 = n17093 ^ n15770;
  assign n18202 = n18201 ^ n16174;
  assign n18204 = n18203 ^ n18202;
  assign n18198 = n18185 ^ n18181;
  assign n18199 = ~n18186 & ~n18198;
  assign n18200 = n18199 ^ n18181;
  assign n18205 = n18204 ^ n18200;
  assign n18195 = n18187 ^ n18179;
  assign n18196 = ~n18188 & ~n18195;
  assign n18197 = n18196 ^ n15122;
  assign n18206 = n18205 ^ n18197;
  assign n18207 = n18206 ^ n14835;
  assign n18208 = ~n18176 & n18189;
  assign n18254 = ~n18207 & n18208;
  assign n18247 = n17089 ^ n16170;
  assign n18248 = n18247 ^ n15323;
  assign n18250 = n18249 ^ n18248;
  assign n18244 = n18203 ^ n18200;
  assign n18245 = ~n18204 & n18244;
  assign n18246 = n18245 ^ n18202;
  assign n18251 = n18250 ^ n18246;
  assign n18252 = n18251 ^ n14831;
  assign n18241 = n18205 ^ n14835;
  assign n18242 = ~n18206 & ~n18241;
  assign n18243 = n18242 ^ n14835;
  assign n18253 = n18252 ^ n18243;
  assign n18255 = n18254 ^ n18253;
  assign n18209 = n18208 ^ n18207;
  assign n18192 = n18190 ^ n1544;
  assign n18193 = ~n18191 & n18192;
  assign n18194 = n18193 ^ n1544;
  assign n18210 = n18209 ^ n18194;
  assign n18234 = n18209 ^ n2561;
  assign n18235 = ~n18210 & n18234;
  assign n18236 = n18235 ^ n2561;
  assign n18240 = n18239 ^ n18236;
  assign n18256 = n18255 ^ n18240;
  assign n18211 = n18210 ^ n2561;
  assign n17826 = n17690 ^ n16932;
  assign n17827 = n17826 ^ n16154;
  assign n18212 = n18211 ^ n17827;
  assign n18228 = n18227 ^ n18224;
  assign n18229 = ~n18225 & ~n18228;
  assign n18230 = n18229 ^ n18227;
  assign n18231 = n18230 ^ n18211;
  assign n18232 = n18212 & n18231;
  assign n18233 = n18232 ^ n17827;
  assign n18257 = n18256 ^ n18233;
  assign n17824 = n16927 ^ n16458;
  assign n17825 = n17824 ^ n17722;
  assign n18280 = n18256 ^ n17825;
  assign n18281 = ~n18257 & ~n18280;
  assign n18282 = n18281 ^ n17825;
  assign n18307 = n18286 ^ n18282;
  assign n18308 = n18306 & ~n18307;
  assign n18309 = n18308 ^ n18284;
  assign n18305 = n17767 ^ n17766;
  assign n18310 = n18309 ^ n18305;
  assign n18303 = n17807 ^ n16148;
  assign n18304 = n18303 ^ n17002;
  assign n18318 = n18305 ^ n18304;
  assign n18319 = ~n18310 & ~n18318;
  assign n18320 = n18319 ^ n18304;
  assign n18335 = n18322 ^ n18320;
  assign n18336 = n18325 & ~n18335;
  assign n18337 = n18336 ^ n18324;
  assign n18340 = n18339 ^ n18337;
  assign n18333 = n16994 ^ n16140;
  assign n18334 = n18333 ^ n17872;
  assign n18398 = n18339 ^ n18334;
  assign n18399 = n18340 & ~n18398;
  assign n18400 = n18399 ^ n18334;
  assign n18440 = n18403 ^ n18400;
  assign n18441 = n18404 & n18440;
  assign n18442 = n18441 ^ n18402;
  assign n18445 = n18444 ^ n18442;
  assign n18446 = n17854 ^ n16127;
  assign n18447 = n18446 ^ n16986;
  assign n18448 = n18447 ^ n18444;
  assign n18449 = n18445 & ~n18448;
  assign n18450 = n18449 ^ n18447;
  assign n18451 = n18450 ^ n18439;
  assign n18452 = n16982 ^ n16122;
  assign n18453 = n18452 ^ n17822;
  assign n18454 = n18453 ^ n18439;
  assign n18455 = ~n18451 & ~n18454;
  assign n18456 = n18455 ^ n18453;
  assign n18457 = n18456 ^ n18435;
  assign n18458 = ~n18438 & ~n18457;
  assign n18459 = n18458 ^ n18437;
  assign n18460 = n18459 ^ n18433;
  assign n18461 = n18434 & ~n18460;
  assign n18462 = n18461 ^ n18431;
  assign n18429 = n17793 ^ n2138;
  assign n18430 = n18429 ^ n17745;
  assign n18463 = n18462 ^ n18430;
  assign n18464 = n17848 ^ n16969;
  assign n18465 = n18464 ^ n16107;
  assign n18466 = n18465 ^ n18430;
  assign n18467 = n18463 & n18466;
  assign n18468 = n18467 ^ n18465;
  assign n18414 = n17796 ^ n17744;
  assign n18469 = n18468 ^ n18414;
  assign n18470 = n17841 ^ n16102;
  assign n18471 = n18470 ^ n16967;
  assign n18472 = n18471 ^ n18414;
  assign n18473 = n18469 & ~n18472;
  assign n18474 = n18473 ^ n18471;
  assign n18475 = n18474 ^ n18427;
  assign n18476 = n18428 & ~n18475;
  assign n18477 = n18476 ^ n17820;
  assign n18478 = n18477 ^ n18422;
  assign n18479 = ~n18425 & n18478;
  assign n18480 = n18479 ^ n18424;
  assign n18421 = n18087 ^ n18076;
  assign n18481 = n18480 ^ n18421;
  assign n18419 = n16952 ^ n16511;
  assign n18420 = n18419 ^ n17828;
  assign n18534 = n18421 ^ n18420;
  assign n18535 = ~n18481 & n18534;
  assign n18536 = n18535 ^ n18420;
  assign n18533 = n18090 ^ n18071;
  assign n18537 = n18536 ^ n18533;
  assign n18531 = n16947 ^ n16655;
  assign n18532 = n18531 ^ n17919;
  assign n18543 = n18533 ^ n18532;
  assign n18544 = n18537 & n18543;
  assign n18545 = n18544 ^ n18532;
  assign n18581 = n18549 ^ n18545;
  assign n18582 = n18580 & ~n18581;
  assign n18583 = n18582 ^ n18547;
  assign n18598 = n18586 ^ n18583;
  assign n18599 = ~n18587 & n18598;
  assign n18600 = n18599 ^ n18585;
  assign n18602 = n18601 ^ n18600;
  assign n18596 = n17341 ^ n16955;
  assign n18597 = n18596 ^ n18147;
  assign n18610 = n18601 ^ n18597;
  assign n18611 = n18602 & ~n18610;
  assign n18612 = n18611 ^ n18597;
  assign n18624 = n18614 ^ n18612;
  assign n18625 = n18616 & n18624;
  assign n18626 = n18625 ^ n18615;
  assign n18640 = n18629 ^ n18626;
  assign n18641 = n18630 & n18640;
  assign n18642 = n18641 ^ n18628;
  assign n18645 = n18644 ^ n18642;
  assign n18638 = n18203 ^ n16418;
  assign n18639 = n18638 ^ n16913;
  assign n18653 = n18644 ^ n18639;
  assign n18654 = n18645 & ~n18653;
  assign n18655 = n18654 ^ n18639;
  assign n18772 = n18658 ^ n18655;
  assign n18773 = ~n18659 & n18772;
  assign n18774 = n18773 ^ n18657;
  assign n18776 = n18775 ^ n18774;
  assign n18770 = n17618 ^ n16430;
  assign n18771 = n18770 ^ n17100;
  assign n18797 = n18775 ^ n18771;
  assign n18798 = n18776 & ~n18797;
  assign n18799 = n18798 ^ n18771;
  assign n18828 = n18802 ^ n18799;
  assign n18829 = ~n18803 & ~n18828;
  assign n18830 = n18829 ^ n18800;
  assign n18880 = n18834 ^ n18830;
  assign n18881 = n18879 & ~n18880;
  assign n18882 = n18881 ^ n18832;
  assign n18884 = n18883 ^ n18882;
  assign n18877 = n17609 ^ n17031;
  assign n18878 = n18877 ^ n16174;
  assign n18981 = n18883 ^ n18878;
  assign n18982 = n18884 & ~n18981;
  assign n18983 = n18982 ^ n18878;
  assign n18988 = n18987 ^ n18983;
  assign n18885 = n18884 ^ n18878;
  assign n18886 = n18885 ^ n15770;
  assign n18833 = n18832 ^ n18830;
  assign n18835 = n18834 ^ n18833;
  assign n18836 = n18835 ^ n15766;
  assign n18804 = n18803 ^ n18799;
  assign n18777 = n18776 ^ n18771;
  assign n18778 = n18777 ^ n15701;
  assign n18660 = n18659 ^ n18655;
  assign n18661 = n18660 ^ n15712;
  assign n18646 = n18645 ^ n18639;
  assign n18647 = n18646 ^ n15707;
  assign n18631 = n18630 ^ n18626;
  assign n18632 = n18631 ^ n16397;
  assign n18617 = n18616 ^ n18612;
  assign n18618 = n18617 ^ n16180;
  assign n18603 = n18602 ^ n18597;
  assign n18606 = n18603 ^ n16184;
  assign n18588 = n18587 ^ n18583;
  assign n18591 = n18588 ^ n16099;
  assign n18548 = n18547 ^ n18545;
  assign n18550 = n18549 ^ n18548;
  assign n18538 = n18537 ^ n18532;
  assign n18482 = n18481 ^ n18420;
  assign n18483 = n18482 ^ n16114;
  assign n18484 = n18477 ^ n18425;
  assign n18485 = n18484 ^ n16119;
  assign n18486 = n18474 ^ n18428;
  assign n18487 = n18486 ^ n16124;
  assign n18488 = n18471 ^ n18469;
  assign n18489 = n18488 ^ n16129;
  assign n18490 = n18465 ^ n18463;
  assign n18491 = n18490 ^ n16133;
  assign n18492 = n18459 ^ n18434;
  assign n18493 = n18492 ^ n16138;
  assign n18494 = n18456 ^ n18437;
  assign n18495 = n18494 ^ n18435;
  assign n18496 = n18495 ^ n16089;
  assign n18497 = n18453 ^ n18451;
  assign n18498 = n18497 ^ n16069;
  assign n18502 = n18447 ^ n18445;
  assign n18405 = n18404 ^ n18400;
  assign n18406 = n18405 ^ n15831;
  assign n18341 = n18340 ^ n18334;
  assign n18342 = n18341 ^ n15310;
  assign n18326 = n18325 ^ n18320;
  assign n18327 = n18326 ^ n15311;
  assign n18311 = n18310 ^ n18304;
  assign n18312 = n18311 ^ n15312;
  assign n18285 = n18284 ^ n18282;
  assign n18287 = n18286 ^ n18285;
  assign n18258 = n18257 ^ n17825;
  assign n18259 = n18258 ^ n15314;
  assign n18260 = n18230 ^ n18212;
  assign n18261 = n18260 ^ n15315;
  assign n18271 = n18270 ^ n18262;
  assign n18272 = ~n18263 & n18271;
  assign n18273 = n18272 ^ n15316;
  assign n18274 = n18273 ^ n18260;
  assign n18275 = n18261 & n18274;
  assign n18276 = n18275 ^ n15315;
  assign n18277 = n18276 ^ n18258;
  assign n18278 = ~n18259 & ~n18277;
  assign n18279 = n18278 ^ n15314;
  assign n18288 = n18287 ^ n18279;
  assign n18300 = n18287 ^ n15313;
  assign n18301 = n18288 & ~n18300;
  assign n18302 = n18301 ^ n15313;
  assign n18315 = n18311 ^ n18302;
  assign n18316 = ~n18312 & ~n18315;
  assign n18317 = n18316 ^ n15312;
  assign n18330 = n18326 ^ n18317;
  assign n18331 = ~n18327 & n18330;
  assign n18332 = n18331 ^ n15311;
  assign n18395 = n18341 ^ n18332;
  assign n18396 = n18342 & ~n18395;
  assign n18397 = n18396 ^ n15310;
  assign n18499 = n18405 ^ n18397;
  assign n18500 = ~n18406 & n18499;
  assign n18501 = n18500 ^ n15831;
  assign n18503 = n18502 ^ n18501;
  assign n18504 = n18502 ^ n15918;
  assign n18505 = n18503 & n18504;
  assign n18506 = n18505 ^ n15918;
  assign n18507 = n18506 ^ n18497;
  assign n18508 = ~n18498 & ~n18507;
  assign n18509 = n18508 ^ n16069;
  assign n18510 = n18509 ^ n18495;
  assign n18511 = ~n18496 & ~n18510;
  assign n18512 = n18511 ^ n16089;
  assign n18513 = n18512 ^ n18492;
  assign n18514 = n18493 & n18513;
  assign n18515 = n18514 ^ n16138;
  assign n18516 = n18515 ^ n18490;
  assign n18517 = ~n18491 & ~n18516;
  assign n18518 = n18517 ^ n16133;
  assign n18519 = n18518 ^ n18488;
  assign n18520 = ~n18489 & n18519;
  assign n18521 = n18520 ^ n16129;
  assign n18522 = n18521 ^ n18486;
  assign n18523 = ~n18487 & ~n18522;
  assign n18524 = n18523 ^ n16124;
  assign n18525 = n18524 ^ n18484;
  assign n18526 = ~n18485 & ~n18525;
  assign n18527 = n18526 ^ n16119;
  assign n18528 = n18527 ^ n18482;
  assign n18529 = ~n18483 & ~n18528;
  assign n18530 = n18529 ^ n16114;
  assign n18539 = n18538 ^ n18530;
  assign n18540 = n18538 ^ n16109;
  assign n18541 = n18539 & ~n18540;
  assign n18542 = n18541 ^ n16109;
  assign n18551 = n18550 ^ n18542;
  assign n18576 = n18550 ^ n16104;
  assign n18577 = ~n18551 & n18576;
  assign n18578 = n18577 ^ n16104;
  assign n18592 = n18588 ^ n18578;
  assign n18593 = ~n18591 & n18592;
  assign n18594 = n18593 ^ n16099;
  assign n18607 = n18603 ^ n18594;
  assign n18608 = n18606 & n18607;
  assign n18609 = n18608 ^ n16184;
  assign n18621 = n18617 ^ n18609;
  assign n18622 = ~n18618 & n18621;
  assign n18623 = n18622 ^ n16180;
  assign n18635 = n18631 ^ n18623;
  assign n18636 = ~n18632 & ~n18635;
  assign n18637 = n18636 ^ n16397;
  assign n18650 = n18646 ^ n18637;
  assign n18651 = ~n18647 & n18650;
  assign n18652 = n18651 ^ n15707;
  assign n18767 = n18660 ^ n18652;
  assign n18768 = ~n18661 & n18767;
  assign n18769 = n18768 ^ n15712;
  assign n18794 = n18777 ^ n18769;
  assign n18795 = ~n18778 & n18794;
  assign n18796 = n18795 ^ n15701;
  assign n18805 = n18804 ^ n18796;
  assign n18825 = n18804 ^ n15738;
  assign n18826 = n18805 & n18825;
  assign n18827 = n18826 ^ n15738;
  assign n18874 = n18835 ^ n18827;
  assign n18875 = n18836 & ~n18874;
  assign n18876 = n18875 ^ n15766;
  assign n18977 = n18885 ^ n18876;
  assign n18978 = ~n18886 & n18977;
  assign n18979 = n18978 ^ n15770;
  assign n18980 = n18979 ^ n15323;
  assign n18989 = n18988 ^ n18980;
  assign n18887 = n18886 ^ n18876;
  assign n18552 = n18551 ^ n16104;
  assign n18553 = n18524 ^ n18485;
  assign n18554 = n18521 ^ n18487;
  assign n18555 = n18506 ^ n18498;
  assign n18289 = n18288 ^ n15313;
  assign n18290 = n18276 ^ n18259;
  assign n18295 = n18293 & ~n18294;
  assign n18296 = n18273 ^ n18261;
  assign n18297 = n18295 & n18296;
  assign n18298 = n18290 & n18297;
  assign n18299 = n18289 & ~n18298;
  assign n18313 = n18312 ^ n18302;
  assign n18314 = ~n18299 & ~n18313;
  assign n18328 = n18327 ^ n18317;
  assign n18329 = ~n18314 & ~n18328;
  assign n18343 = n18342 ^ n18332;
  assign n18394 = n18329 & n18343;
  assign n18407 = n18406 ^ n18397;
  assign n18556 = n18394 & ~n18407;
  assign n18557 = n18503 ^ n15918;
  assign n18558 = ~n18556 & ~n18557;
  assign n18559 = n18555 & ~n18558;
  assign n18560 = n18509 ^ n18496;
  assign n18561 = ~n18559 & n18560;
  assign n18562 = n18512 ^ n18493;
  assign n18563 = ~n18561 & ~n18562;
  assign n18564 = n18515 ^ n18491;
  assign n18565 = n18563 & ~n18564;
  assign n18566 = n18518 ^ n18489;
  assign n18567 = n18565 & n18566;
  assign n18568 = n18554 & n18567;
  assign n18569 = n18553 & ~n18568;
  assign n18570 = n18527 ^ n16114;
  assign n18571 = n18570 ^ n18482;
  assign n18572 = n18569 & ~n18571;
  assign n18573 = n18539 ^ n16109;
  assign n18574 = ~n18572 & ~n18573;
  assign n18575 = n18552 & n18574;
  assign n18579 = n18578 ^ n16099;
  assign n18589 = n18588 ^ n18579;
  assign n18590 = ~n18575 & n18589;
  assign n18595 = n18594 ^ n16184;
  assign n18604 = n18603 ^ n18595;
  assign n18605 = ~n18590 & n18604;
  assign n18619 = n18618 ^ n18609;
  assign n18620 = n18605 & n18619;
  assign n18633 = n18632 ^ n18623;
  assign n18634 = ~n18620 & ~n18633;
  assign n18648 = n18647 ^ n18637;
  assign n18649 = ~n18634 & ~n18648;
  assign n18662 = n18661 ^ n18652;
  assign n18766 = n18649 & ~n18662;
  assign n18779 = n18778 ^ n18769;
  assign n18793 = n18766 & ~n18779;
  assign n18806 = n18805 ^ n15738;
  assign n18824 = ~n18793 & ~n18806;
  assign n18837 = n18836 ^ n18827;
  assign n18888 = ~n18824 & ~n18837;
  assign n18976 = n18887 & n18888;
  assign n18990 = n18989 ^ n18976;
  assign n18991 = n18990 ^ n1520;
  assign n18889 = n18888 ^ n18887;
  assign n18838 = n18837 ^ n18824;
  assign n18807 = n18806 ^ n18793;
  assign n18820 = n18807 ^ n2401;
  assign n18780 = n18779 ^ n18766;
  assign n18781 = n18780 ^ n2388;
  assign n18663 = n18662 ^ n18649;
  assign n2377 = n1351 ^ x390;
  assign n2378 = n2377 ^ n2376;
  assign n2379 = n2378 ^ x326;
  assign n18664 = n18663 ^ n2379;
  assign n18665 = n18648 ^ n18634;
  assign n1296 = n1196 ^ x391;
  assign n1297 = n1296 ^ n1202;
  assign n1298 = n1297 ^ x327;
  assign n18666 = n18665 ^ n1298;
  assign n18667 = n18633 ^ n18620;
  assign n1278 = n1178 ^ x392;
  assign n1279 = n1278 ^ n1272;
  assign n1280 = n1279 ^ x328;
  assign n18668 = n18667 ^ n1280;
  assign n18669 = n18619 ^ n18605;
  assign n18670 = n18669 ^ n1028;
  assign n18671 = n18604 ^ n18590;
  assign n18672 = n18671 ^ n1262;
  assign n18673 = n18589 ^ n18575;
  assign n18674 = n18673 ^ n875;
  assign n18675 = n18574 ^ n18552;
  assign n18676 = n18675 ^ n772;
  assign n18677 = n18573 ^ n18572;
  assign n18678 = n18677 ^ n763;
  assign n18679 = n18571 ^ n18569;
  assign n18680 = n18679 ^ n698;
  assign n18734 = n18568 ^ n18553;
  assign n18681 = n18567 ^ n18554;
  assign n18685 = n18684 ^ n18681;
  assign n18686 = n18566 ^ n18565;
  assign n18690 = n18689 ^ n18686;
  assign n18691 = n18564 ^ n18563;
  assign n18695 = n18694 ^ n18691;
  assign n18696 = n18562 ^ n18561;
  assign n18700 = n18699 ^ n18696;
  assign n18701 = n18560 ^ n18559;
  assign n18702 = n18701 ^ n590;
  assign n18703 = n18558 ^ n18555;
  assign n18707 = n18706 ^ n18703;
  assign n18711 = n18557 ^ n18556;
  assign n18408 = n18407 ^ n18394;
  assign n18344 = n18343 ^ n18329;
  assign n18345 = n18344 ^ n1993;
  assign n18346 = n18328 ^ n18314;
  assign n18347 = n18346 ^ n1838;
  assign n18348 = n18313 ^ n18299;
  assign n18349 = n18348 ^ n1743;
  assign n18350 = n18298 ^ n18289;
  assign n18351 = n18350 ^ n1728;
  assign n18377 = n18297 ^ n18290;
  assign n18352 = n18296 ^ n18295;
  assign n18356 = n18355 ^ n18352;
  assign n18367 = n18366 ^ n18365;
  assign n18371 = n18370 ^ n18366;
  assign n18372 = n18367 & ~n18371;
  assign n18373 = n18372 ^ n18370;
  assign n18374 = n18373 ^ n18352;
  assign n18375 = n18356 & ~n18374;
  assign n18376 = n18375 ^ n18355;
  assign n18378 = n18377 ^ n18376;
  assign n18379 = n18377 ^ n1719;
  assign n18380 = ~n18378 & n18379;
  assign n18381 = n18380 ^ n1719;
  assign n18382 = n18381 ^ n18350;
  assign n18383 = n18351 & ~n18382;
  assign n18384 = n18383 ^ n1728;
  assign n18385 = n18384 ^ n18348;
  assign n18386 = n18349 & ~n18385;
  assign n18387 = n18386 ^ n1743;
  assign n18388 = n18387 ^ n18346;
  assign n18389 = ~n18347 & n18388;
  assign n18390 = n18389 ^ n1838;
  assign n18391 = n18390 ^ n18344;
  assign n18392 = ~n18345 & n18391;
  assign n18393 = n18392 ^ n1993;
  assign n18409 = n18408 ^ n18393;
  assign n18708 = n18408 ^ n1982;
  assign n18709 = ~n18409 & n18708;
  assign n18710 = n18709 ^ n1982;
  assign n18712 = n18711 ^ n18710;
  assign n18713 = n18711 ^ n2181;
  assign n18714 = ~n18712 & n18713;
  assign n18715 = n18714 ^ n2181;
  assign n18716 = n18715 ^ n18703;
  assign n18717 = n18707 & ~n18716;
  assign n18718 = n18717 ^ n18706;
  assign n18719 = n18718 ^ n18701;
  assign n18720 = ~n18702 & n18719;
  assign n18721 = n18720 ^ n590;
  assign n18722 = n18721 ^ n18696;
  assign n18723 = ~n18700 & n18722;
  assign n18724 = n18723 ^ n18699;
  assign n18725 = n18724 ^ n18691;
  assign n18726 = n18695 & ~n18725;
  assign n18727 = n18726 ^ n18694;
  assign n18728 = n18727 ^ n18686;
  assign n18729 = ~n18690 & n18728;
  assign n18730 = n18729 ^ n18689;
  assign n18731 = n18730 ^ n18681;
  assign n18732 = ~n18685 & n18731;
  assign n18733 = n18732 ^ n18684;
  assign n18735 = n18734 ^ n18733;
  assign n684 = n668 ^ x399;
  assign n688 = n687 ^ n684;
  assign n689 = n688 ^ x335;
  assign n18736 = n18734 ^ n689;
  assign n18737 = n18735 & ~n18736;
  assign n18738 = n18737 ^ n689;
  assign n18739 = n18738 ^ n18679;
  assign n18740 = ~n18680 & n18739;
  assign n18741 = n18740 ^ n698;
  assign n18742 = n18741 ^ n18677;
  assign n18743 = ~n18678 & n18742;
  assign n18744 = n18743 ^ n763;
  assign n18745 = n18744 ^ n18675;
  assign n18746 = ~n18676 & n18745;
  assign n18747 = n18746 ^ n772;
  assign n18748 = n18747 ^ n18673;
  assign n18749 = ~n18674 & n18748;
  assign n18750 = n18749 ^ n875;
  assign n18751 = n18750 ^ n18671;
  assign n18752 = n18672 & ~n18751;
  assign n18753 = n18752 ^ n1262;
  assign n18754 = n18753 ^ n18669;
  assign n18755 = ~n18670 & n18754;
  assign n18756 = n18755 ^ n1028;
  assign n18757 = n18756 ^ n1280;
  assign n18758 = n18668 & ~n18757;
  assign n18759 = n18758 ^ n18667;
  assign n18760 = n18759 ^ n18665;
  assign n18761 = ~n18666 & n18760;
  assign n18762 = n18761 ^ n1298;
  assign n18763 = n18762 ^ n18663;
  assign n18764 = n18664 & ~n18763;
  assign n18765 = n18764 ^ n2379;
  assign n18789 = n18765 ^ n2388;
  assign n18790 = n18781 & ~n18789;
  assign n18791 = n18790 ^ n18780;
  assign n18821 = n18807 ^ n18791;
  assign n18822 = n18820 & ~n18821;
  assign n18823 = n18822 ^ n2401;
  assign n18839 = n18838 ^ n18823;
  assign n18871 = n18838 ^ n2478;
  assign n18872 = n18839 & ~n18871;
  assign n18873 = n18872 ^ n2478;
  assign n18890 = n18889 ^ n18873;
  assign n2644 = n2566 ^ x386;
  assign n2645 = n2644 ^ n2471;
  assign n2646 = n2645 ^ x322;
  assign n18973 = n18889 ^ n2646;
  assign n18974 = n18890 & ~n18973;
  assign n18975 = n18974 ^ n2646;
  assign n18992 = n18991 ^ n18975;
  assign n18891 = n18890 ^ n2646;
  assign n18840 = n18839 ^ n2478;
  assign n18792 = n18791 ^ n2401;
  assign n18808 = n18807 ^ n18792;
  assign n18787 = n18305 ^ n17690;
  assign n18788 = n18787 ^ n17017;
  assign n18809 = n18808 ^ n18788;
  assign n18417 = n18286 ^ n17021;
  assign n18418 = n18417 ^ n17644;
  assign n18782 = n18781 ^ n18765;
  assign n18786 = n18418 & n18782;
  assign n18817 = n18788 ^ n18786;
  assign n18818 = n18809 & ~n18817;
  assign n18819 = n18818 ^ n18786;
  assign n18841 = n18840 ^ n18819;
  assign n18815 = n18322 ^ n16937;
  assign n18816 = n18815 ^ n17722;
  assign n18868 = n18840 ^ n18816;
  assign n18869 = n18841 & ~n18868;
  assign n18870 = n18869 ^ n18816;
  assign n18892 = n18891 ^ n18870;
  assign n18866 = n18339 ^ n16932;
  assign n18867 = n18866 ^ n17736;
  assign n18970 = n18891 ^ n18867;
  assign n18971 = n18892 & n18970;
  assign n18972 = n18971 ^ n18867;
  assign n18993 = n18992 ^ n18972;
  assign n18994 = n17807 ^ n16927;
  assign n18995 = n18994 ^ n18403;
  assign n18996 = n18995 ^ n18992;
  assign n18997 = ~n18993 & n18996;
  assign n18998 = n18997 ^ n18995;
  assign n19000 = n18999 ^ n18998;
  assign n19001 = n18444 ^ n17862;
  assign n19002 = n19001 ^ n17135;
  assign n19003 = n19002 ^ n18999;
  assign n19004 = n19000 & n19003;
  assign n19005 = n19004 ^ n19002;
  assign n19006 = n19005 ^ n18968;
  assign n19007 = n18969 & n19006;
  assign n19008 = n19007 ^ n18967;
  assign n19009 = n19008 ^ n18962;
  assign n19010 = ~n18965 & ~n19009;
  assign n19011 = n19010 ^ n18964;
  assign n18958 = n18431 ^ n17854;
  assign n18959 = n18958 ^ n16994;
  assign n18957 = n18373 ^ n18356;
  assign n18960 = n18959 ^ n18957;
  assign n19165 = n19011 ^ n18960;
  assign n19159 = n19008 ^ n18965;
  assign n19141 = n19002 ^ n19000;
  assign n19142 = n19141 ^ n16152;
  assign n19143 = n18995 ^ n18993;
  assign n19144 = n19143 ^ n16458;
  assign n18893 = n18892 ^ n18867;
  assign n18894 = n18893 ^ n16154;
  assign n18842 = n18841 ^ n18816;
  assign n18862 = n18842 ^ n16158;
  assign n18783 = n18782 ^ n18418;
  assign n18784 = n16166 & n18783;
  assign n18785 = n18784 ^ n16162;
  assign n18810 = n18809 ^ n18786;
  assign n18811 = n18810 ^ n18784;
  assign n18812 = ~n18785 & n18811;
  assign n18813 = n18812 ^ n16162;
  assign n18863 = n18842 ^ n18813;
  assign n18864 = ~n18862 & ~n18863;
  assign n18865 = n18864 ^ n16158;
  assign n19145 = n18893 ^ n18865;
  assign n19146 = n18894 & ~n19145;
  assign n19147 = n19146 ^ n16154;
  assign n19148 = n19147 ^ n19143;
  assign n19149 = n19144 & n19148;
  assign n19150 = n19149 ^ n16458;
  assign n19151 = n19150 ^ n19141;
  assign n19152 = n19142 & ~n19151;
  assign n19153 = n19152 ^ n16152;
  assign n19154 = n19153 ^ n16148;
  assign n19155 = n19005 ^ n18969;
  assign n19156 = n19155 ^ n19153;
  assign n19157 = ~n19154 & n19156;
  assign n19158 = n19157 ^ n16148;
  assign n19160 = n19159 ^ n19158;
  assign n19161 = n19159 ^ n16144;
  assign n19162 = ~n19160 & n19161;
  assign n19163 = n19162 ^ n16144;
  assign n19164 = n19163 ^ n16140;
  assign n19264 = n19165 ^ n19164;
  assign n19254 = n19147 ^ n19144;
  assign n18895 = n18894 ^ n18865;
  assign n18814 = n18813 ^ n16158;
  assign n18843 = n18842 ^ n18814;
  assign n18844 = n18783 ^ n16166;
  assign n18845 = n18810 ^ n18785;
  assign n18846 = n18844 & n18845;
  assign n18896 = n18843 & n18846;
  assign n19255 = n18895 & n18896;
  assign n19256 = n19254 & n19255;
  assign n19257 = n19150 ^ n19142;
  assign n19258 = ~n19256 & n19257;
  assign n19259 = n19155 ^ n16148;
  assign n19260 = n19259 ^ n19153;
  assign n19261 = ~n19258 & ~n19260;
  assign n19262 = n19160 ^ n16144;
  assign n19263 = ~n19261 & ~n19262;
  assign n19342 = n19264 ^ n19263;
  assign n19343 = n19342 ^ n1963;
  assign n19366 = n19262 ^ n19261;
  assign n19344 = n19260 ^ n19258;
  assign n19345 = n19344 ^ n1942;
  assign n19346 = n19257 ^ n19256;
  assign n19347 = n19346 ^ n1643;
  assign n19348 = n19255 ^ n19254;
  assign n19352 = n19351 ^ n19348;
  assign n18897 = n18896 ^ n18895;
  assign n19353 = n18897 ^ n1455;
  assign n18847 = n18846 ^ n18843;
  assign n18848 = n18847 ^ n1478;
  assign n18852 = ~n18844 & n18851;
  assign n18853 = n18852 ^ n1505;
  assign n18854 = n18845 ^ n18844;
  assign n18855 = n18854 ^ n18852;
  assign n18856 = n18853 & ~n18855;
  assign n18857 = n18856 ^ n1505;
  assign n18858 = n18857 ^ n18847;
  assign n18859 = n18848 & ~n18858;
  assign n18860 = n18859 ^ n1478;
  assign n19354 = n18897 ^ n18860;
  assign n19355 = n19353 & ~n19354;
  assign n19356 = n19355 ^ n1455;
  assign n19357 = n19356 ^ n19348;
  assign n19358 = n19352 & ~n19357;
  assign n19359 = n19358 ^ n19351;
  assign n19360 = n19359 ^ n19346;
  assign n19361 = n19347 & ~n19360;
  assign n19362 = n19361 ^ n1643;
  assign n19363 = n19362 ^ n19344;
  assign n19364 = n19345 & ~n19363;
  assign n19365 = n19364 ^ n1942;
  assign n19367 = n19366 ^ n19365;
  assign n19368 = n19366 ^ n1948;
  assign n19369 = n19367 & ~n19368;
  assign n19370 = n19369 ^ n1948;
  assign n19371 = n19370 ^ n19342;
  assign n19372 = ~n19343 & n19371;
  assign n19373 = n19372 ^ n1963;
  assign n19779 = n19373 ^ n2094;
  assign n19166 = n19165 ^ n19163;
  assign n19167 = ~n19164 & ~n19166;
  assign n19168 = n19167 ^ n16140;
  assign n19012 = n19011 ^ n18957;
  assign n19013 = n18960 & ~n19012;
  assign n19014 = n19013 ^ n18959;
  assign n18953 = n18430 ^ n17822;
  assign n18954 = n18953 ^ n16992;
  assign n19138 = n19014 ^ n18954;
  assign n18955 = n18378 ^ n1719;
  assign n19139 = n19138 ^ n18955;
  assign n19140 = n19139 ^ n16135;
  assign n19266 = n19168 ^ n19140;
  assign n19265 = n19263 & n19264;
  assign n19374 = n19266 ^ n19265;
  assign n19780 = n19779 ^ n19374;
  assign n18410 = n18409 ^ n1982;
  assign n20891 = n19780 ^ n18410;
  assign n19018 = n18381 ^ n1728;
  assign n19019 = n19018 ^ n18350;
  assign n19531 = n19019 ^ n17862;
  assign n19532 = n19531 ^ n18435;
  assign n19499 = n18955 ^ n18439;
  assign n19500 = n19499 ^ n17807;
  assign n19100 = n18753 ^ n18670;
  assign n19093 = n18750 ^ n18672;
  assign n19086 = n18747 ^ n18674;
  assign n18910 = n18744 ^ n772;
  assign n18911 = n18910 ^ n18675;
  assign n18908 = n18883 ^ n16913;
  assign n18909 = n18908 ^ n17618;
  assign n18912 = n18911 ^ n18909;
  assign n18915 = n18741 ^ n763;
  assign n18916 = n18915 ^ n18677;
  assign n18913 = n18834 ^ n18249;
  assign n18914 = n18913 ^ n17599;
  assign n18917 = n18916 ^ n18914;
  assign n18920 = n18775 ^ n18185;
  assign n18921 = n18920 ^ n17341;
  assign n18919 = n18735 ^ n689;
  assign n18922 = n18921 ^ n18919;
  assign n18924 = n18658 ^ n18165;
  assign n18925 = n18924 ^ n17184;
  assign n18923 = n18730 ^ n18685;
  assign n18926 = n18925 ^ n18923;
  assign n19061 = n18727 ^ n18690;
  assign n18928 = n18629 ^ n18009;
  assign n18929 = n18928 ^ n16947;
  assign n18927 = n18724 ^ n18695;
  assign n18930 = n18929 ^ n18927;
  assign n19051 = n18721 ^ n18700;
  assign n18933 = n18601 ^ n16958;
  assign n18934 = n18933 ^ n17919;
  assign n18931 = n18718 ^ n590;
  assign n18932 = n18931 ^ n18701;
  assign n18935 = n18934 ^ n18932;
  assign n18937 = n18586 ^ n17828;
  assign n18938 = n18937 ^ n16962;
  assign n18936 = n18715 ^ n18707;
  assign n18939 = n18938 ^ n18936;
  assign n18941 = n18549 ^ n16967;
  assign n18942 = n18941 ^ n17832;
  assign n18940 = n18712 ^ n2181;
  assign n18943 = n18942 ^ n18940;
  assign n18944 = n17836 ^ n16969;
  assign n18945 = n18944 ^ n18533;
  assign n18946 = n18945 ^ n18410;
  assign n18947 = n18421 ^ n17841;
  assign n18948 = n18947 ^ n16975;
  assign n18412 = n18390 ^ n1993;
  assign n18413 = n18412 ^ n18344;
  assign n18949 = n18948 ^ n18413;
  assign n19029 = n18387 ^ n18347;
  assign n18950 = n17820 ^ n16982;
  assign n18951 = n18950 ^ n17850;
  assign n18900 = n18384 ^ n18349;
  assign n18952 = n18951 ^ n18900;
  assign n18956 = n18955 ^ n18954;
  assign n19015 = n19014 ^ n18955;
  assign n19016 = n18956 & ~n19015;
  assign n19017 = n19016 ^ n18954;
  assign n19020 = n19019 ^ n19017;
  assign n19021 = n17891 ^ n16986;
  assign n19022 = n19021 ^ n18414;
  assign n19023 = n19022 ^ n19019;
  assign n19024 = ~n19020 & n19023;
  assign n19025 = n19024 ^ n19022;
  assign n19026 = n19025 ^ n18900;
  assign n19027 = ~n18952 & ~n19026;
  assign n19028 = n19027 ^ n18951;
  assign n19030 = n19029 ^ n19028;
  assign n19031 = n18422 ^ n17848;
  assign n19032 = n19031 ^ n16979;
  assign n19033 = n19032 ^ n19029;
  assign n19034 = ~n19030 & n19033;
  assign n19035 = n19034 ^ n19032;
  assign n19036 = n19035 ^ n18413;
  assign n19037 = ~n18949 & ~n19036;
  assign n19038 = n19037 ^ n18948;
  assign n19039 = n19038 ^ n18410;
  assign n19040 = n18946 & ~n19039;
  assign n19041 = n19040 ^ n18945;
  assign n19042 = n19041 ^ n18940;
  assign n19043 = n18943 & ~n19042;
  assign n19044 = n19043 ^ n18942;
  assign n19045 = n19044 ^ n18936;
  assign n19046 = ~n18939 & ~n19045;
  assign n19047 = n19046 ^ n18938;
  assign n19048 = n19047 ^ n18934;
  assign n19049 = n18935 & ~n19048;
  assign n19050 = n19049 ^ n19047;
  assign n19052 = n19051 ^ n19050;
  assign n19053 = n17996 ^ n16952;
  assign n19054 = n19053 ^ n18615;
  assign n19055 = n19054 ^ n19051;
  assign n19056 = ~n19052 & n19055;
  assign n19057 = n19056 ^ n19054;
  assign n19058 = n19057 ^ n18927;
  assign n19059 = ~n18930 & n19058;
  assign n19060 = n19059 ^ n18929;
  assign n19062 = n19061 ^ n19060;
  assign n19063 = n18147 ^ n16941;
  assign n19064 = n19063 ^ n18644;
  assign n19065 = n19064 ^ n19061;
  assign n19066 = ~n19062 & ~n19065;
  assign n19067 = n19066 ^ n19064;
  assign n19068 = n19067 ^ n18923;
  assign n19069 = n18926 & n19068;
  assign n19070 = n19069 ^ n18925;
  assign n19071 = n19070 ^ n18919;
  assign n19072 = ~n18922 & ~n19071;
  assign n19073 = n19072 ^ n18921;
  assign n18918 = n18738 ^ n18680;
  assign n19074 = n19073 ^ n18918;
  assign n19075 = n18800 ^ n17349;
  assign n19076 = n19075 ^ n18203;
  assign n19077 = n19076 ^ n18918;
  assign n19078 = n19074 & ~n19077;
  assign n19079 = n19078 ^ n19076;
  assign n19080 = n19079 ^ n18916;
  assign n19081 = ~n18917 & n19080;
  assign n19082 = n19081 ^ n18914;
  assign n19083 = n19082 ^ n18911;
  assign n19084 = ~n18912 & n19083;
  assign n19085 = n19084 ^ n18909;
  assign n19087 = n19086 ^ n19085;
  assign n19088 = n18984 ^ n17623;
  assign n19089 = n19088 ^ n16908;
  assign n19090 = n19089 ^ n19086;
  assign n19091 = n19087 & ~n19090;
  assign n19092 = n19091 ^ n19089;
  assign n19094 = n19093 ^ n19092;
  assign n19095 = n17612 ^ n17100;
  assign n19096 = n19095 ^ n18215;
  assign n19097 = n19096 ^ n19093;
  assign n19098 = ~n19094 & ~n19097;
  assign n19099 = n19098 ^ n19096;
  assign n19101 = n19100 ^ n19099;
  assign n18906 = n17609 ^ n17093;
  assign n18907 = n18906 ^ n18220;
  assign n19237 = n19100 ^ n18907;
  assign n19238 = ~n19101 & n19237;
  assign n19239 = n19238 ^ n18907;
  assign n19236 = n18756 ^ n18668;
  assign n19240 = n19239 ^ n19236;
  assign n19234 = n17605 ^ n17089;
  assign n19235 = n19234 ^ n18224;
  assign n19241 = n19240 ^ n19235;
  assign n19242 = n19241 ^ n16409;
  assign n19102 = n19101 ^ n18907;
  assign n19103 = n19102 ^ n16413;
  assign n19104 = n19096 ^ n19094;
  assign n19105 = n19104 ^ n16430;
  assign n19106 = n19089 ^ n19087;
  assign n19107 = n19106 ^ n16423;
  assign n19108 = n19082 ^ n18912;
  assign n19109 = n19108 ^ n16418;
  assign n19110 = n19079 ^ n18917;
  assign n19111 = n19110 ^ n16943;
  assign n19112 = n19076 ^ n19074;
  assign n19113 = n19112 ^ n16949;
  assign n19114 = n19070 ^ n18922;
  assign n19115 = n19114 ^ n16955;
  assign n19116 = n19067 ^ n18925;
  assign n19117 = n19116 ^ n18923;
  assign n19118 = n19117 ^ n16901;
  assign n19119 = n19064 ^ n19062;
  assign n19120 = n19119 ^ n16670;
  assign n19202 = n19057 ^ n18930;
  assign n19121 = n19054 ^ n19052;
  assign n19122 = n19121 ^ n16511;
  assign n19123 = n19047 ^ n18935;
  assign n19124 = n19123 ^ n16096;
  assign n19125 = n19044 ^ n18938;
  assign n19126 = n19125 ^ n18936;
  assign n19127 = n19126 ^ n16097;
  assign n19128 = n19041 ^ n18943;
  assign n19129 = n19128 ^ n16102;
  assign n19130 = n19038 ^ n18946;
  assign n19131 = n19130 ^ n16107;
  assign n19132 = n19035 ^ n18949;
  assign n19133 = n19132 ^ n16112;
  assign n19134 = n19032 ^ n19030;
  assign n19135 = n19134 ^ n16117;
  assign n19175 = n19025 ^ n18951;
  assign n19176 = n19175 ^ n18900;
  assign n19136 = n19022 ^ n19020;
  assign n19137 = n19136 ^ n16127;
  assign n19169 = n19168 ^ n19139;
  assign n19170 = n19140 & n19169;
  assign n19171 = n19170 ^ n16135;
  assign n19172 = n19171 ^ n19136;
  assign n19173 = n19137 & ~n19172;
  assign n19174 = n19173 ^ n16127;
  assign n19177 = n19176 ^ n19174;
  assign n19178 = n19176 ^ n16122;
  assign n19179 = n19177 & ~n19178;
  assign n19180 = n19179 ^ n16122;
  assign n19181 = n19180 ^ n19134;
  assign n19182 = n19135 & n19181;
  assign n19183 = n19182 ^ n16117;
  assign n19184 = n19183 ^ n19132;
  assign n19185 = ~n19133 & n19184;
  assign n19186 = n19185 ^ n16112;
  assign n19187 = n19186 ^ n19130;
  assign n19188 = ~n19131 & n19187;
  assign n19189 = n19188 ^ n16107;
  assign n19190 = n19189 ^ n19128;
  assign n19191 = n19129 & n19190;
  assign n19192 = n19191 ^ n16102;
  assign n19193 = n19192 ^ n19126;
  assign n19194 = n19127 & n19193;
  assign n19195 = n19194 ^ n16097;
  assign n19196 = n19195 ^ n19123;
  assign n19197 = ~n19124 & n19196;
  assign n19198 = n19197 ^ n16096;
  assign n19199 = n19198 ^ n19121;
  assign n19200 = ~n19122 & ~n19199;
  assign n19201 = n19200 ^ n16511;
  assign n19203 = n19202 ^ n19201;
  assign n19204 = n19202 ^ n16655;
  assign n19205 = ~n19203 & ~n19204;
  assign n19206 = n19205 ^ n16655;
  assign n19207 = n19206 ^ n19119;
  assign n19208 = n19120 & n19207;
  assign n19209 = n19208 ^ n16670;
  assign n19210 = n19209 ^ n19117;
  assign n19211 = n19118 & ~n19210;
  assign n19212 = n19211 ^ n16901;
  assign n19213 = n19212 ^ n19114;
  assign n19214 = ~n19115 & ~n19213;
  assign n19215 = n19214 ^ n16955;
  assign n19216 = n19215 ^ n19112;
  assign n19217 = ~n19113 & ~n19216;
  assign n19218 = n19217 ^ n16949;
  assign n19219 = n19218 ^ n19110;
  assign n19220 = ~n19111 & n19219;
  assign n19221 = n19220 ^ n16943;
  assign n19222 = n19221 ^ n19108;
  assign n19223 = ~n19109 & n19222;
  assign n19224 = n19223 ^ n16418;
  assign n19225 = n19224 ^ n19106;
  assign n19226 = ~n19107 & n19225;
  assign n19227 = n19226 ^ n16423;
  assign n19228 = n19227 ^ n19104;
  assign n19229 = ~n19105 & n19228;
  assign n19230 = n19229 ^ n16430;
  assign n19231 = n19230 ^ n19102;
  assign n19232 = ~n19103 & n19231;
  assign n19233 = n19232 ^ n16413;
  assign n19243 = n19242 ^ n19233;
  assign n19244 = n19227 ^ n19105;
  assign n19245 = n19224 ^ n19107;
  assign n19246 = n19212 ^ n19115;
  assign n19247 = n19209 ^ n19118;
  assign n19248 = n19195 ^ n19124;
  assign n19249 = n19192 ^ n19127;
  assign n19250 = n19183 ^ n19133;
  assign n19251 = n19180 ^ n16117;
  assign n19252 = n19251 ^ n19134;
  assign n19253 = n19171 ^ n19137;
  assign n19267 = n19265 & n19266;
  assign n19268 = n19253 & ~n19267;
  assign n19269 = n19177 ^ n16122;
  assign n19270 = ~n19268 & n19269;
  assign n19271 = n19252 & ~n19270;
  assign n19272 = ~n19250 & ~n19271;
  assign n19273 = n19186 ^ n19131;
  assign n19274 = n19272 & ~n19273;
  assign n19275 = n19189 ^ n19129;
  assign n19276 = n19274 & n19275;
  assign n19277 = ~n19249 & n19276;
  assign n19278 = n19248 & ~n19277;
  assign n19279 = n19198 ^ n16511;
  assign n19280 = n19279 ^ n19121;
  assign n19281 = n19278 & n19280;
  assign n19282 = n19203 ^ n16655;
  assign n19283 = ~n19281 & n19282;
  assign n19284 = n19206 ^ n16670;
  assign n19285 = n19284 ^ n19119;
  assign n19286 = n19283 & n19285;
  assign n19287 = n19247 & ~n19286;
  assign n19288 = n19246 & ~n19287;
  assign n19289 = n19215 ^ n19113;
  assign n19290 = n19288 & ~n19289;
  assign n19291 = n19218 ^ n19111;
  assign n19292 = ~n19290 & ~n19291;
  assign n19293 = n19221 ^ n19109;
  assign n19294 = ~n19292 & n19293;
  assign n19295 = n19245 & n19294;
  assign n19296 = n19244 & n19295;
  assign n19297 = n19230 ^ n19103;
  assign n19298 = ~n19296 & ~n19297;
  assign n19457 = ~n19243 & ~n19298;
  assign n19468 = n17031 ^ n16931;
  assign n19469 = n19468 ^ n18211;
  assign n19465 = n18759 ^ n1298;
  assign n19466 = n19465 ^ n18665;
  assign n19462 = n19236 ^ n19235;
  assign n19463 = n19240 & ~n19462;
  assign n19464 = n19463 ^ n19235;
  assign n19467 = n19466 ^ n19464;
  assign n19470 = n19469 ^ n19467;
  assign n19458 = n19241 ^ n19233;
  assign n19459 = n19242 & ~n19458;
  assign n19460 = n19459 ^ n16409;
  assign n19461 = n19460 ^ n16174;
  assign n19471 = n19470 ^ n19461;
  assign n19496 = n19457 & n19471;
  assign n19492 = n18762 ^ n2379;
  assign n19493 = n19492 ^ n18663;
  assign n19489 = n18256 ^ n16925;
  assign n19490 = n19489 ^ n17025;
  assign n19486 = n19469 ^ n19466;
  assign n19487 = ~n19467 & n19486;
  assign n19488 = n19487 ^ n19469;
  assign n19491 = n19490 ^ n19488;
  assign n19494 = n19493 ^ n19491;
  assign n19481 = n19470 ^ n16174;
  assign n19482 = n19470 ^ n19460;
  assign n19483 = ~n19481 & n19482;
  assign n19484 = n19483 ^ n16174;
  assign n19485 = n19484 ^ n16170;
  assign n19495 = n19494 ^ n19485;
  assign n19497 = n19496 ^ n19495;
  assign n19472 = n19471 ^ n19457;
  assign n19299 = n19298 ^ n19243;
  assign n19300 = n19299 ^ n2584;
  assign n19449 = n19297 ^ n19296;
  assign n19301 = n19295 ^ n19244;
  assign n2316 = n2276 ^ x421;
  assign n2317 = n2316 ^ n2309;
  assign n2318 = n2317 ^ x357;
  assign n19302 = n19301 ^ n2318;
  assign n19438 = n19294 ^ n19245;
  assign n19303 = n19293 ^ n19292;
  assign n1306 = n1209 ^ x423;
  assign n1310 = n1309 ^ n1306;
  assign n1311 = n1310 ^ x359;
  assign n19304 = n19303 ^ n1311;
  assign n19305 = n19291 ^ n19290;
  assign n19306 = n19305 ^ n1129;
  assign n19427 = n19289 ^ n19288;
  assign n19307 = n19287 ^ n19246;
  assign n19308 = n19307 ^ n968;
  assign n19419 = n19286 ^ n19247;
  assign n19309 = n19285 ^ n19283;
  assign n19310 = n19309 ^ n852;
  assign n19411 = n19282 ^ n19281;
  assign n19403 = n19280 ^ n19278;
  assign n19311 = n19277 ^ n19248;
  assign n19315 = n19314 ^ n19311;
  assign n19316 = n19276 ^ n19249;
  assign n19317 = n19316 ^ n530;
  assign n19319 = n17451 ^ x433;
  assign n19320 = n19319 ^ n575;
  assign n19321 = n19320 ^ x369;
  assign n19318 = n19275 ^ n19274;
  assign n19322 = n19321 ^ n19318;
  assign n19323 = n19273 ^ n19272;
  assign n19324 = n19323 ^ n612;
  assign n19325 = n19271 ^ n19250;
  assign n19329 = n19328 ^ n19325;
  assign n19330 = n19270 ^ n19252;
  assign n19334 = n19333 ^ n19330;
  assign n19335 = n19269 ^ n19268;
  assign n19339 = n19338 ^ n19335;
  assign n19340 = n19267 ^ n19253;
  assign n19341 = n19340 ^ n2107;
  assign n19375 = n19374 ^ n19373;
  assign n19376 = n19374 ^ n2094;
  assign n19377 = n19375 & ~n19376;
  assign n19378 = n19377 ^ n2094;
  assign n19379 = n19378 ^ n19340;
  assign n19380 = ~n19341 & n19379;
  assign n19381 = n19380 ^ n2107;
  assign n19382 = n19381 ^ n19335;
  assign n19383 = n19339 & ~n19382;
  assign n19384 = n19383 ^ n19338;
  assign n19385 = n19384 ^ n19330;
  assign n19386 = ~n19334 & n19385;
  assign n19387 = n19386 ^ n19333;
  assign n19388 = n19387 ^ n19325;
  assign n19389 = ~n19329 & n19388;
  assign n19390 = n19389 ^ n19328;
  assign n19391 = n19390 ^ n19323;
  assign n19392 = n19324 & ~n19391;
  assign n19393 = n19392 ^ n612;
  assign n19394 = n19393 ^ n19318;
  assign n19395 = ~n19322 & n19394;
  assign n19396 = n19395 ^ n19321;
  assign n19397 = n19396 ^ n19316;
  assign n19398 = n19317 & ~n19397;
  assign n19399 = n19398 ^ n530;
  assign n19400 = n19399 ^ n19311;
  assign n19401 = ~n19315 & n19400;
  assign n19402 = n19401 ^ n19314;
  assign n19404 = n19403 ^ n19402;
  assign n19408 = n19407 ^ n19403;
  assign n19409 = ~n19404 & n19408;
  assign n19410 = n19409 ^ n19407;
  assign n19412 = n19411 ^ n19410;
  assign n19413 = n19411 ^ n843;
  assign n19414 = ~n19412 & n19413;
  assign n19415 = n19414 ^ n843;
  assign n19416 = n19415 ^ n19309;
  assign n19417 = ~n19310 & n19416;
  assign n19418 = n19417 ^ n852;
  assign n19420 = n19419 ^ n19418;
  assign n19421 = n19419 ^ n867;
  assign n19422 = n19420 & ~n19421;
  assign n19423 = n19422 ^ n867;
  assign n19424 = n19423 ^ n19307;
  assign n19425 = n19308 & ~n19424;
  assign n19426 = n19425 ^ n968;
  assign n19428 = n19427 ^ n19426;
  assign n19429 = n19427 ^ n1120;
  assign n19430 = ~n19428 & n19429;
  assign n19431 = n19430 ^ n1120;
  assign n19432 = n19431 ^ n19305;
  assign n19433 = n19306 & ~n19432;
  assign n19434 = n19433 ^ n1129;
  assign n19435 = n19434 ^ n19303;
  assign n19436 = n19304 & ~n19435;
  assign n19437 = n19436 ^ n1311;
  assign n19439 = n19438 ^ n19437;
  assign n19440 = n17431 ^ x422;
  assign n19441 = n19440 ^ n1315;
  assign n19442 = n19441 ^ x358;
  assign n19443 = n19442 ^ n19438;
  assign n19444 = n19439 & ~n19443;
  assign n19445 = n19444 ^ n19442;
  assign n19446 = n19445 ^ n19301;
  assign n19447 = ~n19302 & n19446;
  assign n19448 = n19447 ^ n2318;
  assign n19450 = n19449 ^ n19448;
  assign n2593 = n2508 ^ x420;
  assign n2594 = n2593 ^ n1538;
  assign n2595 = n2594 ^ x356;
  assign n19451 = n19449 ^ n2595;
  assign n19452 = ~n19450 & n19451;
  assign n19453 = n19452 ^ n2595;
  assign n19454 = n19453 ^ n19299;
  assign n19455 = ~n19300 & n19454;
  assign n19456 = n19455 ^ n2584;
  assign n19473 = n19472 ^ n19456;
  assign n19474 = n19472 ^ n2608;
  assign n19475 = n19473 & ~n19474;
  assign n19476 = n19475 ^ n2608;
  assign n19480 = n19479 ^ n19476;
  assign n19498 = n19497 ^ n19480;
  assign n19501 = n19500 ^ n19498;
  assign n19520 = n19473 ^ n2608;
  assign n19503 = n18962 ^ n18403;
  assign n19504 = n19503 ^ n17722;
  assign n19502 = n19453 ^ n19300;
  assign n19505 = n19504 ^ n19502;
  assign n19508 = n19445 ^ n19302;
  assign n19509 = n18999 ^ n17644;
  assign n19510 = n19509 ^ n18322;
  assign n19511 = ~n19508 & n19510;
  assign n19506 = n18339 ^ n17690;
  assign n19507 = n19506 ^ n18968;
  assign n19512 = n19511 ^ n19507;
  assign n19513 = n19450 ^ n2595;
  assign n19514 = n19513 ^ n19507;
  assign n19515 = ~n19512 & n19514;
  assign n19516 = n19515 ^ n19511;
  assign n19517 = n19516 ^ n19502;
  assign n19518 = n19505 & n19517;
  assign n19519 = n19518 ^ n19504;
  assign n19521 = n19520 ^ n19519;
  assign n19522 = n18957 ^ n18444;
  assign n19523 = n19522 ^ n17736;
  assign n19524 = n19523 ^ n19519;
  assign n19525 = ~n19521 & n19524;
  assign n19526 = n19525 ^ n19523;
  assign n19527 = n19526 ^ n19498;
  assign n19528 = n19501 & n19527;
  assign n19529 = n19528 ^ n19500;
  assign n18905 = n18851 ^ n18844;
  assign n19530 = n19529 ^ n18905;
  assign n19560 = n19532 ^ n19530;
  assign n19561 = n19560 ^ n17135;
  assign n19562 = n19526 ^ n19501;
  assign n19563 = n19562 ^ n16927;
  assign n19564 = n19523 ^ n19521;
  assign n19565 = n19564 ^ n16932;
  assign n19566 = n19516 ^ n19505;
  assign n19567 = n19566 ^ n16937;
  assign n19568 = n19510 ^ n19508;
  assign n19569 = ~n17021 & ~n19568;
  assign n19570 = n19569 ^ n17017;
  assign n19571 = n19513 ^ n19512;
  assign n19572 = n19571 ^ n19569;
  assign n19573 = ~n19570 & n19572;
  assign n19574 = n19573 ^ n17017;
  assign n19575 = n19574 ^ n19566;
  assign n19576 = ~n19567 & n19575;
  assign n19577 = n19576 ^ n16937;
  assign n19578 = n19577 ^ n19564;
  assign n19579 = n19565 & ~n19578;
  assign n19580 = n19579 ^ n16932;
  assign n19581 = n19580 ^ n19562;
  assign n19582 = n19563 & ~n19581;
  assign n19583 = n19582 ^ n16927;
  assign n19584 = n19583 ^ n19560;
  assign n19585 = ~n19561 & n19584;
  assign n19586 = n19585 ^ n17135;
  assign n19533 = n19532 ^ n18905;
  assign n19534 = n19530 & n19533;
  assign n19535 = n19534 ^ n19532;
  assign n18903 = n18854 ^ n18853;
  assign n18901 = n18900 ^ n18431;
  assign n18902 = n18901 ^ n17872;
  assign n18904 = n18903 ^ n18902;
  assign n19558 = n19535 ^ n18904;
  assign n19559 = n19558 ^ n17002;
  assign n19620 = n19586 ^ n19559;
  assign n19609 = n19580 ^ n19563;
  assign n19610 = n19577 ^ n19565;
  assign n19611 = n19574 ^ n19567;
  assign n19612 = n19568 ^ n17021;
  assign n19613 = n19571 ^ n19570;
  assign n19614 = n19612 & n19613;
  assign n19615 = n19611 & n19614;
  assign n19616 = ~n19610 & n19615;
  assign n19617 = ~n19609 & n19616;
  assign n19618 = n19583 ^ n19561;
  assign n19619 = ~n19617 & ~n19618;
  assign n19667 = n19620 ^ n19619;
  assign n19668 = n19667 ^ n1708;
  assign n19699 = n19618 ^ n19617;
  assign n19669 = n19616 ^ n19609;
  assign n19670 = n19669 ^ n1618;
  assign n19671 = n19615 ^ n19610;
  assign n19672 = n19671 ^ n1609;
  assign n19676 = n19614 ^ n19611;
  assign n19677 = n19676 ^ n19675;
  assign n19681 = ~n19612 & n19680;
  assign n19685 = n19684 ^ n19681;
  assign n19686 = n19613 ^ n19612;
  assign n19687 = n19686 ^ n19681;
  assign n19688 = n19685 & ~n19687;
  assign n19689 = n19688 ^ n19684;
  assign n19690 = n19689 ^ n19676;
  assign n19691 = n19677 & ~n19690;
  assign n19692 = n19691 ^ n19675;
  assign n19693 = n19692 ^ n19671;
  assign n19694 = ~n19672 & n19693;
  assign n19695 = n19694 ^ n1609;
  assign n19696 = n19695 ^ n19669;
  assign n19697 = ~n19670 & n19696;
  assign n19698 = n19697 ^ n1618;
  assign n19700 = n19699 ^ n19698;
  assign n19701 = n19699 ^ n1699;
  assign n19702 = n19700 & ~n19701;
  assign n19703 = n19702 ^ n1699;
  assign n19704 = n19703 ^ n19667;
  assign n19705 = n19668 & ~n19704;
  assign n19706 = n19705 ^ n1708;
  assign n19587 = n19586 ^ n19558;
  assign n19588 = n19559 & ~n19587;
  assign n19589 = n19588 ^ n17002;
  assign n19542 = n19029 ^ n18430;
  assign n19543 = n19542 ^ n17860;
  assign n19539 = n18857 ^ n1478;
  assign n19540 = n19539 ^ n18847;
  assign n19536 = n19535 ^ n18903;
  assign n19537 = n18904 & n19536;
  assign n19538 = n19537 ^ n18902;
  assign n19541 = n19540 ^ n19538;
  assign n19556 = n19543 ^ n19541;
  assign n19557 = n19556 ^ n16998;
  assign n19622 = n19589 ^ n19557;
  assign n19621 = ~n19619 & ~n19620;
  assign n19665 = n19622 ^ n19621;
  assign n19666 = n19665 ^ n1820;
  assign n20370 = n19706 ^ n19666;
  assign n20892 = n20891 ^ n20370;
  assign n20122 = n18962 ^ n18905;
  assign n20123 = n20122 ^ n18322;
  assign n20028 = n19423 ^ n19308;
  assign n20008 = n19420 ^ n867;
  assign n19923 = n19415 ^ n19310;
  assign n19761 = n19093 ^ n18834;
  assign n19762 = n19761 ^ n18185;
  assign n19760 = n19399 ^ n19315;
  assign n19763 = n19762 ^ n19760;
  assign n19765 = n19086 ^ n18165;
  assign n19766 = n19765 ^ n18800;
  assign n19764 = n19396 ^ n19317;
  assign n19767 = n19766 ^ n19764;
  assign n19771 = n18916 ^ n18658;
  assign n19772 = n19771 ^ n18009;
  assign n19769 = n19390 ^ n612;
  assign n19770 = n19769 ^ n19323;
  assign n19773 = n19772 ^ n19770;
  assign n19775 = n18919 ^ n17919;
  assign n19776 = n19775 ^ n18629;
  assign n19774 = n19384 ^ n19334;
  assign n19777 = n19776 ^ n19774;
  assign n19796 = n19381 ^ n19339;
  assign n19737 = n19370 ^ n1963;
  assign n19738 = n19737 ^ n19342;
  assign n19651 = n19367 ^ n1948;
  assign n19637 = n19362 ^ n19345;
  assign n19604 = n19359 ^ n19347;
  assign n19550 = n19356 ^ n19352;
  assign n18861 = n18860 ^ n1455;
  assign n18898 = n18897 ^ n18861;
  assign n18415 = n18414 ^ n18413;
  assign n18416 = n18415 ^ n17854;
  assign n18899 = n18898 ^ n18416;
  assign n19544 = n19543 ^ n19540;
  assign n19545 = ~n19541 & n19544;
  assign n19546 = n19545 ^ n19543;
  assign n19547 = n19546 ^ n18898;
  assign n19548 = ~n18899 & ~n19547;
  assign n19549 = n19548 ^ n18416;
  assign n19551 = n19550 ^ n19549;
  assign n17823 = n17822 ^ n17820;
  assign n18411 = n18410 ^ n17823;
  assign n19601 = n19550 ^ n18411;
  assign n19602 = n19551 & n19601;
  assign n19603 = n19602 ^ n18411;
  assign n19605 = n19604 ^ n19603;
  assign n19599 = n18422 ^ n17891;
  assign n19600 = n19599 ^ n18940;
  assign n19634 = n19604 ^ n19600;
  assign n19635 = ~n19605 & n19634;
  assign n19636 = n19635 ^ n19600;
  assign n19638 = n19637 ^ n19636;
  assign n19632 = n18421 ^ n17850;
  assign n19633 = n19632 ^ n18936;
  assign n19648 = n19637 ^ n19633;
  assign n19649 = ~n19638 & ~n19648;
  assign n19650 = n19649 ^ n19633;
  assign n19652 = n19651 ^ n19650;
  assign n19646 = n18932 ^ n17848;
  assign n19647 = n19646 ^ n18533;
  assign n19734 = n19651 ^ n19647;
  assign n19735 = ~n19652 & n19734;
  assign n19736 = n19735 ^ n19647;
  assign n19739 = n19738 ^ n19736;
  assign n19732 = n19051 ^ n18549;
  assign n19733 = n19732 ^ n17841;
  assign n19781 = n19738 ^ n19733;
  assign n19782 = ~n19739 & n19781;
  assign n19783 = n19782 ^ n19733;
  assign n19784 = n19783 ^ n19780;
  assign n19785 = n18586 ^ n17836;
  assign n19786 = n19785 ^ n18927;
  assign n19787 = n19786 ^ n19780;
  assign n19788 = ~n19784 & n19787;
  assign n19789 = n19788 ^ n19786;
  assign n19778 = n19378 ^ n19341;
  assign n19790 = n19789 ^ n19778;
  assign n19791 = n19061 ^ n17832;
  assign n19792 = n19791 ^ n18601;
  assign n19793 = n19792 ^ n19778;
  assign n19794 = ~n19790 & n19793;
  assign n19795 = n19794 ^ n19792;
  assign n19797 = n19796 ^ n19795;
  assign n19798 = n18923 ^ n17828;
  assign n19799 = n19798 ^ n18615;
  assign n19800 = n19799 ^ n19796;
  assign n19801 = n19797 & n19800;
  assign n19802 = n19801 ^ n19799;
  assign n19803 = n19802 ^ n19774;
  assign n19804 = n19777 & n19803;
  assign n19805 = n19804 ^ n19776;
  assign n19750 = n19387 ^ n19328;
  assign n19751 = n19750 ^ n19325;
  assign n19806 = n19805 ^ n19751;
  assign n19807 = n18918 ^ n17996;
  assign n19808 = n19807 ^ n18644;
  assign n19809 = n19808 ^ n19751;
  assign n19810 = ~n19806 & n19809;
  assign n19811 = n19810 ^ n19808;
  assign n19812 = n19811 ^ n19770;
  assign n19813 = n19773 & n19812;
  assign n19814 = n19813 ^ n19772;
  assign n19768 = n19393 ^ n19322;
  assign n19815 = n19814 ^ n19768;
  assign n19816 = n18775 ^ n18147;
  assign n19817 = n19816 ^ n18911;
  assign n19818 = n19817 ^ n19768;
  assign n19819 = n19815 & ~n19818;
  assign n19820 = n19819 ^ n19817;
  assign n19821 = n19820 ^ n19764;
  assign n19822 = n19767 & ~n19821;
  assign n19823 = n19822 ^ n19766;
  assign n19824 = n19823 ^ n19760;
  assign n19825 = n19763 & n19824;
  assign n19826 = n19825 ^ n19762;
  assign n19759 = n19407 ^ n19404;
  assign n19827 = n19826 ^ n19759;
  assign n19757 = n19100 ^ n18203;
  assign n19758 = n19757 ^ n18883;
  assign n19884 = n19759 ^ n19758;
  assign n19885 = n19827 & ~n19884;
  assign n19886 = n19885 ^ n19758;
  assign n19883 = n19412 ^ n843;
  assign n19887 = n19886 ^ n19883;
  assign n19881 = n18984 ^ n18249;
  assign n19882 = n19881 ^ n19236;
  assign n19920 = n19883 ^ n19882;
  assign n19921 = n19887 & n19920;
  assign n19922 = n19921 ^ n19882;
  assign n19924 = n19923 ^ n19922;
  assign n19918 = n19466 ^ n17618;
  assign n19919 = n19918 ^ n18215;
  assign n20005 = n19923 ^ n19919;
  assign n20006 = n19924 & n20005;
  assign n20007 = n20006 ^ n19919;
  assign n20009 = n20008 ^ n20007;
  assign n20003 = n19493 ^ n18220;
  assign n20004 = n20003 ^ n17623;
  assign n20025 = n20008 ^ n20004;
  assign n20026 = ~n20009 & ~n20025;
  assign n20027 = n20026 ^ n20004;
  assign n20029 = n20028 ^ n20027;
  assign n20023 = n18782 ^ n17612;
  assign n20024 = n20023 ^ n18224;
  assign n20030 = n20029 ^ n20024;
  assign n20031 = n20030 ^ n17100;
  assign n20010 = n20009 ^ n20004;
  assign n20011 = n20010 ^ n16908;
  assign n19925 = n19924 ^ n19919;
  assign n19926 = n19925 ^ n16913;
  assign n19888 = n19887 ^ n19882;
  assign n19889 = n19888 ^ n17599;
  assign n19828 = n19827 ^ n19758;
  assign n19829 = n19828 ^ n17349;
  assign n19830 = n19823 ^ n19763;
  assign n19831 = n19830 ^ n17341;
  assign n19832 = n19820 ^ n19767;
  assign n19833 = n19832 ^ n17184;
  assign n19834 = n19817 ^ n19815;
  assign n19835 = n19834 ^ n16941;
  assign n19836 = n19811 ^ n19773;
  assign n19837 = n19836 ^ n16947;
  assign n19838 = n19808 ^ n19806;
  assign n19839 = n19838 ^ n16952;
  assign n19840 = n19802 ^ n19777;
  assign n19841 = n19840 ^ n16958;
  assign n19842 = n19799 ^ n19797;
  assign n19843 = n19842 ^ n16962;
  assign n19844 = n19792 ^ n19790;
  assign n19845 = n19844 ^ n16967;
  assign n19846 = n19786 ^ n19784;
  assign n19847 = n19846 ^ n16969;
  assign n19740 = n19739 ^ n19733;
  assign n19741 = n19740 ^ n16975;
  assign n19653 = n19652 ^ n19647;
  assign n19654 = n19653 ^ n16979;
  assign n19639 = n19638 ^ n19633;
  assign n19640 = n19639 ^ n16982;
  assign n19606 = n19605 ^ n19600;
  assign n19607 = n19606 ^ n16986;
  assign n19552 = n19551 ^ n18411;
  assign n19553 = n19552 ^ n16992;
  assign n19554 = n19546 ^ n18899;
  assign n19555 = n19554 ^ n16994;
  assign n19590 = n19589 ^ n19556;
  assign n19591 = ~n19557 & n19590;
  assign n19592 = n19591 ^ n16998;
  assign n19593 = n19592 ^ n19554;
  assign n19594 = ~n19555 & ~n19593;
  assign n19595 = n19594 ^ n16994;
  assign n19596 = n19595 ^ n19552;
  assign n19597 = ~n19553 & n19596;
  assign n19598 = n19597 ^ n16992;
  assign n19629 = n19606 ^ n19598;
  assign n19630 = n19607 & ~n19629;
  assign n19631 = n19630 ^ n16986;
  assign n19643 = n19639 ^ n19631;
  assign n19644 = ~n19640 & n19643;
  assign n19645 = n19644 ^ n16982;
  assign n19729 = n19653 ^ n19645;
  assign n19730 = n19654 & n19729;
  assign n19731 = n19730 ^ n16979;
  assign n19848 = n19740 ^ n19731;
  assign n19849 = n19741 & ~n19848;
  assign n19850 = n19849 ^ n16975;
  assign n19851 = n19850 ^ n19846;
  assign n19852 = ~n19847 & ~n19851;
  assign n19853 = n19852 ^ n16969;
  assign n19854 = n19853 ^ n19844;
  assign n19855 = n19845 & n19854;
  assign n19856 = n19855 ^ n16967;
  assign n19857 = n19856 ^ n19842;
  assign n19858 = ~n19843 & ~n19857;
  assign n19859 = n19858 ^ n16962;
  assign n19860 = n19859 ^ n19840;
  assign n19861 = ~n19841 & ~n19860;
  assign n19862 = n19861 ^ n16958;
  assign n19863 = n19862 ^ n19838;
  assign n19864 = n19839 & ~n19863;
  assign n19865 = n19864 ^ n16952;
  assign n19866 = n19865 ^ n19836;
  assign n19867 = n19837 & ~n19866;
  assign n19868 = n19867 ^ n16947;
  assign n19869 = n19868 ^ n19834;
  assign n19870 = n19835 & ~n19869;
  assign n19871 = n19870 ^ n16941;
  assign n19872 = n19871 ^ n19832;
  assign n19873 = n19833 & n19872;
  assign n19874 = n19873 ^ n17184;
  assign n19875 = n19874 ^ n19830;
  assign n19876 = ~n19831 & ~n19875;
  assign n19877 = n19876 ^ n17341;
  assign n19878 = n19877 ^ n19828;
  assign n19879 = ~n19829 & n19878;
  assign n19880 = n19879 ^ n17349;
  assign n19915 = n19888 ^ n19880;
  assign n19916 = ~n19889 & ~n19915;
  assign n19917 = n19916 ^ n17599;
  assign n20000 = n19925 ^ n19917;
  assign n20001 = n19926 & ~n20000;
  assign n20002 = n20001 ^ n16913;
  assign n20020 = n20010 ^ n20002;
  assign n20021 = ~n20011 & ~n20020;
  assign n20022 = n20021 ^ n16908;
  assign n20032 = n20031 ^ n20022;
  assign n20012 = n20011 ^ n20002;
  assign n19890 = n19889 ^ n19880;
  assign n19891 = n19865 ^ n19837;
  assign n19892 = n19862 ^ n19839;
  assign n19893 = n19856 ^ n19843;
  assign n19894 = n19853 ^ n16967;
  assign n19895 = n19894 ^ n19844;
  assign n19742 = n19741 ^ n19731;
  assign n19608 = n19607 ^ n19598;
  assign n19623 = ~n19621 & ~n19622;
  assign n19624 = n19592 ^ n19555;
  assign n19625 = n19623 & ~n19624;
  assign n19626 = n19595 ^ n19553;
  assign n19627 = n19625 & n19626;
  assign n19628 = n19608 & ~n19627;
  assign n19641 = n19640 ^ n19631;
  assign n19642 = ~n19628 & n19641;
  assign n19655 = n19654 ^ n19645;
  assign n19743 = ~n19642 & n19655;
  assign n19896 = n19742 & ~n19743;
  assign n19897 = n19850 ^ n16969;
  assign n19898 = n19897 ^ n19846;
  assign n19899 = n19896 & ~n19898;
  assign n19900 = ~n19895 & n19899;
  assign n19901 = ~n19893 & n19900;
  assign n19902 = n19859 ^ n19841;
  assign n19903 = ~n19901 & ~n19902;
  assign n19904 = ~n19892 & n19903;
  assign n19905 = n19891 & ~n19904;
  assign n19906 = n19868 ^ n19835;
  assign n19907 = n19905 & n19906;
  assign n19908 = n19871 ^ n19833;
  assign n19909 = ~n19907 & ~n19908;
  assign n19910 = n19874 ^ n19831;
  assign n19911 = ~n19909 & n19910;
  assign n19912 = n19877 ^ n19829;
  assign n19913 = n19911 & ~n19912;
  assign n19914 = n19890 & ~n19913;
  assign n19927 = n19926 ^ n19917;
  assign n20013 = ~n19914 & ~n19927;
  assign n20019 = n20012 & n20013;
  assign n20033 = n20032 ^ n20019;
  assign n20014 = n20013 ^ n20012;
  assign n19928 = n19927 ^ n19914;
  assign n1249 = n1152 ^ x455;
  assign n1250 = n1249 ^ n1243;
  assign n1251 = n1250 ^ x391;
  assign n19929 = n19928 ^ n1251;
  assign n19930 = n19913 ^ n19890;
  assign n1234 = n1137 ^ x456;
  assign n1235 = n1234 ^ n1105;
  assign n1236 = n1235 ^ x392;
  assign n19931 = n19930 ^ n1236;
  assign n19989 = n19912 ^ n19911;
  assign n19932 = n19910 ^ n19909;
  assign n19933 = n19932 ^ n1071;
  assign n19981 = n19908 ^ n19907;
  assign n19934 = n19906 ^ n19905;
  assign n19935 = n19934 ^ n758;
  assign n19970 = n19904 ^ n19891;
  assign n19936 = n19903 ^ n19892;
  assign n19937 = n19936 ^ n564;
  assign n19938 = n19902 ^ n19901;
  assign n659 = n643 ^ x463;
  assign n660 = n659 ^ n656;
  assign n661 = n660 ^ x399;
  assign n19939 = n19938 ^ n661;
  assign n19940 = n19900 ^ n19893;
  assign n647 = n634 ^ x464;
  assign n651 = n650 ^ n647;
  assign n652 = n651 ^ x400;
  assign n19941 = n19940 ^ n652;
  assign n19942 = n19899 ^ n19895;
  assign n19946 = n19945 ^ n19942;
  assign n19950 = n19898 ^ n19896;
  assign n19744 = n19743 ^ n19742;
  assign n19748 = n19747 ^ n19744;
  assign n19656 = n19655 ^ n19642;
  assign n19660 = n19659 ^ n19656;
  assign n19661 = n19641 ^ n19628;
  assign n19662 = n19661 ^ n2261;
  assign n19718 = n19627 ^ n19608;
  assign n19663 = n19626 ^ n19625;
  assign n19664 = n19663 ^ n1988;
  assign n19710 = n19624 ^ n19623;
  assign n19707 = n19706 ^ n19665;
  assign n19708 = ~n19666 & n19707;
  assign n19709 = n19708 ^ n1820;
  assign n19711 = n19710 ^ n19709;
  assign n19712 = n19710 ^ n2223;
  assign n19713 = ~n19711 & n19712;
  assign n19714 = n19713 ^ n2223;
  assign n19715 = n19714 ^ n19663;
  assign n19716 = ~n19664 & n19715;
  assign n19717 = n19716 ^ n1988;
  assign n19719 = n19718 ^ n19717;
  assign n19720 = n19718 ^ n2243;
  assign n19721 = n19719 & ~n19720;
  assign n19722 = n19721 ^ n2243;
  assign n19723 = n19722 ^ n19661;
  assign n19724 = n19662 & ~n19723;
  assign n19725 = n19724 ^ n2261;
  assign n19726 = n19725 ^ n19656;
  assign n19727 = ~n19660 & n19726;
  assign n19728 = n19727 ^ n19659;
  assign n19947 = n19744 ^ n19728;
  assign n19948 = n19748 & ~n19947;
  assign n19949 = n19948 ^ n19747;
  assign n19951 = n19950 ^ n19949;
  assign n19955 = n19954 ^ n19950;
  assign n19956 = ~n19951 & n19955;
  assign n19957 = n19956 ^ n19954;
  assign n19958 = n19957 ^ n19942;
  assign n19959 = n19946 & ~n19958;
  assign n19960 = n19959 ^ n19945;
  assign n19961 = n19960 ^ n19940;
  assign n19962 = n19941 & ~n19961;
  assign n19963 = n19962 ^ n652;
  assign n19964 = n19963 ^ n19938;
  assign n19965 = n19939 & ~n19964;
  assign n19966 = n19965 ^ n661;
  assign n19967 = n19966 ^ n19936;
  assign n19968 = ~n19937 & n19967;
  assign n19969 = n19968 ^ n564;
  assign n19971 = n19970 ^ n19969;
  assign n19975 = n19974 ^ n19970;
  assign n19976 = ~n19971 & n19975;
  assign n19977 = n19976 ^ n19974;
  assign n19978 = n19977 ^ n19934;
  assign n19979 = ~n19935 & n19978;
  assign n19980 = n19979 ^ n758;
  assign n19982 = n19981 ^ n19980;
  assign n19983 = n19981 ^ n1085;
  assign n19984 = ~n19982 & n19983;
  assign n19985 = n19984 ^ n1085;
  assign n19986 = n19985 ^ n19932;
  assign n19987 = n19933 & ~n19986;
  assign n19988 = n19987 ^ n1071;
  assign n19990 = n19989 ^ n19988;
  assign n19991 = n19989 ^ n1096;
  assign n19992 = ~n19990 & n19991;
  assign n19993 = n19992 ^ n1096;
  assign n19994 = n19993 ^ n19930;
  assign n19995 = ~n19931 & n19994;
  assign n19996 = n19995 ^ n1236;
  assign n19997 = n19996 ^ n19928;
  assign n19998 = ~n19929 & n19997;
  assign n19999 = n19998 ^ n1251;
  assign n20015 = n20014 ^ n19999;
  assign n20016 = n20014 ^ n2289;
  assign n20017 = n20015 & ~n20016;
  assign n20018 = n20017 ^ n2289;
  assign n20034 = n20033 ^ n20018;
  assign n2346 = n2306 ^ x453;
  assign n2347 = n2346 ^ n2294;
  assign n2348 = n2347 ^ x389;
  assign n20121 = n20034 ^ n2348;
  assign n20182 = n20123 ^ n20121;
  assign n20225 = n20182 ^ n17644;
  assign n20250 = n1523 & n20225;
  assign n20254 = n20253 ^ n20250;
  assign n20047 = n19428 ^ n1120;
  assign n20044 = n20028 ^ n20024;
  assign n20045 = ~n20029 & n20044;
  assign n20046 = n20045 ^ n20024;
  assign n20048 = n20047 ^ n20046;
  assign n20042 = n18808 ^ n18211;
  assign n20043 = n20042 ^ n17609;
  assign n20049 = n20048 ^ n20043;
  assign n20050 = n20049 ^ n17093;
  assign n20039 = n20030 ^ n20022;
  assign n20040 = n20031 & n20039;
  assign n20041 = n20040 ^ n17100;
  assign n20051 = n20050 ^ n20041;
  assign n20038 = n20019 & n20032;
  assign n20052 = n20051 ^ n20038;
  assign n20035 = n20033 ^ n2348;
  assign n20036 = n20034 & ~n20035;
  assign n20037 = n20036 ^ n2348;
  assign n20053 = n20052 ^ n20037;
  assign n20126 = n20053 ^ n2368;
  assign n20124 = ~n20121 & n20123;
  assign n20119 = n18903 ^ n18339;
  assign n20120 = n20119 ^ n18957;
  assign n20125 = n20124 ^ n20120;
  assign n20185 = n20126 ^ n20125;
  assign n20183 = n17644 & ~n20182;
  assign n20184 = n20183 ^ n17690;
  assign n20226 = n20185 ^ n20184;
  assign n20255 = n20226 ^ n20225;
  assign n20256 = n20255 ^ n20250;
  assign n20257 = n20254 & ~n20256;
  assign n20258 = n20257 ^ n20253;
  assign n20186 = n20185 ^ n20183;
  assign n20187 = ~n20184 & ~n20186;
  assign n20188 = n20187 ^ n17690;
  assign n20132 = n18955 ^ n18403;
  assign n20133 = n20132 ^ n19540;
  assign n20066 = n19431 ^ n19306;
  assign n20063 = n20047 ^ n20043;
  assign n20064 = ~n20048 & n20063;
  assign n20065 = n20064 ^ n20043;
  assign n20067 = n20066 ^ n20065;
  assign n20061 = n18840 ^ n17605;
  assign n20062 = n20061 ^ n18256;
  assign n20068 = n20067 ^ n20062;
  assign n20069 = n20068 ^ n17089;
  assign n20058 = n20049 ^ n20041;
  assign n20059 = n20050 & ~n20058;
  assign n20060 = n20059 ^ n17093;
  assign n20070 = n20069 ^ n20060;
  assign n20057 = ~n20038 & n20051;
  assign n20071 = n20070 ^ n20057;
  assign n20054 = n20052 ^ n2368;
  assign n20055 = n20053 & ~n20054;
  assign n20056 = n20055 ^ n2368;
  assign n20072 = n20071 ^ n20056;
  assign n2481 = n2420 ^ x451;
  assign n2485 = n2484 ^ n2481;
  assign n2486 = n2485 ^ x387;
  assign n20130 = n20072 ^ n2486;
  assign n20127 = n20126 ^ n20120;
  assign n20128 = ~n20125 & ~n20127;
  assign n20129 = n20128 ^ n20124;
  assign n20131 = n20130 ^ n20129;
  assign n20180 = n20133 ^ n20131;
  assign n20181 = n20180 ^ n17722;
  assign n20228 = n20188 ^ n20181;
  assign n20227 = ~n20225 & ~n20226;
  assign n20248 = n20228 ^ n20227;
  assign n20249 = n20248 ^ n1436;
  assign n20889 = n20258 ^ n20249;
  assign n20840 = n19738 ^ n18413;
  assign n20320 = n19703 ^ n19668;
  assign n20841 = n20840 ^ n20320;
  assign n20839 = n20255 ^ n20254;
  assign n20842 = n20841 ^ n20839;
  assign n20819 = n19651 ^ n19029;
  assign n20300 = n19700 ^ n1699;
  assign n20820 = n20819 ^ n20300;
  assign n20818 = n20225 ^ n1523;
  assign n20821 = n20820 ^ n20818;
  assign n20700 = n18999 ^ n18286;
  assign n20701 = n20700 ^ n19520;
  assign n20698 = n19996 ^ n19929;
  assign n20448 = n19990 ^ n1096;
  assign n20338 = n19977 ^ n19935;
  assign n20336 = n18782 ^ n18215;
  assign n20084 = n19434 ^ n19304;
  assign n20337 = n20336 ^ n20084;
  assign n20339 = n20338 ^ n20337;
  assign n20341 = n19493 ^ n18984;
  assign n20342 = n20341 ^ n20066;
  assign n20340 = n19974 ^ n19971;
  assign n20343 = n20342 ^ n20340;
  assign n20423 = n19966 ^ n19937;
  assign n20345 = n19236 ^ n18834;
  assign n20346 = n20345 ^ n20028;
  assign n20344 = n19963 ^ n19939;
  assign n20347 = n20346 ^ n20344;
  assign n20349 = n19100 ^ n18800;
  assign n20350 = n20349 ^ n20008;
  assign n20348 = n19960 ^ n19941;
  assign n20351 = n20350 ^ n20348;
  assign n20410 = n19957 ^ n19946;
  assign n20354 = n19954 ^ n19951;
  assign n20352 = n19086 ^ n18658;
  assign n20353 = n20352 ^ n19883;
  assign n20355 = n20354 ^ n20353;
  assign n20358 = n19725 ^ n19660;
  assign n20356 = n18916 ^ n18629;
  assign n20357 = n20356 ^ n19760;
  assign n20359 = n20358 ^ n20357;
  assign n20362 = n19722 ^ n19662;
  assign n20360 = n18918 ^ n18615;
  assign n20361 = n20360 ^ n19764;
  assign n20363 = n20362 ^ n20361;
  assign n20388 = n19719 ^ n2243;
  assign n20365 = n19770 ^ n18586;
  assign n20366 = n20365 ^ n18923;
  assign n20364 = n19714 ^ n19664;
  assign n20367 = n20366 ^ n20364;
  assign n20378 = n19711 ^ n2223;
  assign n20368 = n19774 ^ n18533;
  assign n20369 = n20368 ^ n18927;
  assign n20371 = n20370 ^ n20369;
  assign n20298 = n18932 ^ n18422;
  assign n20299 = n20298 ^ n19778;
  assign n20301 = n20300 ^ n20299;
  assign n20215 = n19695 ^ n19670;
  assign n20165 = n19738 ^ n18414;
  assign n20166 = n20165 ^ n18940;
  assign n20164 = n19692 ^ n19672;
  assign n20167 = n20166 ^ n20164;
  assign n20157 = n19689 ^ n19677;
  assign n19755 = n19686 ^ n19685;
  assign n19753 = n19637 ^ n18431;
  assign n19754 = n19753 ^ n18413;
  assign n19756 = n19755 ^ n19754;
  assign n20147 = n19680 ^ n19612;
  assign n20116 = n18900 ^ n18439;
  assign n20117 = n20116 ^ n19550;
  assign n20076 = ~n20057 & ~n20070;
  assign n20086 = n18891 ^ n18286;
  assign n20087 = n20086 ^ n16931;
  assign n20081 = n20066 ^ n20062;
  assign n20082 = ~n20067 & n20081;
  assign n20083 = n20082 ^ n20062;
  assign n20085 = n20084 ^ n20083;
  assign n20088 = n20087 ^ n20085;
  assign n20077 = n20068 ^ n20060;
  assign n20078 = n20069 & ~n20077;
  assign n20079 = n20078 ^ n17089;
  assign n20080 = n20079 ^ n17031;
  assign n20089 = n20088 ^ n20080;
  assign n20113 = n20076 & n20089;
  assign n20108 = n18992 ^ n18305;
  assign n20109 = n20108 ^ n16925;
  assign n20105 = n20087 ^ n20084;
  assign n20106 = ~n20085 & ~n20105;
  assign n20107 = n20106 ^ n20087;
  assign n20110 = n20109 ^ n20107;
  assign n20104 = n19442 ^ n19439;
  assign n20111 = n20110 ^ n20104;
  assign n20099 = n20088 ^ n17031;
  assign n20100 = n20088 ^ n20079;
  assign n20101 = ~n20099 & n20100;
  assign n20102 = n20101 ^ n17031;
  assign n20103 = n20102 ^ n17025;
  assign n20112 = n20111 ^ n20103;
  assign n20114 = n20113 ^ n20112;
  assign n20090 = n20089 ^ n20076;
  assign n20073 = n20071 ^ n2486;
  assign n20074 = n20072 & ~n20073;
  assign n20075 = n20074 ^ n2486;
  assign n20091 = n20090 ^ n20075;
  assign n1545 = n1544 ^ x450;
  assign n1546 = n1545 ^ n1514;
  assign n1547 = n1546 ^ x386;
  assign n20092 = n20090 ^ n1547;
  assign n20093 = n20091 & ~n20092;
  assign n20094 = n20093 ^ n1547;
  assign n20098 = n20097 ^ n20094;
  assign n20115 = n20114 ^ n20098;
  assign n20118 = n20117 ^ n20115;
  assign n20137 = n20091 ^ n1547;
  assign n20134 = n20133 ^ n20130;
  assign n20135 = n20131 & n20134;
  assign n20136 = n20135 ^ n20133;
  assign n20138 = n20137 ^ n20136;
  assign n20139 = n19019 ^ n18898;
  assign n20140 = n20139 ^ n18444;
  assign n20141 = n20140 ^ n20137;
  assign n20142 = ~n20138 & ~n20141;
  assign n20143 = n20142 ^ n20140;
  assign n20144 = n20143 ^ n20115;
  assign n20145 = n20118 & n20144;
  assign n20146 = n20145 ^ n20117;
  assign n20148 = n20147 ^ n20146;
  assign n20149 = n19604 ^ n18435;
  assign n20150 = n20149 ^ n19029;
  assign n20151 = n20150 ^ n20147;
  assign n20152 = ~n20148 & n20151;
  assign n20153 = n20152 ^ n20150;
  assign n20154 = n20153 ^ n19755;
  assign n20155 = n19756 & n20154;
  assign n20156 = n20155 ^ n19754;
  assign n20158 = n20157 ^ n20156;
  assign n20159 = n19651 ^ n18410;
  assign n20160 = n20159 ^ n18430;
  assign n20161 = n20160 ^ n20157;
  assign n20162 = ~n20158 & ~n20161;
  assign n20163 = n20162 ^ n20160;
  assign n20212 = n20164 ^ n20163;
  assign n20213 = ~n20167 & ~n20212;
  assign n20214 = n20213 ^ n20166;
  assign n20216 = n20215 ^ n20214;
  assign n20210 = n18936 ^ n17820;
  assign n20211 = n20210 ^ n19780;
  assign n20295 = n20215 ^ n20211;
  assign n20296 = n20216 & n20295;
  assign n20297 = n20296 ^ n20211;
  assign n20317 = n20300 ^ n20297;
  assign n20318 = n20301 & ~n20317;
  assign n20319 = n20318 ^ n20299;
  assign n20321 = n20320 ^ n20319;
  assign n20315 = n19796 ^ n18421;
  assign n20316 = n20315 ^ n19051;
  assign n20372 = n20320 ^ n20316;
  assign n20373 = n20321 & ~n20372;
  assign n20374 = n20373 ^ n20316;
  assign n20375 = n20374 ^ n20370;
  assign n20376 = ~n20371 & ~n20375;
  assign n20377 = n20376 ^ n20369;
  assign n20379 = n20378 ^ n20377;
  assign n20380 = n19061 ^ n18549;
  assign n20381 = n20380 ^ n19751;
  assign n20382 = n20381 ^ n20378;
  assign n20383 = ~n20379 & ~n20382;
  assign n20384 = n20383 ^ n20381;
  assign n20385 = n20384 ^ n20364;
  assign n20386 = n20367 & ~n20385;
  assign n20387 = n20386 ^ n20366;
  assign n20389 = n20388 ^ n20387;
  assign n20390 = n18919 ^ n18601;
  assign n20391 = n20390 ^ n19768;
  assign n20392 = n20391 ^ n20388;
  assign n20393 = ~n20389 & ~n20392;
  assign n20394 = n20393 ^ n20391;
  assign n20395 = n20394 ^ n20362;
  assign n20396 = ~n20363 & ~n20395;
  assign n20397 = n20396 ^ n20361;
  assign n20398 = n20397 ^ n20358;
  assign n20399 = n20359 & ~n20398;
  assign n20400 = n20399 ^ n20357;
  assign n19749 = n19748 ^ n19728;
  assign n20401 = n20400 ^ n19749;
  assign n20402 = n18911 ^ n18644;
  assign n20403 = n20402 ^ n19759;
  assign n20404 = n20403 ^ n19749;
  assign n20405 = n20401 & ~n20404;
  assign n20406 = n20405 ^ n20403;
  assign n20407 = n20406 ^ n20354;
  assign n20408 = ~n20355 & n20407;
  assign n20409 = n20408 ^ n20353;
  assign n20411 = n20410 ^ n20409;
  assign n20412 = n19093 ^ n18775;
  assign n20413 = n20412 ^ n19923;
  assign n20414 = n20413 ^ n20410;
  assign n20415 = n20411 & ~n20414;
  assign n20416 = n20415 ^ n20413;
  assign n20417 = n20416 ^ n20348;
  assign n20418 = n20351 & n20417;
  assign n20419 = n20418 ^ n20350;
  assign n20420 = n20419 ^ n20344;
  assign n20421 = n20347 & ~n20420;
  assign n20422 = n20421 ^ n20346;
  assign n20424 = n20423 ^ n20422;
  assign n20425 = n19466 ^ n18883;
  assign n20426 = n20425 ^ n20047;
  assign n20427 = n20426 ^ n20423;
  assign n20428 = n20424 & ~n20427;
  assign n20429 = n20428 ^ n20426;
  assign n20430 = n20429 ^ n20340;
  assign n20431 = n20343 & ~n20430;
  assign n20432 = n20431 ^ n20342;
  assign n20433 = n20432 ^ n20338;
  assign n20434 = n20339 & n20433;
  assign n20435 = n20434 ^ n20337;
  assign n20335 = n19982 ^ n1085;
  assign n20436 = n20435 ^ n20335;
  assign n20437 = n18808 ^ n18220;
  assign n20438 = n20437 ^ n20104;
  assign n20439 = n20438 ^ n20335;
  assign n20440 = n20436 & n20439;
  assign n20441 = n20440 ^ n20438;
  assign n20334 = n19985 ^ n19933;
  assign n20442 = n20441 ^ n20334;
  assign n20443 = n18840 ^ n18224;
  assign n20444 = n20443 ^ n19508;
  assign n20445 = n20444 ^ n20334;
  assign n20446 = ~n20442 & n20445;
  assign n20447 = n20446 ^ n20444;
  assign n20449 = n20448 ^ n20447;
  assign n20332 = n18891 ^ n18211;
  assign n20333 = n20332 ^ n19513;
  assign n20541 = n20448 ^ n20333;
  assign n20542 = ~n20449 & ~n20541;
  assign n20543 = n20542 ^ n20333;
  assign n20540 = n19993 ^ n19931;
  assign n20544 = n20543 ^ n20540;
  assign n20538 = n18992 ^ n18256;
  assign n20539 = n20538 ^ n19502;
  assign n20695 = n20540 ^ n20539;
  assign n20696 = ~n20544 & ~n20695;
  assign n20697 = n20696 ^ n20539;
  assign n20699 = n20698 ^ n20697;
  assign n20702 = n20701 ^ n20699;
  assign n20545 = n20544 ^ n20539;
  assign n20546 = n20545 ^ n17605;
  assign n20450 = n20449 ^ n20333;
  assign n20451 = n20450 ^ n17609;
  assign n20452 = n20444 ^ n20442;
  assign n20453 = n20452 ^ n17612;
  assign n20454 = n20438 ^ n20436;
  assign n20455 = n20454 ^ n17623;
  assign n20456 = n20432 ^ n20339;
  assign n20457 = n20456 ^ n17618;
  assign n20458 = n20429 ^ n20343;
  assign n20459 = n20458 ^ n18249;
  assign n20460 = n20426 ^ n20424;
  assign n20461 = n20460 ^ n18203;
  assign n20462 = n20419 ^ n20347;
  assign n20463 = n20462 ^ n18185;
  assign n20464 = n20416 ^ n20351;
  assign n20465 = n20464 ^ n18165;
  assign n20466 = n20413 ^ n20411;
  assign n20467 = n20466 ^ n18147;
  assign n20468 = n20406 ^ n20355;
  assign n20469 = n20468 ^ n18009;
  assign n20470 = n20403 ^ n20401;
  assign n20471 = n20470 ^ n17996;
  assign n20472 = n20397 ^ n20359;
  assign n20473 = n20472 ^ n17919;
  assign n20474 = n20394 ^ n20363;
  assign n20475 = n20474 ^ n17828;
  assign n20476 = n20391 ^ n20389;
  assign n20477 = n20476 ^ n17832;
  assign n20478 = n20384 ^ n20367;
  assign n20479 = n20478 ^ n17836;
  assign n20480 = n20381 ^ n20379;
  assign n20481 = n20480 ^ n17841;
  assign n20482 = n20374 ^ n20371;
  assign n20483 = n20482 ^ n17848;
  assign n20322 = n20321 ^ n20316;
  assign n20323 = n20322 ^ n17850;
  assign n20302 = n20301 ^ n20297;
  assign n20303 = n20302 ^ n17891;
  assign n20217 = n20216 ^ n20211;
  assign n20218 = n20217 ^ n17822;
  assign n20168 = n20167 ^ n20163;
  assign n20169 = n20168 ^ n17854;
  assign n20170 = n20160 ^ n20158;
  assign n20171 = n20170 ^ n17860;
  assign n20172 = n20153 ^ n19756;
  assign n20173 = n20172 ^ n17872;
  assign n20174 = n20150 ^ n20148;
  assign n20175 = n20174 ^ n17862;
  assign n20176 = n20143 ^ n20118;
  assign n20177 = n20176 ^ n17807;
  assign n20178 = n20140 ^ n20138;
  assign n20179 = n20178 ^ n17736;
  assign n20189 = n20188 ^ n20180;
  assign n20190 = ~n20181 & n20189;
  assign n20191 = n20190 ^ n17722;
  assign n20192 = n20191 ^ n20178;
  assign n20193 = ~n20179 & n20192;
  assign n20194 = n20193 ^ n17736;
  assign n20195 = n20194 ^ n20176;
  assign n20196 = ~n20177 & n20195;
  assign n20197 = n20196 ^ n17807;
  assign n20198 = n20197 ^ n20174;
  assign n20199 = n20175 & ~n20198;
  assign n20200 = n20199 ^ n17862;
  assign n20201 = n20200 ^ n20172;
  assign n20202 = n20173 & ~n20201;
  assign n20203 = n20202 ^ n17872;
  assign n20204 = n20203 ^ n20170;
  assign n20205 = n20171 & ~n20204;
  assign n20206 = n20205 ^ n17860;
  assign n20207 = n20206 ^ n20168;
  assign n20208 = ~n20169 & n20207;
  assign n20209 = n20208 ^ n17854;
  assign n20292 = n20217 ^ n20209;
  assign n20293 = n20218 & n20292;
  assign n20294 = n20293 ^ n17822;
  assign n20312 = n20302 ^ n20294;
  assign n20313 = n20303 & n20312;
  assign n20314 = n20313 ^ n17891;
  assign n20484 = n20322 ^ n20314;
  assign n20485 = ~n20323 & n20484;
  assign n20486 = n20485 ^ n17850;
  assign n20487 = n20486 ^ n20482;
  assign n20488 = ~n20483 & n20487;
  assign n20489 = n20488 ^ n17848;
  assign n20490 = n20489 ^ n20480;
  assign n20491 = n20481 & ~n20490;
  assign n20492 = n20491 ^ n17841;
  assign n20493 = n20492 ^ n20478;
  assign n20494 = n20479 & ~n20493;
  assign n20495 = n20494 ^ n17836;
  assign n20496 = n20495 ^ n20476;
  assign n20497 = n20477 & n20496;
  assign n20498 = n20497 ^ n17832;
  assign n20499 = n20498 ^ n20474;
  assign n20500 = n20475 & n20499;
  assign n20501 = n20500 ^ n17828;
  assign n20502 = n20501 ^ n20472;
  assign n20503 = n20473 & ~n20502;
  assign n20504 = n20503 ^ n17919;
  assign n20505 = n20504 ^ n20470;
  assign n20506 = n20471 & n20505;
  assign n20507 = n20506 ^ n17996;
  assign n20508 = n20507 ^ n20468;
  assign n20509 = ~n20469 & ~n20508;
  assign n20510 = n20509 ^ n18009;
  assign n20511 = n20510 ^ n20466;
  assign n20512 = ~n20467 & n20511;
  assign n20513 = n20512 ^ n18147;
  assign n20514 = n20513 ^ n20464;
  assign n20515 = n20465 & ~n20514;
  assign n20516 = n20515 ^ n18165;
  assign n20517 = n20516 ^ n20462;
  assign n20518 = ~n20463 & n20517;
  assign n20519 = n20518 ^ n18185;
  assign n20520 = n20519 ^ n20460;
  assign n20521 = n20461 & ~n20520;
  assign n20522 = n20521 ^ n18203;
  assign n20523 = n20522 ^ n20458;
  assign n20524 = n20459 & n20523;
  assign n20525 = n20524 ^ n18249;
  assign n20526 = n20525 ^ n20456;
  assign n20527 = ~n20457 & ~n20526;
  assign n20528 = n20527 ^ n17618;
  assign n20529 = n20528 ^ n20454;
  assign n20530 = n20455 & ~n20529;
  assign n20531 = n20530 ^ n17623;
  assign n20532 = n20531 ^ n20452;
  assign n20533 = n20453 & n20532;
  assign n20534 = n20533 ^ n17612;
  assign n20535 = n20534 ^ n20450;
  assign n20536 = ~n20451 & n20535;
  assign n20537 = n20536 ^ n17609;
  assign n20691 = n20545 ^ n20537;
  assign n20692 = ~n20546 & ~n20691;
  assign n20693 = n20692 ^ n17605;
  assign n20694 = n20693 ^ n16931;
  assign n20703 = n20702 ^ n20694;
  assign n20547 = n20546 ^ n20537;
  assign n20548 = n20531 ^ n20453;
  assign n20549 = n20510 ^ n20467;
  assign n20550 = n20504 ^ n20471;
  assign n20551 = n20501 ^ n20473;
  assign n20552 = n20498 ^ n20475;
  assign n20553 = n20489 ^ n20481;
  assign n20554 = n20486 ^ n20483;
  assign n20304 = n20303 ^ n20294;
  assign n20219 = n20218 ^ n20209;
  assign n20220 = n20206 ^ n20169;
  assign n20221 = n20203 ^ n20171;
  assign n20222 = n20200 ^ n20173;
  assign n20223 = n20197 ^ n20175;
  assign n20224 = n20191 ^ n20179;
  assign n20229 = n20227 & n20228;
  assign n20230 = n20224 & n20229;
  assign n20231 = n20194 ^ n20177;
  assign n20232 = n20230 & n20231;
  assign n20233 = n20223 & ~n20232;
  assign n20234 = ~n20222 & ~n20233;
  assign n20235 = n20221 & ~n20234;
  assign n20236 = ~n20220 & n20235;
  assign n20305 = n20219 & n20236;
  assign n20311 = n20304 & ~n20305;
  assign n20324 = n20323 ^ n20314;
  assign n20555 = ~n20311 & ~n20324;
  assign n20556 = n20554 & ~n20555;
  assign n20557 = n20553 & ~n20556;
  assign n20558 = n20492 ^ n20479;
  assign n20559 = n20557 & n20558;
  assign n20560 = n20495 ^ n20477;
  assign n20561 = n20559 & n20560;
  assign n20562 = ~n20552 & n20561;
  assign n20563 = ~n20551 & ~n20562;
  assign n20564 = ~n20550 & n20563;
  assign n20565 = n20507 ^ n20469;
  assign n20566 = ~n20564 & n20565;
  assign n20567 = ~n20549 & n20566;
  assign n20568 = n20513 ^ n20465;
  assign n20569 = ~n20567 & ~n20568;
  assign n20570 = n20516 ^ n20463;
  assign n20571 = ~n20569 & ~n20570;
  assign n20572 = n20519 ^ n20461;
  assign n20573 = n20571 & n20572;
  assign n20574 = n20522 ^ n20459;
  assign n20575 = ~n20573 & ~n20574;
  assign n20576 = n20525 ^ n20457;
  assign n20577 = ~n20575 & n20576;
  assign n20578 = n20528 ^ n20455;
  assign n20579 = n20577 & n20578;
  assign n20580 = n20548 & n20579;
  assign n20581 = n20534 ^ n20451;
  assign n20582 = ~n20580 & ~n20581;
  assign n20704 = n20547 & ~n20582;
  assign n20770 = n20703 & n20704;
  assign n20767 = n20015 ^ n2289;
  assign n20764 = n18968 ^ n18305;
  assign n20765 = n20764 ^ n19498;
  assign n20761 = n20701 ^ n20698;
  assign n20762 = n20699 & ~n20761;
  assign n20763 = n20762 ^ n20701;
  assign n20766 = n20765 ^ n20763;
  assign n20768 = n20767 ^ n20766;
  assign n20756 = n20702 ^ n16931;
  assign n20757 = n20702 ^ n20693;
  assign n20758 = n20756 & ~n20757;
  assign n20759 = n20758 ^ n16931;
  assign n20760 = n20759 ^ n16925;
  assign n20769 = n20768 ^ n20760;
  assign n20771 = n20770 ^ n20769;
  assign n20705 = n20704 ^ n20703;
  assign n20583 = n20582 ^ n20547;
  assign n20584 = n20583 ^ n2466;
  assign n20683 = n20581 ^ n20580;
  assign n20585 = n20579 ^ n20548;
  assign n2453 = n2379 ^ x485;
  assign n2454 = n2453 ^ n2452;
  assign n2455 = n2454 ^ x421;
  assign n20586 = n20585 ^ n2455;
  assign n20675 = n20578 ^ n20577;
  assign n20587 = n20576 ^ n20575;
  assign n1386 = n1280 ^ x487;
  assign n1387 = n1386 ^ n1380;
  assign n1388 = n1387 ^ x423;
  assign n20588 = n20587 ^ n1388;
  assign n20589 = n20574 ^ n20573;
  assign n20590 = n20589 ^ n1115;
  assign n20664 = n20572 ^ n20571;
  assign n20591 = n20570 ^ n20569;
  assign n20592 = n20591 ^ n951;
  assign n20656 = n20568 ^ n20567;
  assign n20593 = n20566 ^ n20549;
  assign n20594 = n20593 ^ n823;
  assign n20648 = n20565 ^ n20564;
  assign n20595 = n20563 ^ n20550;
  assign n742 = n689 ^ x494;
  assign n746 = n745 ^ n742;
  assign n747 = n746 ^ x430;
  assign n20596 = n20595 ^ n747;
  assign n20597 = n20562 ^ n20551;
  assign n20601 = n20600 ^ n20597;
  assign n20602 = n20561 ^ n20552;
  assign n20606 = n20605 ^ n20602;
  assign n20607 = n20560 ^ n20559;
  assign n20611 = n20610 ^ n20607;
  assign n20628 = n20558 ^ n20557;
  assign n20612 = n20556 ^ n20553;
  assign n20613 = n20612 ^ n596;
  assign n20614 = n20555 ^ n20554;
  assign n20618 = n20617 ^ n20614;
  assign n20325 = n20324 ^ n20311;
  assign n20329 = n20328 ^ n20325;
  assign n20306 = n20305 ^ n20304;
  assign n20237 = n20236 ^ n20219;
  assign n20238 = n20237 ^ n2083;
  assign n20284 = n20235 ^ n20220;
  assign n20239 = n20234 ^ n20221;
  assign n20240 = n20239 ^ n1809;
  assign n20241 = n20233 ^ n20222;
  assign n20242 = n20241 ^ n1794;
  assign n20273 = n20232 ^ n20223;
  assign n20246 = n20231 ^ n20230;
  assign n20247 = n20246 ^ n20245;
  assign n20262 = n20229 ^ n20224;
  assign n20259 = n20258 ^ n20248;
  assign n20260 = n20249 & ~n20259;
  assign n20261 = n20260 ^ n1436;
  assign n20263 = n20262 ^ n20261;
  assign n20267 = n20266 ^ n20262;
  assign n20268 = ~n20263 & n20267;
  assign n20269 = n20268 ^ n20266;
  assign n20270 = n20269 ^ n20246;
  assign n20271 = n20247 & ~n20270;
  assign n20272 = n20271 ^ n20245;
  assign n20274 = n20273 ^ n20272;
  assign n20275 = n20273 ^ n1785;
  assign n20276 = ~n20274 & n20275;
  assign n20277 = n20276 ^ n1785;
  assign n20278 = n20277 ^ n20241;
  assign n20279 = n20242 & ~n20278;
  assign n20280 = n20279 ^ n1794;
  assign n20281 = n20280 ^ n20239;
  assign n20282 = n20240 & ~n20281;
  assign n20283 = n20282 ^ n1809;
  assign n20285 = n20284 ^ n20283;
  assign n20286 = n20284 ^ n1922;
  assign n20287 = ~n20285 & n20286;
  assign n20288 = n20287 ^ n1922;
  assign n20289 = n20288 ^ n20237;
  assign n20290 = ~n20238 & n20289;
  assign n20291 = n20290 ^ n2083;
  assign n20307 = n20306 ^ n20291;
  assign n20308 = n20306 ^ n2072;
  assign n20309 = n20307 & ~n20308;
  assign n20310 = n20309 ^ n2072;
  assign n20619 = n20325 ^ n20310;
  assign n20620 = ~n20329 & n20619;
  assign n20621 = n20620 ^ n20328;
  assign n20622 = n20621 ^ n20614;
  assign n20623 = ~n20618 & n20622;
  assign n20624 = n20623 ^ n20617;
  assign n20625 = n20624 ^ n20612;
  assign n20626 = n20613 & ~n20625;
  assign n20627 = n20626 ^ n596;
  assign n20629 = n20628 ^ n20627;
  assign n20633 = n20632 ^ n20628;
  assign n20634 = n20629 & ~n20633;
  assign n20635 = n20634 ^ n20632;
  assign n20636 = n20635 ^ n20607;
  assign n20637 = ~n20611 & n20636;
  assign n20638 = n20637 ^ n20610;
  assign n20639 = n20638 ^ n20602;
  assign n20640 = n20606 & ~n20639;
  assign n20641 = n20640 ^ n20605;
  assign n20642 = n20641 ^ n20597;
  assign n20643 = n20601 & ~n20642;
  assign n20644 = n20643 ^ n20600;
  assign n20645 = n20644 ^ n20595;
  assign n20646 = ~n20596 & n20645;
  assign n20647 = n20646 ^ n747;
  assign n20649 = n20648 ^ n20647;
  assign n20650 = n20648 ^ n733;
  assign n20651 = ~n20649 & n20650;
  assign n20652 = n20651 ^ n733;
  assign n20653 = n20652 ^ n20593;
  assign n20654 = n20594 & ~n20653;
  assign n20655 = n20654 ^ n823;
  assign n20657 = n20656 ^ n20655;
  assign n20658 = n20656 ^ n832;
  assign n20659 = ~n20657 & n20658;
  assign n20660 = n20659 ^ n832;
  assign n20661 = n20660 ^ n20591;
  assign n20662 = ~n20592 & n20661;
  assign n20663 = n20662 ^ n951;
  assign n20665 = n20664 ^ n20663;
  assign n20666 = n20664 ^ n1370;
  assign n20667 = n20665 & ~n20666;
  assign n20668 = n20667 ^ n1370;
  assign n20669 = n20668 ^ n20589;
  assign n20670 = n20590 & ~n20669;
  assign n20671 = n20670 ^ n1115;
  assign n20672 = n20671 ^ n20587;
  assign n20673 = n20588 & ~n20672;
  assign n20674 = n20673 ^ n1388;
  assign n20676 = n20675 ^ n20674;
  assign n1404 = n1298 ^ x486;
  assign n1405 = n1404 ^ n1304;
  assign n1406 = n1405 ^ x422;
  assign n20677 = n20675 ^ n1406;
  assign n20678 = n20676 & ~n20677;
  assign n20679 = n20678 ^ n1406;
  assign n20680 = n20679 ^ n20585;
  assign n20681 = ~n20586 & n20680;
  assign n20682 = n20681 ^ n2455;
  assign n20684 = n20683 ^ n20682;
  assign n20685 = n20683 ^ n2440;
  assign n20686 = ~n20684 & n20685;
  assign n20687 = n20686 ^ n2440;
  assign n20688 = n20687 ^ n20583;
  assign n20689 = n20584 & ~n20688;
  assign n20690 = n20689 ^ n2466;
  assign n20706 = n20705 ^ n20690;
  assign n20752 = n20705 ^ n2553;
  assign n20753 = n20706 & ~n20752;
  assign n20754 = n20753 ^ n2553;
  assign n2650 = n2646 ^ x481;
  assign n2651 = n2650 ^ n2546;
  assign n2652 = n2651 ^ x417;
  assign n20755 = n20754 ^ n2652;
  assign n20772 = n20771 ^ n20755;
  assign n20722 = n20687 ^ n20584;
  assign n20713 = n19540 ^ n18962;
  assign n20714 = n20713 ^ n20147;
  assign n20715 = n20679 ^ n20586;
  assign n20716 = n20714 & ~n20715;
  assign n20711 = n18957 ^ n18898;
  assign n20712 = n20711 ^ n19755;
  assign n20717 = n20716 ^ n20712;
  assign n20718 = n20684 ^ n2440;
  assign n20719 = n20718 ^ n20712;
  assign n20720 = n20717 & ~n20719;
  assign n20721 = n20720 ^ n20716;
  assign n20723 = n20722 ^ n20721;
  assign n20724 = n19550 ^ n18955;
  assign n20725 = n20724 ^ n20157;
  assign n20726 = n20725 ^ n20722;
  assign n20727 = ~n20723 & n20726;
  assign n20728 = n20727 ^ n20725;
  assign n20708 = n19604 ^ n19019;
  assign n20709 = n20708 ^ n20164;
  assign n20748 = n20728 ^ n20709;
  assign n20707 = n20706 ^ n2553;
  assign n20749 = n20728 ^ n20707;
  assign n20750 = ~n20748 & n20749;
  assign n20751 = n20750 ^ n20709;
  assign n20773 = n20772 ^ n20751;
  assign n20746 = n19637 ^ n18900;
  assign n20747 = n20746 ^ n20215;
  assign n20815 = n20772 ^ n20747;
  assign n20816 = n20773 & ~n20815;
  assign n20817 = n20816 ^ n20747;
  assign n20836 = n20818 ^ n20817;
  assign n20837 = ~n20821 & n20836;
  assign n20838 = n20837 ^ n20820;
  assign n20886 = n20839 ^ n20838;
  assign n20887 = n20842 & n20886;
  assign n20888 = n20887 ^ n20841;
  assign n20890 = n20889 ^ n20888;
  assign n21009 = n20892 ^ n20890;
  assign n21010 = n21009 ^ n18430;
  assign n20843 = n20842 ^ n20838;
  assign n20844 = n20843 ^ n18431;
  assign n20822 = n20821 ^ n20817;
  assign n20823 = n20822 ^ n18435;
  assign n20774 = n20773 ^ n20747;
  assign n20775 = n20774 ^ n18439;
  assign n20710 = n20709 ^ n20707;
  assign n20729 = n20728 ^ n20710;
  assign n20730 = n20729 ^ n18444;
  assign n20731 = n20725 ^ n20723;
  assign n20732 = n20731 ^ n18403;
  assign n20733 = n20715 ^ n20714;
  assign n20734 = n18322 & ~n20733;
  assign n20735 = n20734 ^ n18339;
  assign n20736 = n20718 ^ n20717;
  assign n20737 = n20736 ^ n20734;
  assign n20738 = ~n20735 & ~n20737;
  assign n20739 = n20738 ^ n18339;
  assign n20740 = n20739 ^ n20731;
  assign n20741 = ~n20732 & n20740;
  assign n20742 = n20741 ^ n18403;
  assign n20743 = n20742 ^ n20729;
  assign n20744 = n20730 & n20743;
  assign n20745 = n20744 ^ n18444;
  assign n20812 = n20774 ^ n20745;
  assign n20813 = ~n20775 & ~n20812;
  assign n20814 = n20813 ^ n18439;
  assign n20833 = n20822 ^ n20814;
  assign n20834 = n20823 & n20833;
  assign n20835 = n20834 ^ n18435;
  assign n21011 = n20843 ^ n20835;
  assign n21012 = n20844 & n21011;
  assign n21013 = n21012 ^ n18431;
  assign n21014 = n21013 ^ n21009;
  assign n21015 = n21010 & n21014;
  assign n21016 = n21015 ^ n18430;
  assign n20893 = n20892 ^ n20889;
  assign n20894 = ~n20890 & n20893;
  assign n20895 = n20894 ^ n20892;
  assign n20883 = n19778 ^ n18940;
  assign n20884 = n20883 ^ n20378;
  assign n20882 = n20266 ^ n20263;
  assign n20885 = n20884 ^ n20882;
  assign n21007 = n20895 ^ n20885;
  assign n21008 = n21007 ^ n18414;
  assign n21085 = n21016 ^ n21008;
  assign n20845 = n20844 ^ n20835;
  assign n20776 = n20775 ^ n20745;
  assign n20777 = n20739 ^ n20732;
  assign n20778 = n20733 ^ n18322;
  assign n20779 = n20736 ^ n20735;
  assign n20780 = ~n20778 & ~n20779;
  assign n20781 = n20777 & n20780;
  assign n20782 = n20742 ^ n20730;
  assign n20783 = n20781 & ~n20782;
  assign n20811 = ~n20776 & n20783;
  assign n20824 = n20823 ^ n20814;
  assign n20846 = ~n20811 & n20824;
  assign n21082 = n20845 & ~n20846;
  assign n21083 = n21013 ^ n21010;
  assign n21084 = ~n21082 & n21083;
  assign n21169 = n21085 ^ n21084;
  assign n21161 = n21083 ^ n21082;
  assign n21162 = n21161 ^ n2032;
  assign n20847 = n20846 ^ n20845;
  assign n20848 = n20847 ^ n1694;
  assign n20825 = n20824 ^ n20811;
  assign n20784 = n20783 ^ n20776;
  assign n20785 = n20784 ^ n1601;
  assign n20786 = n20782 ^ n20781;
  assign n20787 = n20786 ^ n1484;
  assign n20788 = n20780 ^ n20777;
  assign n20789 = n20788 ^ n1508;
  assign n20793 = n20778 & n20792;
  assign n20797 = n20796 ^ n20793;
  assign n20798 = n20779 ^ n20778;
  assign n20799 = n20798 ^ n20793;
  assign n20800 = n20797 & ~n20799;
  assign n20801 = n20800 ^ n20796;
  assign n20802 = n20801 ^ n20788;
  assign n20803 = n20789 & ~n20802;
  assign n20804 = n20803 ^ n1508;
  assign n20805 = n20804 ^ n20786;
  assign n20806 = ~n20787 & n20805;
  assign n20807 = n20806 ^ n1484;
  assign n20808 = n20807 ^ n20784;
  assign n20809 = ~n20785 & n20808;
  assign n20810 = n20809 ^ n1601;
  assign n20826 = n20825 ^ n20810;
  assign n20830 = n20829 ^ n20825;
  assign n20831 = ~n20826 & n20830;
  assign n20832 = n20831 ^ n20829;
  assign n21163 = n20847 ^ n20832;
  assign n21164 = ~n20848 & n21163;
  assign n21165 = n21164 ^ n1694;
  assign n21166 = n21165 ^ n21161;
  assign n21167 = n21162 & ~n21166;
  assign n21168 = n21167 ^ n2032;
  assign n21170 = n21169 ^ n21168;
  assign n21171 = n21169 ^ n2038;
  assign n21172 = ~n21170 & n21171;
  assign n21173 = n21172 ^ n2038;
  assign n21086 = n21084 & ~n21085;
  assign n21017 = n21016 ^ n21007;
  assign n21018 = n21008 & n21017;
  assign n21019 = n21018 ^ n18414;
  assign n20901 = n19796 ^ n18936;
  assign n20902 = n20901 ^ n20364;
  assign n20899 = n20269 ^ n20247;
  assign n20896 = n20895 ^ n20882;
  assign n20897 = ~n20885 & ~n20896;
  assign n20898 = n20897 ^ n20884;
  assign n20900 = n20899 ^ n20898;
  assign n21005 = n20902 ^ n20900;
  assign n21006 = n21005 ^ n17820;
  assign n21081 = n21019 ^ n21006;
  assign n21159 = n21086 ^ n21081;
  assign n21160 = n21159 ^ n2053;
  assign n21631 = n21173 ^ n21160;
  assign n20934 = n20288 ^ n20238;
  assign n22599 = n21631 ^ n20934;
  assign n21360 = n20300 ^ n19604;
  assign n21361 = n21360 ^ n20882;
  assign n21318 = n20668 ^ n20590;
  assign n21268 = n20660 ^ n20592;
  assign n21249 = n20657 ^ n832;
  assign n21120 = n20652 ^ n20594;
  assign n21070 = n20649 ^ n733;
  assign n20975 = n20644 ^ n20596;
  assign n20863 = n20066 ^ n19236;
  assign n20864 = n20863 ^ n20334;
  assign n20862 = n20641 ^ n20601;
  assign n20865 = n20864 ^ n20862;
  assign n20867 = n20047 ^ n19100;
  assign n20868 = n20867 ^ n20335;
  assign n20866 = n20638 ^ n20606;
  assign n20869 = n20868 ^ n20866;
  assign n20962 = n20635 ^ n20611;
  assign n20871 = n20008 ^ n19086;
  assign n20872 = n20871 ^ n20340;
  assign n20870 = n20632 ^ n20629;
  assign n20873 = n20872 ^ n20870;
  assign n20877 = n20621 ^ n20618;
  assign n20875 = n19883 ^ n18916;
  assign n20876 = n20875 ^ n20344;
  assign n20878 = n20877 ^ n20876;
  assign n20879 = n19759 ^ n18918;
  assign n20880 = n20879 ^ n20348;
  assign n20330 = n20329 ^ n20310;
  assign n20881 = n20880 ^ n20330;
  assign n20927 = n20285 ^ n1922;
  assign n20920 = n20280 ^ n20240;
  assign n20913 = n20277 ^ n20242;
  assign n20906 = n20274 ^ n1785;
  assign n20903 = n20902 ^ n20899;
  assign n20904 = n20900 & ~n20903;
  assign n20905 = n20904 ^ n20902;
  assign n20907 = n20906 ^ n20905;
  assign n20908 = n19774 ^ n18932;
  assign n20909 = n20908 ^ n20388;
  assign n20910 = n20909 ^ n20906;
  assign n20911 = n20907 & ~n20910;
  assign n20912 = n20911 ^ n20909;
  assign n20914 = n20913 ^ n20912;
  assign n20915 = n19751 ^ n19051;
  assign n20916 = n20915 ^ n20362;
  assign n20917 = n20916 ^ n20913;
  assign n20918 = n20914 & n20917;
  assign n20919 = n20918 ^ n20916;
  assign n20921 = n20920 ^ n20919;
  assign n20922 = n19770 ^ n18927;
  assign n20923 = n20922 ^ n20358;
  assign n20924 = n20923 ^ n20920;
  assign n20925 = ~n20921 & ~n20924;
  assign n20926 = n20925 ^ n20923;
  assign n20928 = n20927 ^ n20926;
  assign n20929 = n19768 ^ n19061;
  assign n20930 = n20929 ^ n19749;
  assign n20931 = n20930 ^ n20927;
  assign n20932 = n20928 & n20931;
  assign n20933 = n20932 ^ n20930;
  assign n20935 = n20934 ^ n20933;
  assign n20936 = n19764 ^ n18923;
  assign n20937 = n20936 ^ n20354;
  assign n20938 = n20937 ^ n20934;
  assign n20939 = n20935 & n20938;
  assign n20940 = n20939 ^ n20937;
  assign n20852 = n20307 ^ n2072;
  assign n20941 = n20940 ^ n20852;
  assign n20942 = n19760 ^ n18919;
  assign n20943 = n20942 ^ n20410;
  assign n20944 = n20943 ^ n20852;
  assign n20945 = ~n20941 & ~n20944;
  assign n20946 = n20945 ^ n20943;
  assign n20947 = n20946 ^ n20330;
  assign n20948 = n20881 & n20947;
  assign n20949 = n20948 ^ n20880;
  assign n20950 = n20949 ^ n20877;
  assign n20951 = n20878 & ~n20950;
  assign n20952 = n20951 ^ n20876;
  assign n20874 = n20624 ^ n20613;
  assign n20953 = n20952 ^ n20874;
  assign n20954 = n19923 ^ n18911;
  assign n20955 = n20954 ^ n20423;
  assign n20956 = n20955 ^ n20874;
  assign n20957 = n20953 & ~n20956;
  assign n20958 = n20957 ^ n20955;
  assign n20959 = n20958 ^ n20870;
  assign n20960 = ~n20873 & ~n20959;
  assign n20961 = n20960 ^ n20872;
  assign n20963 = n20962 ^ n20961;
  assign n20964 = n20028 ^ n19093;
  assign n20965 = n20964 ^ n20338;
  assign n20966 = n20965 ^ n20962;
  assign n20967 = n20963 & n20966;
  assign n20968 = n20967 ^ n20965;
  assign n20969 = n20968 ^ n20866;
  assign n20970 = ~n20869 & n20969;
  assign n20971 = n20970 ^ n20868;
  assign n20972 = n20971 ^ n20862;
  assign n20973 = n20865 & n20972;
  assign n20974 = n20973 ^ n20864;
  assign n20976 = n20975 ^ n20974;
  assign n20860 = n20084 ^ n19466;
  assign n20861 = n20860 ^ n20448;
  assign n21067 = n20975 ^ n20861;
  assign n21068 = n20976 & n21067;
  assign n21069 = n21068 ^ n20861;
  assign n21071 = n21070 ^ n21069;
  assign n21065 = n20104 ^ n19493;
  assign n21066 = n21065 ^ n20540;
  assign n21117 = n21070 ^ n21066;
  assign n21118 = n21071 & n21117;
  assign n21119 = n21118 ^ n21066;
  assign n21121 = n21120 ^ n21119;
  assign n21115 = n19508 ^ n18782;
  assign n21116 = n21115 ^ n20698;
  assign n21246 = n21120 ^ n21116;
  assign n21247 = ~n21121 & n21246;
  assign n21248 = n21247 ^ n21116;
  assign n21250 = n21249 ^ n21248;
  assign n21244 = n19513 ^ n18808;
  assign n21245 = n21244 ^ n20767;
  assign n21265 = n21249 ^ n21245;
  assign n21266 = ~n21250 & ~n21265;
  assign n21267 = n21266 ^ n21245;
  assign n21269 = n21268 ^ n21267;
  assign n21263 = n19502 ^ n18840;
  assign n21264 = n21263 ^ n20121;
  assign n21293 = n21268 ^ n21264;
  assign n21294 = ~n21269 & n21293;
  assign n21295 = n21294 ^ n21264;
  assign n21292 = n20665 ^ n1370;
  assign n21296 = n21295 ^ n21292;
  assign n21290 = n19520 ^ n18891;
  assign n21291 = n21290 ^ n20126;
  assign n21315 = n21292 ^ n21291;
  assign n21316 = ~n21296 & n21315;
  assign n21317 = n21316 ^ n21291;
  assign n21319 = n21318 ^ n21317;
  assign n21313 = n19498 ^ n18992;
  assign n21314 = n21313 ^ n20130;
  assign n21320 = n21319 ^ n21314;
  assign n21321 = n21320 ^ n18256;
  assign n21297 = n21296 ^ n21291;
  assign n21298 = n21297 ^ n18211;
  assign n21270 = n21269 ^ n21264;
  assign n21271 = n21270 ^ n18224;
  assign n21251 = n21250 ^ n21245;
  assign n21252 = n21251 ^ n18220;
  assign n21122 = n21121 ^ n21116;
  assign n21123 = n21122 ^ n18215;
  assign n21072 = n21071 ^ n21066;
  assign n21073 = n21072 ^ n18984;
  assign n20977 = n20976 ^ n20861;
  assign n20978 = n20977 ^ n18883;
  assign n20979 = n20971 ^ n20865;
  assign n20980 = n20979 ^ n18834;
  assign n20981 = n20968 ^ n20869;
  assign n20982 = n20981 ^ n18800;
  assign n20983 = n20965 ^ n20963;
  assign n20984 = n20983 ^ n18775;
  assign n20985 = n20958 ^ n20873;
  assign n20986 = n20985 ^ n18658;
  assign n20987 = n20955 ^ n20953;
  assign n20988 = n20987 ^ n18644;
  assign n20989 = n20949 ^ n20878;
  assign n20990 = n20989 ^ n18629;
  assign n20991 = n20946 ^ n20881;
  assign n20992 = n20991 ^ n18615;
  assign n20993 = n20943 ^ n20941;
  assign n20994 = n20993 ^ n18601;
  assign n20995 = n20937 ^ n20935;
  assign n20996 = n20995 ^ n18586;
  assign n20997 = n20930 ^ n20928;
  assign n20998 = n20997 ^ n18549;
  assign n20999 = n20923 ^ n20921;
  assign n21000 = n20999 ^ n18533;
  assign n21001 = n20916 ^ n20914;
  assign n21002 = n21001 ^ n18421;
  assign n21003 = n20909 ^ n20907;
  assign n21004 = n21003 ^ n18422;
  assign n21020 = n21019 ^ n21005;
  assign n21021 = n21006 & n21020;
  assign n21022 = n21021 ^ n17820;
  assign n21023 = n21022 ^ n21003;
  assign n21024 = ~n21004 & ~n21023;
  assign n21025 = n21024 ^ n18422;
  assign n21026 = n21025 ^ n21001;
  assign n21027 = ~n21002 & ~n21026;
  assign n21028 = n21027 ^ n18421;
  assign n21029 = n21028 ^ n20999;
  assign n21030 = n21000 & n21029;
  assign n21031 = n21030 ^ n18533;
  assign n21032 = n21031 ^ n20997;
  assign n21033 = n20998 & ~n21032;
  assign n21034 = n21033 ^ n18549;
  assign n21035 = n21034 ^ n20995;
  assign n21036 = n20996 & n21035;
  assign n21037 = n21036 ^ n18586;
  assign n21038 = n21037 ^ n20993;
  assign n21039 = n20994 & ~n21038;
  assign n21040 = n21039 ^ n18601;
  assign n21041 = n21040 ^ n20991;
  assign n21042 = n20992 & ~n21041;
  assign n21043 = n21042 ^ n18615;
  assign n21044 = n21043 ^ n20989;
  assign n21045 = n20990 & n21044;
  assign n21046 = n21045 ^ n18629;
  assign n21047 = n21046 ^ n20987;
  assign n21048 = n20988 & n21047;
  assign n21049 = n21048 ^ n18644;
  assign n21050 = n21049 ^ n20985;
  assign n21051 = n20986 & ~n21050;
  assign n21052 = n21051 ^ n18658;
  assign n21053 = n21052 ^ n20983;
  assign n21054 = n20984 & ~n21053;
  assign n21055 = n21054 ^ n18775;
  assign n21056 = n21055 ^ n20981;
  assign n21057 = n20982 & ~n21056;
  assign n21058 = n21057 ^ n18800;
  assign n21059 = n21058 ^ n20979;
  assign n21060 = ~n20980 & n21059;
  assign n21061 = n21060 ^ n18834;
  assign n21062 = n21061 ^ n20977;
  assign n21063 = ~n20978 & ~n21062;
  assign n21064 = n21063 ^ n18883;
  assign n21112 = n21072 ^ n21064;
  assign n21113 = ~n21073 & ~n21112;
  assign n21114 = n21113 ^ n18984;
  assign n21241 = n21122 ^ n21114;
  assign n21242 = ~n21123 & ~n21241;
  assign n21243 = n21242 ^ n18215;
  assign n21260 = n21251 ^ n21243;
  assign n21261 = n21252 & ~n21260;
  assign n21262 = n21261 ^ n18220;
  assign n21287 = n21270 ^ n21262;
  assign n21288 = ~n21271 & ~n21287;
  assign n21289 = n21288 ^ n18224;
  assign n21310 = n21297 ^ n21289;
  assign n21311 = ~n21298 & n21310;
  assign n21312 = n21311 ^ n18211;
  assign n21322 = n21321 ^ n21312;
  assign n21299 = n21298 ^ n21289;
  assign n21272 = n21271 ^ n21262;
  assign n21253 = n21252 ^ n21243;
  assign n21074 = n21073 ^ n21064;
  assign n21075 = n21058 ^ n20980;
  assign n21076 = n21055 ^ n20982;
  assign n21077 = n21046 ^ n20988;
  assign n21078 = n21040 ^ n20992;
  assign n21079 = n21031 ^ n20998;
  assign n21080 = n21022 ^ n21004;
  assign n21087 = n21081 & n21086;
  assign n21088 = ~n21080 & ~n21087;
  assign n21089 = n21025 ^ n21002;
  assign n21090 = ~n21088 & ~n21089;
  assign n21091 = n21028 ^ n21000;
  assign n21092 = ~n21090 & n21091;
  assign n21093 = n21079 & ~n21092;
  assign n21094 = n21034 ^ n18586;
  assign n21095 = n21094 ^ n20995;
  assign n21096 = n21093 & n21095;
  assign n21097 = n21037 ^ n20994;
  assign n21098 = n21096 & ~n21097;
  assign n21099 = ~n21078 & n21098;
  assign n21100 = n21043 ^ n20990;
  assign n21101 = ~n21099 & n21100;
  assign n21102 = ~n21077 & n21101;
  assign n21103 = n21049 ^ n20986;
  assign n21104 = ~n21102 & ~n21103;
  assign n21105 = n21052 ^ n20984;
  assign n21106 = n21104 & ~n21105;
  assign n21107 = n21076 & ~n21106;
  assign n21108 = n21075 & ~n21107;
  assign n21109 = n21061 ^ n20978;
  assign n21110 = n21108 & n21109;
  assign n21111 = n21074 & ~n21110;
  assign n21124 = n21123 ^ n21114;
  assign n21254 = ~n21111 & n21124;
  assign n21273 = n21253 & n21254;
  assign n21300 = ~n21272 & n21273;
  assign n21323 = ~n21299 & ~n21300;
  assign n21352 = n21322 & ~n21323;
  assign n21348 = n18999 ^ n18905;
  assign n21349 = n21348 ^ n20137;
  assign n21346 = n20671 ^ n20588;
  assign n21343 = n21318 ^ n21314;
  assign n21344 = n21319 & n21343;
  assign n21345 = n21344 ^ n21314;
  assign n21347 = n21346 ^ n21345;
  assign n21350 = n21349 ^ n21347;
  assign n21339 = n21320 ^ n21312;
  assign n21340 = ~n21321 & n21339;
  assign n21341 = n21340 ^ n18256;
  assign n21342 = n21341 ^ n18286;
  assign n21351 = n21350 ^ n21342;
  assign n21353 = n21352 ^ n21351;
  assign n21324 = n21323 ^ n21322;
  assign n21301 = n21300 ^ n21299;
  assign n21274 = n21273 ^ n21272;
  assign n21255 = n21254 ^ n21253;
  assign n21125 = n21124 ^ n21111;
  assign n21126 = n21125 ^ n1228;
  assign n21127 = n21110 ^ n21074;
  assign n1217 = n1207 ^ n1120;
  assign n1218 = n1217 ^ n1055;
  assign n1219 = n1218 ^ x456;
  assign n21128 = n21127 ^ n1219;
  assign n21230 = n21109 ^ n21108;
  assign n21129 = n21107 ^ n21075;
  assign n937 = n896 ^ n867;
  assign n938 = n937 ^ n918;
  assign n939 = n938 ^ x458;
  assign n21130 = n21129 ^ n939;
  assign n21222 = n21106 ^ n21076;
  assign n21131 = n21105 ^ n21104;
  assign n21132 = n21131 ^ n928;
  assign n21211 = n21103 ^ n21102;
  assign n21133 = n21101 ^ n21077;
  assign n21137 = n21136 ^ n21133;
  assign n21138 = n21100 ^ n21099;
  assign n21139 = n21138 ^ n539;
  assign n21141 = n19321 ^ n12450;
  assign n21142 = n21141 ^ n625;
  assign n21143 = n21142 ^ x464;
  assign n21140 = n21098 ^ n21078;
  assign n21144 = n21143 ^ n21140;
  assign n21145 = n21097 ^ n21096;
  assign n21146 = n21145 ^ n621;
  assign n21191 = n21095 ^ n21093;
  assign n21147 = n21092 ^ n21079;
  assign n21151 = n21150 ^ n21147;
  assign n21152 = n21091 ^ n21090;
  assign n21156 = n21155 ^ n21152;
  assign n21157 = n21089 ^ n21088;
  assign n21158 = n21157 ^ n2214;
  assign n21177 = n21087 ^ n21080;
  assign n21174 = n21173 ^ n21159;
  assign n21175 = ~n21160 & n21174;
  assign n21176 = n21175 ^ n2053;
  assign n21178 = n21177 ^ n21176;
  assign n21179 = n21177 ^ n2199;
  assign n21180 = ~n21178 & n21179;
  assign n21181 = n21180 ^ n2199;
  assign n21182 = n21181 ^ n21157;
  assign n21183 = ~n21158 & n21182;
  assign n21184 = n21183 ^ n2214;
  assign n21185 = n21184 ^ n21152;
  assign n21186 = ~n21156 & n21185;
  assign n21187 = n21186 ^ n21155;
  assign n21188 = n21187 ^ n21147;
  assign n21189 = n21151 & ~n21188;
  assign n21190 = n21189 ^ n21150;
  assign n21192 = n21191 ^ n21190;
  assign n21196 = n21195 ^ n21191;
  assign n21197 = n21192 & ~n21196;
  assign n21198 = n21197 ^ n21195;
  assign n21199 = n21198 ^ n21145;
  assign n21200 = n21146 & ~n21199;
  assign n21201 = n21200 ^ n621;
  assign n21202 = n21201 ^ n21140;
  assign n21203 = n21144 & ~n21202;
  assign n21204 = n21203 ^ n21143;
  assign n21205 = n21204 ^ n21138;
  assign n21206 = ~n21139 & n21205;
  assign n21207 = n21206 ^ n539;
  assign n21208 = n21207 ^ n21133;
  assign n21209 = ~n21137 & n21208;
  assign n21210 = n21209 ^ n21136;
  assign n21212 = n21211 ^ n21210;
  assign n21216 = n21215 ^ n21211;
  assign n21217 = n21212 & ~n21216;
  assign n21218 = n21217 ^ n21215;
  assign n21219 = n21218 ^ n21131;
  assign n21220 = n21132 & ~n21219;
  assign n21221 = n21220 ^ n928;
  assign n21223 = n21222 ^ n21221;
  assign n21224 = n21222 ^ n914;
  assign n21225 = n21223 & ~n21224;
  assign n21226 = n21225 ^ n914;
  assign n21227 = n21226 ^ n21129;
  assign n21228 = n21130 & ~n21227;
  assign n21229 = n21228 ^ n939;
  assign n21231 = n21230 ^ n21229;
  assign n21232 = n21230 ^ n1051;
  assign n21233 = n21231 & ~n21232;
  assign n21234 = n21233 ^ n1051;
  assign n21235 = n21234 ^ n21127;
  assign n21236 = ~n21128 & n21235;
  assign n21237 = n21236 ^ n1219;
  assign n21238 = n21237 ^ n21125;
  assign n21239 = n21126 & ~n21238;
  assign n21240 = n21239 ^ n1228;
  assign n21256 = n21255 ^ n21240;
  assign n2268 = n2267 ^ n1311;
  assign n2272 = n2271 ^ n2268;
  assign n2273 = n2272 ^ x454;
  assign n21257 = n21255 ^ n2273;
  assign n21258 = n21256 & ~n21257;
  assign n21259 = n21258 ^ n2273;
  assign n21275 = n21274 ^ n21259;
  assign n21276 = n19442 ^ n1535;
  assign n21277 = n21276 ^ n2281;
  assign n21278 = n21277 ^ x453;
  assign n21284 = n21278 ^ n21274;
  assign n21285 = ~n21275 & n21284;
  assign n21286 = n21285 ^ n21278;
  assign n21302 = n21301 ^ n21286;
  assign n2361 = n2360 ^ n2318;
  assign n2362 = n2361 ^ n2351;
  assign n2363 = n2362 ^ x452;
  assign n21307 = n21301 ^ n2363;
  assign n21308 = ~n21302 & n21307;
  assign n21309 = n21308 ^ n2363;
  assign n21325 = n21324 ^ n21309;
  assign n21326 = n2595 ^ n2522;
  assign n21327 = n21326 ^ n1541;
  assign n21328 = n21327 ^ x451;
  assign n21336 = n21328 ^ n21324;
  assign n21337 = ~n21325 & n21336;
  assign n21338 = n21337 ^ n21328;
  assign n21354 = n21353 ^ n21338;
  assign n21358 = n21357 ^ n21354;
  assign n21329 = n21328 ^ n21325;
  assign n21279 = n21278 ^ n21275;
  assign n21280 = n20157 ^ n19540;
  assign n21281 = n21280 ^ n20818;
  assign n21282 = n21279 & n21281;
  assign n20858 = n20164 ^ n18898;
  assign n20859 = n20858 ^ n20839;
  assign n21283 = n21282 ^ n20859;
  assign n21303 = n21302 ^ n2363;
  assign n21304 = n21303 ^ n20859;
  assign n21305 = ~n21283 & n21304;
  assign n21306 = n21305 ^ n21282;
  assign n21330 = n21329 ^ n21306;
  assign n21331 = n20215 ^ n19550;
  assign n21332 = n21331 ^ n20889;
  assign n21333 = n21332 ^ n21329;
  assign n21334 = ~n21330 & ~n21333;
  assign n21335 = n21334 ^ n21332;
  assign n21359 = n21358 ^ n21335;
  assign n21447 = n21361 ^ n21359;
  assign n21448 = n21447 ^ n19019;
  assign n21449 = n21332 ^ n21330;
  assign n21450 = n21449 ^ n18955;
  assign n21451 = n21281 ^ n21279;
  assign n21452 = ~n18962 & n21451;
  assign n21453 = n21452 ^ n18957;
  assign n21454 = n21303 ^ n21283;
  assign n21455 = n21454 ^ n21452;
  assign n21456 = n21453 & n21455;
  assign n21457 = n21456 ^ n18957;
  assign n21458 = n21457 ^ n21449;
  assign n21459 = ~n21450 & n21458;
  assign n21460 = n21459 ^ n18955;
  assign n21461 = n21460 ^ n21447;
  assign n21462 = ~n21448 & n21461;
  assign n21463 = n21462 ^ n19019;
  assign n21390 = n20320 ^ n19637;
  assign n21391 = n21390 ^ n20899;
  assign n21386 = n21351 & n21352;
  assign n21383 = n20676 ^ n1406;
  assign n21380 = n18968 ^ n18903;
  assign n21381 = n21380 ^ n20115;
  assign n21377 = n21349 ^ n21346;
  assign n21378 = ~n21347 & n21377;
  assign n21379 = n21378 ^ n21349;
  assign n21382 = n21381 ^ n21379;
  assign n21384 = n21383 ^ n21382;
  assign n21372 = n21350 ^ n18286;
  assign n21373 = n21350 ^ n21341;
  assign n21374 = ~n21372 & ~n21373;
  assign n21375 = n21374 ^ n18286;
  assign n21376 = n21375 ^ n18305;
  assign n21385 = n21384 ^ n21376;
  assign n21387 = n21386 ^ n21385;
  assign n21365 = n21357 ^ n21353;
  assign n21366 = n21354 & ~n21365;
  assign n21367 = n21366 ^ n21357;
  assign n21371 = n21370 ^ n21367;
  assign n21388 = n21387 ^ n21371;
  assign n21362 = n21361 ^ n21358;
  assign n21363 = ~n21359 & n21362;
  assign n21364 = n21363 ^ n21361;
  assign n21389 = n21388 ^ n21364;
  assign n21445 = n21391 ^ n21389;
  assign n21446 = n21445 ^ n18900;
  assign n21501 = n21463 ^ n21446;
  assign n21502 = n21460 ^ n21448;
  assign n21503 = n21457 ^ n21450;
  assign n21504 = n21451 ^ n18962;
  assign n21505 = n21454 ^ n21453;
  assign n21506 = ~n21504 & ~n21505;
  assign n21507 = ~n21503 & n21506;
  assign n21508 = ~n21502 & n21507;
  assign n21509 = ~n21501 & n21508;
  assign n21464 = n21463 ^ n21445;
  assign n21465 = ~n21446 & n21464;
  assign n21466 = n21465 ^ n18900;
  assign n21397 = n20370 ^ n19651;
  assign n21398 = n21397 ^ n20906;
  assign n21395 = n20792 ^ n20778;
  assign n21392 = n21391 ^ n21388;
  assign n21393 = n21389 & n21392;
  assign n21394 = n21393 ^ n21391;
  assign n21396 = n21395 ^ n21394;
  assign n21443 = n21398 ^ n21396;
  assign n21444 = n21443 ^ n19029;
  assign n21510 = n21466 ^ n21444;
  assign n21511 = ~n21509 & n21510;
  assign n21467 = n21466 ^ n21443;
  assign n21468 = ~n21444 & ~n21467;
  assign n21469 = n21468 ^ n19029;
  assign n21403 = n20378 ^ n19738;
  assign n21404 = n21403 ^ n20913;
  assign n21399 = n21398 ^ n21395;
  assign n21400 = ~n21396 & n21399;
  assign n21401 = n21400 ^ n21398;
  assign n20857 = n20798 ^ n20797;
  assign n21402 = n21401 ^ n20857;
  assign n21441 = n21404 ^ n21402;
  assign n21442 = n21441 ^ n18413;
  assign n21500 = n21469 ^ n21442;
  assign n21552 = n21511 ^ n21500;
  assign n21553 = n21552 ^ n1765;
  assign n21587 = n21510 ^ n21509;
  assign n21554 = n21508 ^ n21501;
  assign n21555 = n21554 ^ n1667;
  assign n21559 = n21507 ^ n21502;
  assign n21560 = n21559 ^ n21558;
  assign n21561 = n21506 ^ n21503;
  assign n21565 = n21564 ^ n21561;
  assign n21569 = n21504 & n21568;
  assign n21573 = n21572 ^ n21569;
  assign n21574 = n21505 ^ n21504;
  assign n21575 = n21574 ^ n21572;
  assign n21576 = n21573 & ~n21575;
  assign n21577 = n21576 ^ n21569;
  assign n21578 = n21577 ^ n21561;
  assign n21579 = ~n21565 & n21578;
  assign n21580 = n21579 ^ n21564;
  assign n21581 = n21580 ^ n21559;
  assign n21582 = ~n21560 & n21581;
  assign n21583 = n21582 ^ n21558;
  assign n21584 = n21583 ^ n21554;
  assign n21585 = ~n21555 & n21584;
  assign n21586 = n21585 ^ n1667;
  assign n21588 = n21587 ^ n21586;
  assign n21589 = n21587 ^ n1676;
  assign n21590 = ~n21588 & n21589;
  assign n21591 = n21590 ^ n1676;
  assign n21592 = n21591 ^ n21552;
  assign n21593 = n21553 & ~n21592;
  assign n21594 = n21593 ^ n1765;
  assign n21470 = n21469 ^ n21441;
  assign n21471 = n21442 & ~n21470;
  assign n21472 = n21471 ^ n18413;
  assign n21409 = n20364 ^ n19780;
  assign n21410 = n21409 ^ n20920;
  assign n21405 = n21404 ^ n20857;
  assign n21406 = ~n21402 & ~n21405;
  assign n21407 = n21406 ^ n21404;
  assign n20856 = n20801 ^ n20789;
  assign n21408 = n21407 ^ n20856;
  assign n21439 = n21410 ^ n21408;
  assign n21440 = n21439 ^ n18410;
  assign n21513 = n21472 ^ n21440;
  assign n21512 = ~n21500 & ~n21511;
  assign n21550 = n21513 ^ n21512;
  assign n21551 = n21550 ^ n1774;
  assign n21663 = n21594 ^ n21551;
  assign n22600 = n22599 ^ n21663;
  assign n21931 = n21226 ^ n21130;
  assign n21911 = n21223 ^ n914;
  assign n21809 = n20121 ^ n19508;
  assign n21810 = n21809 ^ n21346;
  assign n21808 = n21218 ^ n21132;
  assign n21811 = n21810 ^ n21808;
  assign n21749 = n20767 ^ n20104;
  assign n21750 = n21749 ^ n21318;
  assign n21748 = n21215 ^ n21212;
  assign n21751 = n21750 ^ n21748;
  assign n21741 = n21207 ^ n21137;
  assign n21687 = n20540 ^ n20066;
  assign n21688 = n21687 ^ n21268;
  assign n21646 = n21204 ^ n21139;
  assign n21689 = n21688 ^ n21646;
  assign n21692 = n21201 ^ n21144;
  assign n21690 = n20448 ^ n20047;
  assign n21691 = n21690 ^ n21249;
  assign n21693 = n21692 ^ n21691;
  assign n21695 = n20335 ^ n20008;
  assign n21696 = n21695 ^ n21070;
  assign n21694 = n21195 ^ n21192;
  assign n21697 = n21696 ^ n21694;
  assign n21698 = n20340 ^ n19883;
  assign n21699 = n21698 ^ n20862;
  assign n21661 = n21184 ^ n21156;
  assign n21700 = n21699 ^ n21661;
  assign n21702 = n20423 ^ n19759;
  assign n21703 = n21702 ^ n20866;
  assign n21701 = n21181 ^ n21158;
  assign n21704 = n21703 ^ n21701;
  assign n21632 = n20348 ^ n19764;
  assign n21633 = n21632 ^ n20870;
  assign n21634 = n21633 ^ n21631;
  assign n21492 = n20354 ^ n19770;
  assign n21493 = n21492 ^ n20877;
  assign n21491 = n21165 ^ n21162;
  assign n21494 = n21493 ^ n21491;
  assign n20851 = n20358 ^ n19774;
  assign n20853 = n20852 ^ n20851;
  assign n20850 = n20829 ^ n20826;
  assign n20854 = n20853 ^ n20850;
  assign n21420 = n20807 ^ n20785;
  assign n21411 = n21410 ^ n20856;
  assign n21412 = n21408 & n21411;
  assign n21413 = n21412 ^ n21410;
  assign n20855 = n20804 ^ n20787;
  assign n21414 = n21413 ^ n20855;
  assign n21415 = n20388 ^ n19778;
  assign n21416 = n21415 ^ n20927;
  assign n21417 = n21416 ^ n20855;
  assign n21418 = n21414 & ~n21417;
  assign n21419 = n21418 ^ n21416;
  assign n21421 = n21420 ^ n21419;
  assign n21422 = n20362 ^ n19796;
  assign n21423 = n21422 ^ n20934;
  assign n21424 = n21423 ^ n21420;
  assign n21425 = n21421 & n21424;
  assign n21426 = n21425 ^ n21423;
  assign n21427 = n21426 ^ n20850;
  assign n21428 = ~n20854 & n21427;
  assign n21429 = n21428 ^ n20853;
  assign n20849 = n20848 ^ n20832;
  assign n21430 = n21429 ^ n20849;
  assign n19752 = n19751 ^ n19749;
  assign n20331 = n20330 ^ n19752;
  assign n21488 = n20849 ^ n20331;
  assign n21489 = ~n21430 & ~n21488;
  assign n21490 = n21489 ^ n20331;
  assign n21528 = n21491 ^ n21490;
  assign n21529 = ~n21494 & ~n21528;
  assign n21530 = n21529 ^ n21493;
  assign n21527 = n21170 ^ n2038;
  assign n21531 = n21530 ^ n21527;
  assign n21525 = n20410 ^ n19768;
  assign n21526 = n21525 ^ n20874;
  assign n21628 = n21527 ^ n21526;
  assign n21629 = n21531 & ~n21628;
  assign n21630 = n21629 ^ n21526;
  assign n21705 = n21631 ^ n21630;
  assign n21706 = n21634 & ~n21705;
  assign n21707 = n21706 ^ n21633;
  assign n21666 = n21178 ^ n2199;
  assign n21708 = n21707 ^ n21666;
  assign n21709 = n20344 ^ n19760;
  assign n21710 = n21709 ^ n20962;
  assign n21711 = n21710 ^ n21666;
  assign n21712 = n21708 & n21711;
  assign n21713 = n21712 ^ n21710;
  assign n21714 = n21713 ^ n21701;
  assign n21715 = n21704 & n21714;
  assign n21716 = n21715 ^ n21703;
  assign n21717 = n21716 ^ n21661;
  assign n21718 = ~n21700 & ~n21717;
  assign n21719 = n21718 ^ n21699;
  assign n21656 = n21187 ^ n21151;
  assign n21720 = n21719 ^ n21656;
  assign n21721 = n20338 ^ n19923;
  assign n21722 = n21721 ^ n20975;
  assign n21723 = n21722 ^ n21656;
  assign n21724 = ~n21720 & ~n21723;
  assign n21725 = n21724 ^ n21722;
  assign n21726 = n21725 ^ n21694;
  assign n21727 = n21697 & ~n21726;
  assign n21728 = n21727 ^ n21696;
  assign n21652 = n21198 ^ n21146;
  assign n21729 = n21728 ^ n21652;
  assign n21730 = n20334 ^ n20028;
  assign n21731 = n21730 ^ n21120;
  assign n21732 = n21731 ^ n21652;
  assign n21733 = n21729 & n21732;
  assign n21734 = n21733 ^ n21731;
  assign n21735 = n21734 ^ n21692;
  assign n21736 = n21693 & ~n21735;
  assign n21737 = n21736 ^ n21691;
  assign n21738 = n21737 ^ n21646;
  assign n21739 = ~n21689 & n21738;
  assign n21740 = n21739 ^ n21688;
  assign n21742 = n21741 ^ n21740;
  assign n21743 = n20698 ^ n20084;
  assign n21744 = n21743 ^ n21292;
  assign n21745 = n21744 ^ n21741;
  assign n21746 = n21742 & ~n21745;
  assign n21747 = n21746 ^ n21744;
  assign n21805 = n21748 ^ n21747;
  assign n21806 = ~n21751 & n21805;
  assign n21807 = n21806 ^ n21750;
  assign n21908 = n21808 ^ n21807;
  assign n21909 = n21811 & ~n21908;
  assign n21910 = n21909 ^ n21810;
  assign n21912 = n21911 ^ n21910;
  assign n21906 = n20126 ^ n19513;
  assign n21907 = n21906 ^ n21383;
  assign n21928 = n21911 ^ n21907;
  assign n21929 = n21912 & ~n21928;
  assign n21930 = n21929 ^ n21907;
  assign n21932 = n21931 ^ n21930;
  assign n21926 = n20130 ^ n19502;
  assign n21927 = n21926 ^ n20715;
  assign n21933 = n21932 ^ n21927;
  assign n21934 = n21933 ^ n18840;
  assign n21913 = n21912 ^ n21907;
  assign n21914 = n21913 ^ n18808;
  assign n21812 = n21811 ^ n21807;
  assign n21813 = n21812 ^ n18782;
  assign n21752 = n21751 ^ n21747;
  assign n21753 = n21752 ^ n19493;
  assign n21754 = n21744 ^ n21742;
  assign n21755 = n21754 ^ n19466;
  assign n21756 = n21737 ^ n21689;
  assign n21757 = n21756 ^ n19236;
  assign n21758 = n21734 ^ n21693;
  assign n21759 = n21758 ^ n19100;
  assign n21760 = n21731 ^ n21729;
  assign n21761 = n21760 ^ n19093;
  assign n21762 = n21725 ^ n21697;
  assign n21763 = n21762 ^ n19086;
  assign n21764 = n21722 ^ n21720;
  assign n21765 = n21764 ^ n18911;
  assign n21766 = n21716 ^ n21700;
  assign n21767 = n21766 ^ n18916;
  assign n21768 = n21713 ^ n21704;
  assign n21769 = n21768 ^ n18918;
  assign n21770 = n21710 ^ n21708;
  assign n21771 = n21770 ^ n18919;
  assign n21635 = n21634 ^ n21630;
  assign n21636 = n21635 ^ n18923;
  assign n21532 = n21531 ^ n21526;
  assign n21533 = n21532 ^ n19061;
  assign n21495 = n21494 ^ n21490;
  assign n21496 = n21495 ^ n18927;
  assign n21431 = n21430 ^ n20331;
  assign n21432 = n21431 ^ n19051;
  assign n21433 = n21426 ^ n20854;
  assign n21434 = n21433 ^ n18932;
  assign n21435 = n21423 ^ n21421;
  assign n21436 = n21435 ^ n18936;
  assign n21437 = n21416 ^ n21414;
  assign n21438 = n21437 ^ n18940;
  assign n21473 = n21472 ^ n21439;
  assign n21474 = ~n21440 & ~n21473;
  assign n21475 = n21474 ^ n18410;
  assign n21476 = n21475 ^ n21437;
  assign n21477 = ~n21438 & n21476;
  assign n21478 = n21477 ^ n18940;
  assign n21479 = n21478 ^ n21435;
  assign n21480 = n21436 & ~n21479;
  assign n21481 = n21480 ^ n18936;
  assign n21482 = n21481 ^ n21433;
  assign n21483 = ~n21434 & ~n21482;
  assign n21484 = n21483 ^ n18932;
  assign n21485 = n21484 ^ n21431;
  assign n21486 = ~n21432 & n21485;
  assign n21487 = n21486 ^ n19051;
  assign n21522 = n21495 ^ n21487;
  assign n21523 = ~n21496 & ~n21522;
  assign n21524 = n21523 ^ n18927;
  assign n21625 = n21532 ^ n21524;
  assign n21626 = ~n21533 & ~n21625;
  assign n21627 = n21626 ^ n19061;
  assign n21772 = n21635 ^ n21627;
  assign n21773 = n21636 & ~n21772;
  assign n21774 = n21773 ^ n18923;
  assign n21775 = n21774 ^ n21770;
  assign n21776 = n21771 & ~n21775;
  assign n21777 = n21776 ^ n18919;
  assign n21778 = n21777 ^ n21768;
  assign n21779 = ~n21769 & n21778;
  assign n21780 = n21779 ^ n18918;
  assign n21781 = n21780 ^ n21766;
  assign n21782 = ~n21767 & n21781;
  assign n21783 = n21782 ^ n18916;
  assign n21784 = n21783 ^ n21764;
  assign n21785 = n21765 & ~n21784;
  assign n21786 = n21785 ^ n18911;
  assign n21787 = n21786 ^ n21762;
  assign n21788 = n21763 & ~n21787;
  assign n21789 = n21788 ^ n19086;
  assign n21790 = n21789 ^ n21760;
  assign n21791 = ~n21761 & ~n21790;
  assign n21792 = n21791 ^ n19093;
  assign n21793 = n21792 ^ n21758;
  assign n21794 = ~n21759 & ~n21793;
  assign n21795 = n21794 ^ n19100;
  assign n21796 = n21795 ^ n21756;
  assign n21797 = ~n21757 & ~n21796;
  assign n21798 = n21797 ^ n19236;
  assign n21799 = n21798 ^ n21754;
  assign n21800 = n21755 & n21799;
  assign n21801 = n21800 ^ n19466;
  assign n21802 = n21801 ^ n21752;
  assign n21803 = ~n21753 & ~n21802;
  assign n21804 = n21803 ^ n19493;
  assign n21903 = n21812 ^ n21804;
  assign n21904 = n21813 & ~n21903;
  assign n21905 = n21904 ^ n18782;
  assign n21923 = n21913 ^ n21905;
  assign n21924 = ~n21914 & n21923;
  assign n21925 = n21924 ^ n18808;
  assign n21935 = n21934 ^ n21925;
  assign n21915 = n21914 ^ n21905;
  assign n21814 = n21813 ^ n21804;
  assign n21815 = n21801 ^ n21753;
  assign n21816 = n21792 ^ n21759;
  assign n21817 = n21789 ^ n21761;
  assign n21818 = n21786 ^ n21763;
  assign n21819 = n21783 ^ n21765;
  assign n21820 = n21777 ^ n21769;
  assign n21821 = n21774 ^ n21771;
  assign n21637 = n21636 ^ n21627;
  assign n21497 = n21496 ^ n21487;
  assign n21498 = n21484 ^ n21432;
  assign n21499 = n21481 ^ n21434;
  assign n21514 = ~n21512 & ~n21513;
  assign n21515 = n21475 ^ n21438;
  assign n21516 = n21514 & n21515;
  assign n21517 = n21478 ^ n21436;
  assign n21518 = n21516 & ~n21517;
  assign n21519 = ~n21499 & ~n21518;
  assign n21520 = ~n21498 & ~n21519;
  assign n21521 = n21497 & ~n21520;
  assign n21534 = n21533 ^ n21524;
  assign n21638 = ~n21521 & n21534;
  assign n21822 = n21637 & n21638;
  assign n21823 = n21821 & n21822;
  assign n21824 = ~n21820 & n21823;
  assign n21825 = n21780 ^ n21767;
  assign n21826 = ~n21824 & n21825;
  assign n21827 = ~n21819 & n21826;
  assign n21828 = n21818 & ~n21827;
  assign n21829 = ~n21817 & n21828;
  assign n21830 = ~n21816 & ~n21829;
  assign n21831 = n21795 ^ n21757;
  assign n21832 = ~n21830 & ~n21831;
  assign n21833 = n21798 ^ n21755;
  assign n21834 = n21832 & ~n21833;
  assign n21835 = n21815 & ~n21834;
  assign n21916 = ~n21814 & ~n21835;
  assign n21922 = n21915 & n21916;
  assign n21936 = n21935 ^ n21922;
  assign n21937 = n21936 ^ n2336;
  assign n21917 = n21916 ^ n21915;
  assign n21836 = n21835 ^ n21814;
  assign n1342 = n1323 ^ n1236;
  assign n1343 = n1342 ^ n1196;
  assign n1344 = n1343 ^ x487;
  assign n21837 = n21836 ^ n1344;
  assign n21838 = n21834 ^ n21815;
  assign n21839 = n21838 ^ n1186;
  assign n21892 = n21833 ^ n21832;
  assign n21840 = n21831 ^ n21830;
  assign n21841 = n21840 ^ n1165;
  assign n21884 = n21829 ^ n21816;
  assign n21842 = n21828 ^ n21817;
  assign n21846 = n21845 ^ n21842;
  assign n21876 = n21827 ^ n21818;
  assign n21847 = n21826 ^ n21819;
  assign n677 = n661 ^ n553;
  assign n678 = n677 ^ n674;
  assign n679 = n678 ^ x494;
  assign n21848 = n21847 ^ n679;
  assign n21849 = n21825 ^ n21824;
  assign n665 = n652 ^ n547;
  assign n669 = n668 ^ n665;
  assign n670 = n669 ^ x495;
  assign n21850 = n21849 ^ n670;
  assign n21851 = n21823 ^ n21820;
  assign n21855 = n21854 ^ n21851;
  assign n21856 = n21822 ^ n21821;
  assign n21860 = n21859 ^ n21856;
  assign n21639 = n21638 ^ n21637;
  assign n21535 = n21534 ^ n21521;
  assign n21539 = n21538 ^ n21535;
  assign n21540 = n21520 ^ n21497;
  assign n21544 = n21543 ^ n21540;
  assign n21545 = n21519 ^ n21498;
  assign n21549 = n21548 ^ n21545;
  assign n21611 = n21518 ^ n21499;
  assign n21603 = n21517 ^ n21516;
  assign n21598 = n21515 ^ n21514;
  assign n21595 = n21594 ^ n21550;
  assign n21596 = ~n21551 & n21595;
  assign n21597 = n21596 ^ n1774;
  assign n21599 = n21598 ^ n21597;
  assign n21600 = n21598 ^ n1908;
  assign n21601 = n21599 & ~n21600;
  assign n21602 = n21601 ^ n1908;
  assign n21604 = n21603 ^ n21602;
  assign n21608 = n21607 ^ n21603;
  assign n21609 = ~n21604 & n21608;
  assign n21610 = n21609 ^ n21607;
  assign n21612 = n21611 ^ n21610;
  assign n21613 = n21611 ^ n2078;
  assign n21614 = ~n21612 & n21613;
  assign n21615 = n21614 ^ n2078;
  assign n21616 = n21615 ^ n21545;
  assign n21617 = ~n21549 & n21616;
  assign n21618 = n21617 ^ n21548;
  assign n21619 = n21618 ^ n21540;
  assign n21620 = ~n21544 & n21619;
  assign n21621 = n21620 ^ n21543;
  assign n21622 = n21621 ^ n21535;
  assign n21623 = n21539 & ~n21622;
  assign n21624 = n21623 ^ n21538;
  assign n21640 = n21639 ^ n21624;
  assign n21861 = n21643 ^ n21639;
  assign n21862 = n21640 & ~n21861;
  assign n21863 = n21862 ^ n21643;
  assign n21864 = n21863 ^ n21856;
  assign n21865 = ~n21860 & n21864;
  assign n21866 = n21865 ^ n21859;
  assign n21867 = n21866 ^ n21851;
  assign n21868 = n21855 & ~n21867;
  assign n21869 = n21868 ^ n21854;
  assign n21870 = n21869 ^ n21849;
  assign n21871 = ~n21850 & n21870;
  assign n21872 = n21871 ^ n670;
  assign n21873 = n21872 ^ n21847;
  assign n21874 = ~n21848 & n21873;
  assign n21875 = n21874 ^ n679;
  assign n21877 = n21876 ^ n21875;
  assign n21878 = n21876 ^ n720;
  assign n21879 = ~n21877 & n21878;
  assign n21880 = n21879 ^ n720;
  assign n21881 = n21880 ^ n21842;
  assign n21882 = n21846 & ~n21881;
  assign n21883 = n21882 ^ n21845;
  assign n21885 = n21884 ^ n21883;
  assign n21886 = n21884 ^ n818;
  assign n21887 = ~n21885 & n21886;
  assign n21888 = n21887 ^ n818;
  assign n21889 = n21888 ^ n21840;
  assign n21890 = ~n21841 & n21889;
  assign n21891 = n21890 ^ n1165;
  assign n21893 = n21892 ^ n21891;
  assign n21894 = n21892 ^ n1171;
  assign n21895 = ~n21893 & n21894;
  assign n21896 = n21895 ^ n1171;
  assign n21897 = n21896 ^ n21838;
  assign n21898 = ~n21839 & n21897;
  assign n21899 = n21898 ^ n1186;
  assign n21900 = n21899 ^ n21836;
  assign n21901 = ~n21837 & n21900;
  assign n21902 = n21901 ^ n1344;
  assign n21918 = n21917 ^ n21902;
  assign n1357 = n1335 ^ n1251;
  assign n1358 = n1357 ^ n1351;
  assign n1359 = n1358 ^ x486;
  assign n21919 = n21917 ^ n1359;
  assign n21920 = n21918 & ~n21919;
  assign n21921 = n21920 ^ n1359;
  assign n21938 = n21937 ^ n21921;
  assign n21685 = n20889 ^ n20157;
  assign n21686 = n21685 ^ n21395;
  assign n22150 = n21938 ^ n21686;
  assign n22237 = n22150 ^ n19540;
  assign n22390 = n2652 ^ n1463;
  assign n22391 = n22390 ^ n2627;
  assign n22392 = n22391 ^ n1487;
  assign n22393 = ~n22237 & n22392;
  assign n22394 = n22393 ^ n1526;
  assign n21957 = n21922 & ~n21935;
  assign n21950 = n21931 ^ n21927;
  assign n21951 = ~n21932 & ~n21950;
  assign n21952 = n21951 ^ n21927;
  assign n21949 = n21231 ^ n1051;
  assign n21953 = n21952 ^ n21949;
  assign n21947 = n20137 ^ n19520;
  assign n21948 = n21947 ^ n20718;
  assign n21954 = n21953 ^ n21948;
  assign n21955 = n21954 ^ n18891;
  assign n21944 = n21933 ^ n21925;
  assign n21945 = n21934 & n21944;
  assign n21946 = n21945 ^ n18840;
  assign n21956 = n21955 ^ n21946;
  assign n21958 = n21957 ^ n21956;
  assign n21941 = n21936 ^ n21921;
  assign n21942 = n21937 & ~n21941;
  assign n21943 = n21942 ^ n2336;
  assign n21959 = n21958 ^ n21943;
  assign n2415 = n2414 ^ n2348;
  assign n2416 = n2415 ^ n2343;
  assign n2417 = n2416 ^ x484;
  assign n21960 = n21959 ^ n2417;
  assign n21939 = n21686 & n21938;
  assign n21683 = n20882 ^ n20164;
  assign n21684 = n21683 ^ n20857;
  assign n21940 = n21939 ^ n21684;
  assign n22153 = n21960 ^ n21940;
  assign n22151 = n19540 & n22150;
  assign n22152 = n22151 ^ n18898;
  assign n22238 = n22153 ^ n22152;
  assign n22395 = n22238 ^ n22237;
  assign n22396 = n22395 ^ n1526;
  assign n22397 = n22394 & ~n22396;
  assign n22398 = n22397 ^ n22393;
  assign n22239 = n22237 & n22238;
  assign n22154 = n22153 ^ n22151;
  assign n22155 = n22152 & ~n22154;
  assign n22156 = n22155 ^ n18898;
  assign n21985 = n20899 ^ n20215;
  assign n21986 = n21985 ^ n20856;
  assign n21974 = n21949 ^ n21948;
  assign n21975 = ~n21953 & ~n21974;
  assign n21976 = n21975 ^ n21948;
  assign n21973 = n21234 ^ n21128;
  assign n21977 = n21976 ^ n21973;
  assign n21971 = n20115 ^ n19498;
  assign n21972 = n21971 ^ n20722;
  assign n21978 = n21977 ^ n21972;
  assign n21979 = n21978 ^ n18992;
  assign n21968 = n21954 ^ n21946;
  assign n21969 = ~n21955 & n21968;
  assign n21970 = n21969 ^ n18891;
  assign n21980 = n21979 ^ n21970;
  assign n21967 = n21956 & ~n21957;
  assign n21981 = n21980 ^ n21967;
  assign n21982 = n21981 ^ n2411;
  assign n21964 = n21958 ^ n2417;
  assign n21965 = n21959 & ~n21964;
  assign n21966 = n21965 ^ n2417;
  assign n21983 = n21982 ^ n21966;
  assign n21961 = n21960 ^ n21684;
  assign n21962 = ~n21940 & ~n21961;
  assign n21963 = n21962 ^ n21939;
  assign n21984 = n21983 ^ n21963;
  assign n22148 = n21986 ^ n21984;
  assign n22149 = n22148 ^ n19550;
  assign n22236 = n22156 ^ n22149;
  assign n22385 = n22239 ^ n22236;
  assign n22389 = n22388 ^ n22385;
  assign n22598 = n22398 ^ n22389;
  assign n22601 = n22600 ^ n22598;
  assign n22603 = n21527 ^ n20927;
  assign n22067 = n21591 ^ n21553;
  assign n22604 = n22603 ^ n22067;
  assign n22602 = n22395 ^ n22394;
  assign n22605 = n22604 ^ n22602;
  assign n22607 = n21491 ^ n20920;
  assign n21668 = n21588 ^ n1676;
  assign n22608 = n22607 ^ n21668;
  assign n22606 = n22392 ^ n22237;
  assign n22609 = n22608 ^ n22606;
  assign n22686 = n20913 ^ n20849;
  assign n22057 = n21583 ^ n21555;
  assign n22687 = n22686 ^ n22057;
  assign n22678 = n20839 ^ n19755;
  assign n22679 = n22678 ^ n21388;
  assign n22646 = n20818 ^ n20147;
  assign n22647 = n22646 ^ n21358;
  assign n22645 = n21899 ^ n21837;
  assign n22648 = n22647 ^ n22645;
  assign n22615 = n20707 ^ n20137;
  assign n22616 = n22615 ^ n21303;
  assign n22614 = n21893 ^ n1171;
  assign n22617 = n22616 ^ n22614;
  assign n22519 = n20722 ^ n20130;
  assign n22520 = n22519 ^ n21279;
  assign n22518 = n21888 ^ n21841;
  assign n22521 = n22520 ^ n22518;
  assign n22338 = n20718 ^ n20126;
  assign n22026 = n21256 ^ n2273;
  assign n22339 = n22338 ^ n22026;
  assign n22337 = n21885 ^ n818;
  assign n22340 = n22339 ^ n22337;
  assign n22324 = n20715 ^ n20121;
  assign n22001 = n21237 ^ n21126;
  assign n22325 = n22324 ^ n22001;
  assign n22323 = n21880 ^ n21846;
  assign n22326 = n22325 ^ n22323;
  assign n22310 = n21383 ^ n20767;
  assign n22311 = n22310 ^ n21973;
  assign n22309 = n21877 ^ n720;
  assign n22312 = n22311 ^ n22309;
  assign n22295 = n21346 ^ n20698;
  assign n22296 = n22295 ^ n21949;
  assign n22294 = n21872 ^ n21848;
  assign n22297 = n22296 ^ n22294;
  assign n22225 = n21866 ^ n21855;
  assign n22114 = n21268 ^ n20334;
  assign n22115 = n22114 ^ n21808;
  assign n22113 = n21863 ^ n21860;
  assign n22116 = n22115 ^ n22113;
  assign n22100 = n21621 ^ n21539;
  assign n21648 = n21618 ^ n21544;
  assign n21645 = n21070 ^ n20340;
  assign n21647 = n21646 ^ n21645;
  assign n21649 = n21648 ^ n21647;
  assign n22090 = n21615 ^ n21549;
  assign n21651 = n20862 ^ n20344;
  assign n21653 = n21652 ^ n21651;
  assign n21650 = n21612 ^ n2078;
  assign n21654 = n21653 ^ n21650;
  assign n22080 = n21607 ^ n21604;
  assign n21658 = n21599 ^ n1908;
  assign n21655 = n20962 ^ n20410;
  assign n21657 = n21656 ^ n21655;
  assign n21659 = n21658 ^ n21657;
  assign n21660 = n20870 ^ n20354;
  assign n21662 = n21661 ^ n21660;
  assign n21664 = n21663 ^ n21662;
  assign n21665 = n20877 ^ n20358;
  assign n21667 = n21666 ^ n21665;
  assign n21669 = n21668 ^ n21667;
  assign n21671 = n20852 ^ n20388;
  assign n21672 = n21671 ^ n21527;
  assign n21670 = n21580 ^ n21560;
  assign n21673 = n21672 ^ n21670;
  assign n21676 = n20927 ^ n20378;
  assign n21677 = n21676 ^ n20849;
  assign n21675 = n21574 ^ n21573;
  assign n21678 = n21677 ^ n21675;
  assign n21680 = n20920 ^ n20850;
  assign n21681 = n21680 ^ n20370;
  assign n21679 = n21568 ^ n21504;
  assign n21682 = n21681 ^ n21679;
  assign n22029 = n21380 ^ n19755;
  assign n22030 = n22029 ^ n20772;
  assign n21996 = ~n21967 & ~n21980;
  assign n22006 = n20147 ^ n18905;
  assign n22007 = n22006 ^ n20707;
  assign n22002 = n21973 ^ n21972;
  assign n22003 = n21977 & n22002;
  assign n22004 = n22003 ^ n21972;
  assign n22005 = n22004 ^ n22001;
  assign n22008 = n22007 ^ n22005;
  assign n21997 = n21978 ^ n21970;
  assign n21998 = ~n21979 & n21997;
  assign n21999 = n21998 ^ n18992;
  assign n22000 = n21999 ^ n18999;
  assign n22009 = n22008 ^ n22000;
  assign n22027 = n21996 & n22009;
  assign n22028 = n22027 ^ n22026;
  assign n22031 = n22030 ^ n22028;
  assign n1548 = n1547 ^ n1424;
  assign n1549 = n1548 ^ n1517;
  assign n1550 = n1549 ^ x481;
  assign n22032 = n22031 ^ n1550;
  assign n22010 = n22009 ^ n21996;
  assign n21993 = n21981 ^ n21966;
  assign n21994 = ~n21982 & n21993;
  assign n21995 = n21994 ^ n2411;
  assign n22011 = n22010 ^ n21995;
  assign n2563 = n2559 ^ n2486;
  assign n2567 = n2566 ^ n2563;
  assign n2568 = n2567 ^ x482;
  assign n22023 = n22010 ^ n2568;
  assign n22024 = n22011 & ~n22023;
  assign n22025 = n22024 ^ n2568;
  assign n22033 = n22032 ^ n22025;
  assign n22019 = n22008 ^ n18999;
  assign n22020 = n22008 ^ n21999;
  assign n22021 = n22019 & n22020;
  assign n22022 = n22021 ^ n18999;
  assign n22034 = n22033 ^ n22022;
  assign n22016 = n22007 ^ n22001;
  assign n22017 = n22005 & ~n22016;
  assign n22018 = n22017 ^ n22007;
  assign n22035 = n22034 ^ n22018;
  assign n21990 = n20906 ^ n20300;
  assign n21991 = n21990 ^ n20855;
  assign n21987 = n21986 ^ n21983;
  assign n21988 = n21984 & n21987;
  assign n21989 = n21988 ^ n21986;
  assign n21992 = n21991 ^ n21989;
  assign n22012 = n22011 ^ n2568;
  assign n22013 = n22012 ^ n21989;
  assign n22014 = ~n21992 & ~n22013;
  assign n22015 = n22014 ^ n21991;
  assign n22036 = n22035 ^ n22015;
  assign n22037 = n20913 ^ n20320;
  assign n22038 = n22037 ^ n21420;
  assign n22039 = n22038 ^ n22035;
  assign n22040 = ~n22036 & ~n22039;
  assign n22041 = n22040 ^ n22038;
  assign n22042 = n22041 ^ n21679;
  assign n22043 = ~n21682 & n22042;
  assign n22044 = n22043 ^ n21681;
  assign n22045 = n22044 ^ n21675;
  assign n22046 = ~n21678 & n22045;
  assign n22047 = n22046 ^ n21677;
  assign n21674 = n21577 ^ n21565;
  assign n22048 = n22047 ^ n21674;
  assign n22049 = n20934 ^ n20364;
  assign n22050 = n22049 ^ n21491;
  assign n22051 = n22050 ^ n21674;
  assign n22052 = ~n22048 & ~n22051;
  assign n22053 = n22052 ^ n22050;
  assign n22054 = n22053 ^ n21670;
  assign n22055 = ~n21673 & n22054;
  assign n22056 = n22055 ^ n21672;
  assign n22058 = n22057 ^ n22056;
  assign n22059 = n21631 ^ n20330;
  assign n22060 = n22059 ^ n20362;
  assign n22061 = n22060 ^ n22057;
  assign n22062 = n22058 & ~n22061;
  assign n22063 = n22062 ^ n22060;
  assign n22064 = n22063 ^ n21668;
  assign n22065 = n21669 & ~n22064;
  assign n22066 = n22065 ^ n21667;
  assign n22068 = n22067 ^ n22066;
  assign n22069 = n20874 ^ n19749;
  assign n22070 = n22069 ^ n21701;
  assign n22071 = n22070 ^ n22067;
  assign n22072 = ~n22068 & ~n22071;
  assign n22073 = n22072 ^ n22070;
  assign n22074 = n22073 ^ n21662;
  assign n22075 = ~n21664 & n22074;
  assign n22076 = n22075 ^ n21663;
  assign n22077 = n22076 ^ n21658;
  assign n22078 = n21659 & ~n22077;
  assign n22079 = n22078 ^ n21657;
  assign n22081 = n22080 ^ n22079;
  assign n22082 = n20866 ^ n20348;
  assign n22083 = n22082 ^ n21694;
  assign n22084 = n22083 ^ n22080;
  assign n22085 = n22081 & ~n22084;
  assign n22086 = n22085 ^ n22083;
  assign n22087 = n22086 ^ n21650;
  assign n22088 = n21654 & n22087;
  assign n22089 = n22088 ^ n21653;
  assign n22091 = n22090 ^ n22089;
  assign n22092 = n20975 ^ n20423;
  assign n22093 = n22092 ^ n21692;
  assign n22094 = n22093 ^ n22090;
  assign n22095 = n22091 & ~n22094;
  assign n22096 = n22095 ^ n22093;
  assign n22097 = n22096 ^ n21647;
  assign n22098 = n21649 & n22097;
  assign n22099 = n22098 ^ n21648;
  assign n22101 = n22100 ^ n22099;
  assign n22102 = n21120 ^ n20338;
  assign n22103 = n22102 ^ n21741;
  assign n22104 = n22103 ^ n22100;
  assign n22105 = n22101 & n22104;
  assign n22106 = n22105 ^ n22103;
  assign n21644 = n21643 ^ n21640;
  assign n22107 = n22106 ^ n21644;
  assign n22108 = n21249 ^ n20335;
  assign n22109 = n22108 ^ n21748;
  assign n22110 = n22109 ^ n21644;
  assign n22111 = n22107 & n22110;
  assign n22112 = n22111 ^ n22109;
  assign n22222 = n22113 ^ n22112;
  assign n22223 = n22116 & ~n22222;
  assign n22224 = n22223 ^ n22115;
  assign n22226 = n22225 ^ n22224;
  assign n22220 = n21292 ^ n20448;
  assign n22221 = n22220 ^ n21911;
  assign n22280 = n22225 ^ n22221;
  assign n22281 = n22226 & n22280;
  assign n22282 = n22281 ^ n22221;
  assign n22279 = n21869 ^ n21850;
  assign n22283 = n22282 ^ n22279;
  assign n22277 = n21318 ^ n20540;
  assign n22278 = n22277 ^ n21931;
  assign n22291 = n22279 ^ n22278;
  assign n22292 = n22283 & n22291;
  assign n22293 = n22292 ^ n22278;
  assign n22306 = n22296 ^ n22293;
  assign n22307 = ~n22297 & n22306;
  assign n22308 = n22307 ^ n22294;
  assign n22320 = n22309 ^ n22308;
  assign n22321 = ~n22312 & n22320;
  assign n22322 = n22321 ^ n22311;
  assign n22334 = n22323 ^ n22322;
  assign n22335 = n22326 & n22334;
  assign n22336 = n22335 ^ n22325;
  assign n22515 = n22337 ^ n22336;
  assign n22516 = n22340 & ~n22515;
  assign n22517 = n22516 ^ n22339;
  assign n22618 = n22520 ^ n22517;
  assign n22619 = n22521 & n22618;
  assign n22620 = n22619 ^ n22518;
  assign n22631 = n22620 ^ n22614;
  assign n22632 = n22617 & n22631;
  assign n22633 = n22632 ^ n22616;
  assign n22551 = n21896 ^ n21839;
  assign n22634 = n22633 ^ n22551;
  assign n22629 = n20772 ^ n20115;
  assign n22630 = n22629 ^ n21329;
  assign n22642 = n22630 ^ n22551;
  assign n22643 = n22634 & n22642;
  assign n22644 = n22643 ^ n22630;
  assign n22675 = n22645 ^ n22644;
  assign n22676 = ~n22648 & ~n22675;
  assign n22677 = n22676 ^ n22647;
  assign n22680 = n22679 ^ n22677;
  assign n22544 = n21918 ^ n1359;
  assign n22681 = n22680 ^ n22544;
  assign n22649 = n22648 ^ n22644;
  assign n22650 = n22649 ^ n18905;
  assign n22635 = n22634 ^ n22630;
  assign n22636 = n22635 ^ n19498;
  assign n22621 = n22620 ^ n22617;
  assign n22522 = n22521 ^ n22517;
  assign n22610 = n22522 ^ n19502;
  assign n22341 = n22340 ^ n22336;
  assign n22342 = n22341 ^ n19513;
  assign n22327 = n22326 ^ n22322;
  assign n22328 = n22327 ^ n19508;
  assign n22313 = n22312 ^ n22308;
  assign n22316 = n22313 ^ n20104;
  assign n22298 = n22297 ^ n22293;
  assign n22299 = n22298 ^ n20084;
  assign n22284 = n22283 ^ n22278;
  assign n22287 = n22284 ^ n20066;
  assign n22227 = n22226 ^ n22221;
  assign n22117 = n22116 ^ n22112;
  assign n22118 = n22117 ^ n20028;
  assign n22119 = n22109 ^ n22107;
  assign n22120 = n22119 ^ n20008;
  assign n22121 = n22103 ^ n22101;
  assign n22122 = n22121 ^ n19923;
  assign n22206 = n22096 ^ n21649;
  assign n22123 = n22093 ^ n22091;
  assign n22124 = n22123 ^ n19759;
  assign n22125 = n22086 ^ n21654;
  assign n22126 = n22125 ^ n19760;
  assign n22127 = n22083 ^ n22081;
  assign n22128 = n22127 ^ n19764;
  assign n22192 = n22076 ^ n21659;
  assign n22129 = n22070 ^ n22068;
  assign n22130 = n22129 ^ n19751;
  assign n22131 = n22063 ^ n21669;
  assign n22132 = n22131 ^ n19774;
  assign n22133 = n22060 ^ n22058;
  assign n22134 = n22133 ^ n19796;
  assign n22135 = n22053 ^ n21673;
  assign n22136 = n22135 ^ n19778;
  assign n22137 = n22050 ^ n22048;
  assign n22138 = n22137 ^ n19780;
  assign n22139 = n22044 ^ n21678;
  assign n22140 = n22139 ^ n19738;
  assign n22141 = n22041 ^ n21682;
  assign n22142 = n22141 ^ n19651;
  assign n22143 = n22038 ^ n22036;
  assign n22144 = n22143 ^ n19637;
  assign n22145 = n22012 ^ n21991;
  assign n22146 = n22145 ^ n21989;
  assign n22147 = n22146 ^ n19604;
  assign n22157 = n22156 ^ n22148;
  assign n22158 = n22149 & ~n22157;
  assign n22159 = n22158 ^ n19550;
  assign n22160 = n22159 ^ n22146;
  assign n22161 = n22147 & ~n22160;
  assign n22162 = n22161 ^ n19604;
  assign n22163 = n22162 ^ n22143;
  assign n22164 = ~n22144 & n22163;
  assign n22165 = n22164 ^ n19637;
  assign n22166 = n22165 ^ n22141;
  assign n22167 = ~n22142 & ~n22166;
  assign n22168 = n22167 ^ n19651;
  assign n22169 = n22168 ^ n22139;
  assign n22170 = ~n22140 & n22169;
  assign n22171 = n22170 ^ n19738;
  assign n22172 = n22171 ^ n22137;
  assign n22173 = ~n22138 & n22172;
  assign n22174 = n22173 ^ n19780;
  assign n22175 = n22174 ^ n22135;
  assign n22176 = n22136 & ~n22175;
  assign n22177 = n22176 ^ n19778;
  assign n22178 = n22177 ^ n22133;
  assign n22179 = ~n22134 & ~n22178;
  assign n22180 = n22179 ^ n19796;
  assign n22181 = n22180 ^ n22131;
  assign n22182 = ~n22132 & ~n22181;
  assign n22183 = n22182 ^ n19774;
  assign n22184 = n22183 ^ n22129;
  assign n22185 = n22130 & ~n22184;
  assign n22186 = n22185 ^ n19751;
  assign n22187 = n22186 ^ n19770;
  assign n22188 = n22073 ^ n21664;
  assign n22189 = n22188 ^ n22186;
  assign n22190 = ~n22187 & n22189;
  assign n22191 = n22190 ^ n19770;
  assign n22193 = n22192 ^ n22191;
  assign n22194 = n22192 ^ n19768;
  assign n22195 = n22193 & n22194;
  assign n22196 = n22195 ^ n19768;
  assign n22197 = n22196 ^ n22127;
  assign n22198 = n22128 & n22197;
  assign n22199 = n22198 ^ n19764;
  assign n22200 = n22199 ^ n22125;
  assign n22201 = n22126 & n22200;
  assign n22202 = n22201 ^ n19760;
  assign n22203 = n22202 ^ n22123;
  assign n22204 = ~n22124 & ~n22203;
  assign n22205 = n22204 ^ n19759;
  assign n22207 = n22206 ^ n22205;
  assign n22208 = n22206 ^ n19883;
  assign n22209 = ~n22207 & n22208;
  assign n22210 = n22209 ^ n19883;
  assign n22211 = n22210 ^ n22121;
  assign n22212 = n22122 & n22211;
  assign n22213 = n22212 ^ n19923;
  assign n22214 = n22213 ^ n22119;
  assign n22215 = ~n22120 & n22214;
  assign n22216 = n22215 ^ n20008;
  assign n22217 = n22216 ^ n22117;
  assign n22218 = ~n22118 & ~n22217;
  assign n22219 = n22218 ^ n20028;
  assign n22228 = n22227 ^ n22219;
  assign n22273 = n22227 ^ n20047;
  assign n22274 = n22228 & ~n22273;
  assign n22275 = n22274 ^ n20047;
  assign n22288 = n22284 ^ n22275;
  assign n22289 = n22287 & ~n22288;
  assign n22290 = n22289 ^ n20066;
  assign n22302 = n22298 ^ n22290;
  assign n22303 = n22299 & ~n22302;
  assign n22304 = n22303 ^ n20084;
  assign n22317 = n22313 ^ n22304;
  assign n22318 = ~n22316 & ~n22317;
  assign n22319 = n22318 ^ n20104;
  assign n22331 = n22327 ^ n22319;
  assign n22332 = n22328 & ~n22331;
  assign n22333 = n22332 ^ n19508;
  assign n22511 = n22341 ^ n22333;
  assign n22512 = n22342 & n22511;
  assign n22513 = n22512 ^ n19513;
  assign n22611 = n22522 ^ n22513;
  assign n22612 = ~n22610 & ~n22611;
  assign n22613 = n22612 ^ n19502;
  assign n22622 = n22621 ^ n22613;
  assign n22626 = n22621 ^ n19520;
  assign n22627 = ~n22622 & n22626;
  assign n22628 = n22627 ^ n19520;
  assign n22639 = n22635 ^ n22628;
  assign n22640 = n22636 & n22639;
  assign n22641 = n22640 ^ n19498;
  assign n22671 = n22649 ^ n22641;
  assign n22672 = ~n22650 & ~n22671;
  assign n22673 = n22672 ^ n18905;
  assign n22674 = n22673 ^ n18903;
  assign n22682 = n22681 ^ n22674;
  assign n22623 = n22622 ^ n19520;
  assign n22514 = n22513 ^ n19502;
  assign n22523 = n22522 ^ n22514;
  assign n22229 = n22228 ^ n20047;
  assign n22230 = n22213 ^ n22120;
  assign n22231 = n22210 ^ n22122;
  assign n22232 = n22207 ^ n19883;
  assign n22233 = n22202 ^ n22124;
  assign n22234 = n22196 ^ n22128;
  assign n22235 = n22193 ^ n19768;
  assign n22240 = n22236 & n22239;
  assign n22241 = n22159 ^ n22147;
  assign n22242 = n22240 & n22241;
  assign n22243 = n22162 ^ n22144;
  assign n22244 = n22242 & ~n22243;
  assign n22245 = n22165 ^ n22142;
  assign n22246 = ~n22244 & n22245;
  assign n22247 = n22168 ^ n22140;
  assign n22248 = ~n22246 & n22247;
  assign n22249 = n22171 ^ n22138;
  assign n22250 = ~n22248 & ~n22249;
  assign n22251 = n22174 ^ n22136;
  assign n22252 = n22250 & n22251;
  assign n22253 = n22177 ^ n22134;
  assign n22254 = n22252 & ~n22253;
  assign n22255 = n22180 ^ n22132;
  assign n22256 = ~n22254 & ~n22255;
  assign n22257 = n22183 ^ n22130;
  assign n22258 = ~n22256 & n22257;
  assign n22259 = n22188 ^ n19770;
  assign n22260 = n22259 ^ n22186;
  assign n22261 = ~n22258 & ~n22260;
  assign n22262 = ~n22235 & ~n22261;
  assign n22263 = n22234 & n22262;
  assign n22264 = n22199 ^ n22126;
  assign n22265 = n22263 & ~n22264;
  assign n22266 = ~n22233 & n22265;
  assign n22267 = n22232 & ~n22266;
  assign n22268 = n22231 & n22267;
  assign n22269 = ~n22230 & ~n22268;
  assign n22270 = n22216 ^ n22118;
  assign n22271 = n22269 & ~n22270;
  assign n22272 = ~n22229 & ~n22271;
  assign n22276 = n22275 ^ n20066;
  assign n22285 = n22284 ^ n22276;
  assign n22286 = ~n22272 & ~n22285;
  assign n22300 = n22299 ^ n22290;
  assign n22301 = n22286 & ~n22300;
  assign n22305 = n22304 ^ n20104;
  assign n22314 = n22313 ^ n22305;
  assign n22315 = ~n22301 & ~n22314;
  assign n22329 = n22328 ^ n22319;
  assign n22330 = ~n22315 & n22329;
  assign n22343 = n22342 ^ n22333;
  assign n22524 = n22330 & n22343;
  assign n22624 = n22523 & n22524;
  assign n22625 = ~n22623 & ~n22624;
  assign n22637 = n22636 ^ n22628;
  assign n22638 = ~n22625 & n22637;
  assign n22651 = n22650 ^ n22641;
  assign n22670 = n22638 & n22651;
  assign n22683 = n22682 ^ n22670;
  assign n22652 = n22651 ^ n22638;
  assign n22653 = n22652 ^ n2539;
  assign n22654 = n22637 ^ n22625;
  assign n22655 = n22654 ^ n2523;
  assign n22659 = n22624 ^ n22623;
  assign n22526 = n2383 ^ n1406;
  assign n22527 = n22526 ^ n2276;
  assign n22528 = n22527 ^ n1535;
  assign n22525 = n22524 ^ n22523;
  assign n22529 = n22528 ^ n22525;
  assign n22345 = n2376 ^ n1388;
  assign n22346 = n22345 ^ n17431;
  assign n22347 = n22346 ^ n2267;
  assign n22344 = n22343 ^ n22330;
  assign n22348 = n22347 ^ n22344;
  assign n22349 = n22329 ^ n22315;
  assign n1203 = n1202 ^ n1115;
  assign n1210 = n1209 ^ n1203;
  assign n1214 = n1213 ^ n1210;
  assign n22350 = n22349 ^ n1214;
  assign n22351 = n22314 ^ n22301;
  assign n22355 = n22354 ^ n22351;
  assign n22356 = n22300 ^ n22286;
  assign n22357 = n22356 ^ n1038;
  assign n22358 = n22285 ^ n22272;
  assign n22359 = n22358 ^ n897;
  assign n22491 = n22271 ^ n22229;
  assign n22486 = n22270 ^ n22269;
  assign n22473 = n22267 ^ n22231;
  assign n22360 = n22266 ^ n22232;
  assign n22364 = n22363 ^ n22360;
  assign n22365 = n22265 ^ n22233;
  assign n22369 = n22368 ^ n22365;
  assign n22459 = n22264 ^ n22263;
  assign n22454 = n22262 ^ n22234;
  assign n22446 = n22261 ^ n22235;
  assign n22438 = n22260 ^ n22258;
  assign n22370 = n22255 ^ n22254;
  assign n22371 = n22370 ^ n2188;
  assign n22372 = n22253 ^ n22252;
  assign n22373 = n22372 ^ n2012;
  assign n22374 = n22251 ^ n22250;
  assign n22375 = n22374 ^ n1890;
  assign n22376 = n22249 ^ n22248;
  assign n22377 = n22376 ^ n1872;
  assign n22416 = n22247 ^ n22246;
  assign n22408 = n22245 ^ n22244;
  assign n22378 = n22243 ^ n22242;
  assign n22382 = n22381 ^ n22378;
  assign n22383 = n22241 ^ n22240;
  assign n22384 = n22383 ^ n1445;
  assign n22399 = n22398 ^ n22385;
  assign n22400 = n22389 & ~n22399;
  assign n22401 = n22400 ^ n22388;
  assign n22402 = n22401 ^ n22383;
  assign n22403 = n22384 & ~n22402;
  assign n22404 = n22403 ^ n1445;
  assign n22405 = n22404 ^ n22378;
  assign n22406 = ~n22382 & n22405;
  assign n22407 = n22406 ^ n22381;
  assign n22409 = n22408 ^ n22407;
  assign n22413 = n22412 ^ n22408;
  assign n22414 = ~n22409 & n22413;
  assign n22415 = n22414 ^ n22412;
  assign n22417 = n22416 ^ n22415;
  assign n22418 = n22416 ^ n1860;
  assign n22419 = n22417 & ~n22418;
  assign n22420 = n22419 ^ n1860;
  assign n22421 = n22420 ^ n22376;
  assign n22422 = ~n22377 & n22421;
  assign n22423 = n22422 ^ n1872;
  assign n22424 = n22423 ^ n22374;
  assign n22425 = ~n22375 & n22424;
  assign n22426 = n22425 ^ n1890;
  assign n22427 = n22426 ^ n22372;
  assign n22428 = n22373 & ~n22427;
  assign n22429 = n22428 ^ n2012;
  assign n22430 = n22429 ^ n22370;
  assign n22431 = n22371 & ~n22430;
  assign n22432 = n22431 ^ n2188;
  assign n22433 = n22432 ^ n2174;
  assign n22434 = n22257 ^ n22256;
  assign n22435 = n22434 ^ n22432;
  assign n22436 = n22433 & ~n22435;
  assign n22437 = n22436 ^ n2174;
  assign n22439 = n22438 ^ n22437;
  assign n22443 = n22442 ^ n22437;
  assign n22444 = ~n22439 & n22443;
  assign n22445 = n22444 ^ n22442;
  assign n22447 = n22446 ^ n22445;
  assign n22451 = n22450 ^ n22446;
  assign n22452 = n22447 & ~n22451;
  assign n22453 = n22452 ^ n22450;
  assign n22455 = n22454 ^ n22453;
  assign n22456 = n22454 ^ n605;
  assign n22457 = n22455 & ~n22456;
  assign n22458 = n22457 ^ n605;
  assign n22460 = n22459 ^ n22458;
  assign n22461 = n20632 ^ n13810;
  assign n22462 = n22461 ^ n17451;
  assign n22463 = n22462 ^ n522;
  assign n22464 = n22463 ^ n22459;
  assign n22465 = ~n22460 & n22464;
  assign n22466 = n22465 ^ n22463;
  assign n22467 = n22466 ^ n22365;
  assign n22468 = n22369 & ~n22467;
  assign n22469 = n22468 ^ n22368;
  assign n22470 = n22469 ^ n22360;
  assign n22471 = ~n22364 & n22470;
  assign n22472 = n22471 ^ n22363;
  assign n22474 = n22473 ^ n22472;
  assign n22478 = n22477 ^ n22472;
  assign n22479 = ~n22474 & n22478;
  assign n22480 = n22479 ^ n22477;
  assign n777 = n747 ^ n705;
  assign n784 = n783 ^ n777;
  assign n788 = n787 ^ n784;
  assign n22481 = n22480 ^ n788;
  assign n22482 = n22268 ^ n22230;
  assign n22483 = n22482 ^ n788;
  assign n22484 = n22481 & n22483;
  assign n22485 = n22484 ^ n22480;
  assign n22487 = n22486 ^ n22485;
  assign n22488 = n22486 ^ n800;
  assign n22489 = ~n22487 & n22488;
  assign n22490 = n22489 ^ n800;
  assign n22492 = n22491 ^ n22490;
  assign n22493 = n22491 ^ n882;
  assign n22494 = ~n22492 & n22493;
  assign n22495 = n22494 ^ n882;
  assign n22496 = n22495 ^ n22358;
  assign n22497 = ~n22359 & n22496;
  assign n22498 = n22497 ^ n897;
  assign n22499 = n22498 ^ n22356;
  assign n22500 = n22357 & ~n22499;
  assign n22501 = n22500 ^ n1038;
  assign n22502 = n22501 ^ n22354;
  assign n22503 = n22355 & ~n22502;
  assign n22504 = n22503 ^ n22351;
  assign n22505 = n22504 ^ n22349;
  assign n22506 = n22350 & ~n22505;
  assign n22507 = n22506 ^ n1214;
  assign n22508 = n22507 ^ n22344;
  assign n22509 = ~n22348 & n22508;
  assign n22510 = n22509 ^ n22347;
  assign n22656 = n22525 ^ n22510;
  assign n22657 = ~n22529 & n22656;
  assign n22658 = n22657 ^ n22528;
  assign n22660 = n22659 ^ n22658;
  assign n2509 = n2455 ^ n2395;
  assign n2510 = n2509 ^ n2508;
  assign n2511 = n2510 ^ n2360;
  assign n22661 = n22659 ^ n2511;
  assign n22662 = ~n22660 & n22661;
  assign n22663 = n22662 ^ n2511;
  assign n22664 = n22663 ^ n2523;
  assign n22665 = n22655 & ~n22664;
  assign n22666 = n22665 ^ n22654;
  assign n22667 = n22666 ^ n22652;
  assign n22668 = ~n22653 & n22667;
  assign n22669 = n22668 ^ n2539;
  assign n22684 = n22683 ^ n22669;
  assign n22685 = n22684 ^ n2634;
  assign n22688 = n22687 ^ n22685;
  assign n22691 = n22666 ^ n22653;
  assign n22689 = n20906 ^ n20850;
  assign n22690 = n22689 ^ n21670;
  assign n22692 = n22691 ^ n22690;
  assign n22694 = n21420 ^ n20899;
  assign n22695 = n22694 ^ n21674;
  assign n22693 = n22663 ^ n22655;
  assign n22696 = n22695 ^ n22693;
  assign n22530 = n22529 ^ n22510;
  assign n22531 = n20889 ^ n20856;
  assign n22532 = n22531 ^ n21679;
  assign n22699 = ~n22530 & n22532;
  assign n22697 = n20882 ^ n20855;
  assign n22698 = n22697 ^ n21675;
  assign n22700 = n22699 ^ n22698;
  assign n22701 = n22660 ^ n2511;
  assign n22702 = n22701 ^ n22698;
  assign n22703 = ~n22700 & n22702;
  assign n22704 = n22703 ^ n22699;
  assign n22705 = n22704 ^ n22693;
  assign n22706 = n22696 & ~n22705;
  assign n22707 = n22706 ^ n22695;
  assign n22708 = n22707 ^ n22690;
  assign n22709 = n22692 & n22708;
  assign n22710 = n22709 ^ n22691;
  assign n22711 = n22710 ^ n22685;
  assign n22712 = ~n22688 & ~n22711;
  assign n22713 = n22712 ^ n22687;
  assign n22714 = n22713 ^ n22606;
  assign n22715 = ~n22609 & n22714;
  assign n22716 = n22715 ^ n22608;
  assign n22717 = n22716 ^ n22602;
  assign n22718 = n22605 & ~n22717;
  assign n22719 = n22718 ^ n22604;
  assign n22720 = n22719 ^ n22598;
  assign n22721 = ~n22601 & ~n22720;
  assign n22722 = n22721 ^ n22600;
  assign n22595 = n21666 ^ n20852;
  assign n22596 = n22595 ^ n21658;
  assign n22540 = n22401 ^ n22384;
  assign n22597 = n22596 ^ n22540;
  assign n22844 = n22722 ^ n22597;
  assign n22845 = n22844 ^ n20388;
  assign n22880 = n22719 ^ n22601;
  assign n22846 = n22716 ^ n22604;
  assign n22847 = n22846 ^ n22602;
  assign n22848 = n22847 ^ n20378;
  assign n22849 = n22713 ^ n22609;
  assign n22850 = n22849 ^ n20370;
  assign n22851 = n22710 ^ n22687;
  assign n22852 = n22851 ^ n22685;
  assign n22853 = n22852 ^ n20320;
  assign n22533 = n22532 ^ n22530;
  assign n22854 = n20157 & ~n22533;
  assign n22855 = n22854 ^ n20164;
  assign n22856 = n22701 ^ n22700;
  assign n22857 = n22856 ^ n22854;
  assign n22858 = ~n22855 & n22857;
  assign n22859 = n22858 ^ n20164;
  assign n22860 = n22859 ^ n20215;
  assign n22861 = n22704 ^ n22695;
  assign n22862 = n22861 ^ n22693;
  assign n22863 = n22862 ^ n22859;
  assign n22864 = n22860 & n22863;
  assign n22865 = n22864 ^ n20215;
  assign n22866 = n22865 ^ n20300;
  assign n22867 = n22707 ^ n22692;
  assign n22868 = n22867 ^ n22865;
  assign n22869 = n22866 & n22868;
  assign n22870 = n22869 ^ n20300;
  assign n22871 = n22870 ^ n22852;
  assign n22872 = n22853 & n22871;
  assign n22873 = n22872 ^ n20320;
  assign n22874 = n22873 ^ n22849;
  assign n22875 = n22850 & n22874;
  assign n22876 = n22875 ^ n20370;
  assign n22877 = n22876 ^ n22847;
  assign n22878 = n22848 & n22877;
  assign n22879 = n22878 ^ n20378;
  assign n22881 = n22880 ^ n22879;
  assign n22882 = n22879 ^ n20364;
  assign n22883 = n22881 & ~n22882;
  assign n22884 = n22883 ^ n20364;
  assign n22885 = n22884 ^ n22844;
  assign n22886 = n22845 & ~n22885;
  assign n22887 = n22886 ^ n20388;
  assign n22985 = n22887 ^ n20362;
  assign n22723 = n22722 ^ n22540;
  assign n22724 = n22597 & n22723;
  assign n22725 = n22724 ^ n22596;
  assign n22592 = n21701 ^ n20330;
  assign n22593 = n22592 ^ n22080;
  assign n22591 = n22404 ^ n22382;
  assign n22594 = n22593 ^ n22591;
  assign n22842 = n22725 ^ n22594;
  assign n22986 = n22985 ^ n22842;
  assign n22966 = n22884 ^ n22845;
  assign n22967 = n22870 ^ n22853;
  assign n22534 = n22533 ^ n20157;
  assign n22968 = n22856 ^ n22855;
  assign n22969 = ~n22534 & n22968;
  assign n22970 = n22862 ^ n20215;
  assign n22971 = n22970 ^ n22859;
  assign n22972 = n22969 & n22971;
  assign n22973 = n22867 ^ n20300;
  assign n22974 = n22973 ^ n22865;
  assign n22975 = n22972 & n22974;
  assign n22976 = ~n22967 & n22975;
  assign n22977 = n22873 ^ n20370;
  assign n22978 = n22977 ^ n22849;
  assign n22979 = ~n22976 & ~n22978;
  assign n22980 = n22876 ^ n22848;
  assign n22981 = ~n22979 & ~n22980;
  assign n22982 = n22881 ^ n20364;
  assign n22983 = ~n22981 & ~n22982;
  assign n22984 = n22966 & n22983;
  assign n23093 = n22986 ^ n22984;
  assign n23094 = n23093 ^ n2131;
  assign n23095 = n22983 ^ n22966;
  assign n23096 = n23095 ^ n2121;
  assign n23137 = n22982 ^ n22981;
  assign n23097 = n22980 ^ n22979;
  assign n23101 = n23100 ^ n23097;
  assign n23102 = n22978 ^ n22976;
  assign n23103 = n23102 ^ n1653;
  assign n23104 = n22974 ^ n22972;
  assign n23105 = n23104 ^ n1579;
  assign n23115 = n22971 ^ n22969;
  assign n23109 = n22534 & n22537;
  assign n23110 = n23109 ^ n23108;
  assign n23111 = n22968 ^ n22534;
  assign n23112 = n23111 ^ n23108;
  assign n23113 = n23110 & n23112;
  assign n23114 = n23113 ^ n23109;
  assign n23116 = n23115 ^ n23114;
  assign n23120 = n23119 ^ n23115;
  assign n23121 = ~n23116 & n23120;
  assign n23122 = n23121 ^ n23119;
  assign n23123 = n23122 ^ n23104;
  assign n23124 = n23105 & ~n23123;
  assign n23125 = n23124 ^ n1579;
  assign n23126 = n23125 ^ n1591;
  assign n23127 = n22975 ^ n22967;
  assign n23128 = n23127 ^ n23125;
  assign n23129 = n23126 & n23128;
  assign n23130 = n23129 ^ n1591;
  assign n23131 = n23130 ^ n1653;
  assign n23132 = ~n23103 & ~n23131;
  assign n23133 = n23132 ^ n23102;
  assign n23134 = n23133 ^ n23097;
  assign n23135 = n23101 & n23134;
  assign n23136 = n23135 ^ n23100;
  assign n23138 = n23137 ^ n23136;
  assign n23139 = n23137 ^ n1760;
  assign n23140 = n23138 & ~n23139;
  assign n23141 = n23140 ^ n1760;
  assign n23142 = n23141 ^ n23095;
  assign n23143 = ~n23096 & n23142;
  assign n23144 = n23143 ^ n2121;
  assign n23145 = n23144 ^ n23093;
  assign n23146 = n23094 & ~n23145;
  assign n23147 = n23146 ^ n2131;
  assign n22731 = n21661 ^ n20877;
  assign n22732 = n22731 ^ n21650;
  assign n22729 = n22412 ^ n22409;
  assign n22726 = n22725 ^ n22591;
  assign n22727 = ~n22594 & n22726;
  assign n22728 = n22727 ^ n22593;
  assign n22730 = n22729 ^ n22728;
  assign n22891 = n22732 ^ n22730;
  assign n22843 = n22842 ^ n20362;
  assign n22888 = n22887 ^ n22842;
  assign n22889 = ~n22843 & ~n22888;
  assign n22890 = n22889 ^ n20362;
  assign n22892 = n22891 ^ n22890;
  assign n22988 = n22892 ^ n20358;
  assign n22987 = n22984 & ~n22986;
  assign n23091 = n22988 ^ n22987;
  assign n23092 = n23091 ^ n2146;
  assign n23493 = n23147 ^ n23092;
  assign n23494 = n23493 ^ n21648;
  assign n22573 = n22442 ^ n22439;
  assign n23495 = n23494 ^ n22573;
  assign n23244 = n22057 ^ n21420;
  assign n23245 = n23244 ^ n22598;
  assign n23042 = n21278 ^ n1538;
  assign n23043 = n23042 ^ n2323;
  assign n23044 = n23043 ^ n2414;
  assign n22556 = n21973 ^ n21318;
  assign n22557 = n22556 ^ n22518;
  assign n22555 = n22469 ^ n22364;
  assign n22558 = n22557 ^ n22555;
  assign n22560 = n21949 ^ n21292;
  assign n22561 = n22560 ^ n22337;
  assign n22559 = n22466 ^ n22369;
  assign n22562 = n22561 ^ n22559;
  assign n22564 = n21931 ^ n21268;
  assign n22565 = n22564 ^ n22323;
  assign n22563 = n22463 ^ n22460;
  assign n22566 = n22565 ^ n22563;
  assign n22768 = n22455 ^ n605;
  assign n22568 = n21808 ^ n21120;
  assign n22569 = n22568 ^ n22294;
  assign n22567 = n22450 ^ n22447;
  assign n22570 = n22569 ^ n22567;
  assign n22571 = n21748 ^ n21070;
  assign n22572 = n22571 ^ n22279;
  assign n22574 = n22573 ^ n22572;
  assign n22577 = n22434 ^ n22433;
  assign n22575 = n21741 ^ n20975;
  assign n22576 = n22575 ^ n22225;
  assign n22578 = n22577 ^ n22576;
  assign n22581 = n22429 ^ n22371;
  assign n22579 = n21646 ^ n20862;
  assign n22580 = n22579 ^ n22113;
  assign n22582 = n22581 ^ n22580;
  assign n22585 = n22426 ^ n22373;
  assign n22583 = n21692 ^ n20866;
  assign n22584 = n22583 ^ n21644;
  assign n22586 = n22585 ^ n22584;
  assign n22746 = n22423 ^ n22375;
  assign n22589 = n22420 ^ n22377;
  assign n22587 = n21694 ^ n20870;
  assign n22588 = n22587 ^ n21648;
  assign n22590 = n22589 ^ n22588;
  assign n22736 = n22417 ^ n1860;
  assign n22733 = n22732 ^ n22729;
  assign n22734 = ~n22730 & n22733;
  assign n22735 = n22734 ^ n22732;
  assign n22737 = n22736 ^ n22735;
  assign n22738 = n21656 ^ n20874;
  assign n22739 = n22738 ^ n22090;
  assign n22740 = n22739 ^ n22736;
  assign n22741 = n22737 & n22740;
  assign n22742 = n22741 ^ n22739;
  assign n22743 = n22742 ^ n22589;
  assign n22744 = n22590 & ~n22743;
  assign n22745 = n22744 ^ n22588;
  assign n22747 = n22746 ^ n22745;
  assign n22748 = n21652 ^ n20962;
  assign n22749 = n22748 ^ n22100;
  assign n22750 = n22749 ^ n22746;
  assign n22751 = ~n22747 & n22750;
  assign n22752 = n22751 ^ n22749;
  assign n22753 = n22752 ^ n22585;
  assign n22754 = ~n22586 & n22753;
  assign n22755 = n22754 ^ n22584;
  assign n22756 = n22755 ^ n22581;
  assign n22757 = n22582 & n22756;
  assign n22758 = n22757 ^ n22580;
  assign n22759 = n22758 ^ n22577;
  assign n22760 = n22578 & ~n22759;
  assign n22761 = n22760 ^ n22576;
  assign n22762 = n22761 ^ n22572;
  assign n22763 = n22574 & ~n22762;
  assign n22764 = n22763 ^ n22573;
  assign n22765 = n22764 ^ n22567;
  assign n22766 = n22570 & n22765;
  assign n22767 = n22766 ^ n22569;
  assign n22769 = n22768 ^ n22767;
  assign n22770 = n21911 ^ n21249;
  assign n22771 = n22770 ^ n22309;
  assign n22772 = n22771 ^ n22768;
  assign n22773 = ~n22769 & n22772;
  assign n22774 = n22773 ^ n22771;
  assign n22775 = n22774 ^ n22565;
  assign n22776 = ~n22566 & ~n22775;
  assign n22777 = n22776 ^ n22563;
  assign n22778 = n22777 ^ n22559;
  assign n22779 = n22562 & ~n22778;
  assign n22780 = n22779 ^ n22561;
  assign n22781 = n22780 ^ n22555;
  assign n22782 = ~n22558 & n22781;
  assign n22783 = n22782 ^ n22557;
  assign n22554 = n22477 ^ n22474;
  assign n22784 = n22783 ^ n22554;
  assign n22785 = n22001 ^ n21346;
  assign n22786 = n22785 ^ n22614;
  assign n22787 = n22786 ^ n22554;
  assign n22788 = ~n22784 & n22787;
  assign n22789 = n22788 ^ n22786;
  assign n22550 = n22026 ^ n21383;
  assign n22552 = n22551 ^ n22550;
  assign n22549 = n22482 ^ n22481;
  assign n22553 = n22552 ^ n22549;
  assign n22813 = n22789 ^ n22553;
  assign n22814 = n22813 ^ n20767;
  assign n22815 = n22786 ^ n22784;
  assign n22816 = n22815 ^ n20698;
  assign n22817 = n22780 ^ n22557;
  assign n22818 = n22817 ^ n22555;
  assign n22819 = n22818 ^ n20540;
  assign n22820 = n22777 ^ n22562;
  assign n22821 = n22820 ^ n20448;
  assign n22822 = n22774 ^ n22566;
  assign n22823 = n22822 ^ n20334;
  assign n22824 = n22771 ^ n22769;
  assign n22825 = n22824 ^ n20335;
  assign n22917 = n22764 ^ n22570;
  assign n22826 = n22761 ^ n22574;
  assign n22827 = n22826 ^ n20340;
  assign n22828 = n22758 ^ n22576;
  assign n22829 = n22828 ^ n22577;
  assign n22830 = n22829 ^ n20423;
  assign n22831 = n22755 ^ n22582;
  assign n22832 = n22831 ^ n20344;
  assign n22833 = n22752 ^ n22586;
  assign n22834 = n22833 ^ n20348;
  assign n22835 = n22749 ^ n22747;
  assign n22836 = n22835 ^ n20410;
  assign n22837 = n22742 ^ n22588;
  assign n22838 = n22837 ^ n22589;
  assign n22839 = n22838 ^ n20354;
  assign n22840 = n22739 ^ n22737;
  assign n22841 = n22840 ^ n19749;
  assign n22893 = n22891 ^ n20358;
  assign n22894 = ~n22892 & ~n22893;
  assign n22895 = n22894 ^ n20358;
  assign n22896 = n22895 ^ n22840;
  assign n22897 = n22841 & n22896;
  assign n22898 = n22897 ^ n19749;
  assign n22899 = n22898 ^ n22838;
  assign n22900 = ~n22839 & n22899;
  assign n22901 = n22900 ^ n20354;
  assign n22902 = n22901 ^ n22835;
  assign n22903 = ~n22836 & n22902;
  assign n22904 = n22903 ^ n20410;
  assign n22905 = n22904 ^ n22833;
  assign n22906 = n22834 & ~n22905;
  assign n22907 = n22906 ^ n20348;
  assign n22908 = n22907 ^ n22831;
  assign n22909 = ~n22832 & n22908;
  assign n22910 = n22909 ^ n20344;
  assign n22911 = n22910 ^ n22829;
  assign n22912 = ~n22830 & ~n22911;
  assign n22913 = n22912 ^ n20423;
  assign n22914 = n22913 ^ n22826;
  assign n22915 = n22827 & n22914;
  assign n22916 = n22915 ^ n20340;
  assign n22918 = n22917 ^ n22916;
  assign n22919 = n22917 ^ n20338;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = n22920 ^ n20338;
  assign n22922 = n22921 ^ n22824;
  assign n22923 = ~n22825 & ~n22922;
  assign n22924 = n22923 ^ n20335;
  assign n22925 = n22924 ^ n22822;
  assign n22926 = n22823 & ~n22925;
  assign n22927 = n22926 ^ n20334;
  assign n22928 = n22927 ^ n22820;
  assign n22929 = n22821 & ~n22928;
  assign n22930 = n22929 ^ n20448;
  assign n22931 = n22930 ^ n22818;
  assign n22932 = n22819 & n22931;
  assign n22933 = n22932 ^ n20540;
  assign n22934 = n22933 ^ n22815;
  assign n22935 = ~n22816 & n22934;
  assign n22936 = n22935 ^ n20698;
  assign n22937 = n22936 ^ n22813;
  assign n22938 = ~n22814 & n22937;
  assign n22939 = n22938 ^ n20767;
  assign n22959 = n22939 ^ n20121;
  assign n22794 = n21279 ^ n20715;
  assign n22795 = n22794 ^ n22645;
  assign n22790 = n22789 ^ n22552;
  assign n22791 = n22553 & n22790;
  assign n22792 = n22791 ^ n22549;
  assign n22547 = n22485 ^ n800;
  assign n22548 = n22547 ^ n22486;
  assign n22793 = n22792 ^ n22548;
  assign n22811 = n22795 ^ n22793;
  assign n22960 = n22959 ^ n22811;
  assign n22961 = n22913 ^ n20340;
  assign n22962 = n22961 ^ n22826;
  assign n22963 = n22907 ^ n22832;
  assign n22964 = n22898 ^ n20354;
  assign n22965 = n22964 ^ n22838;
  assign n22989 = ~n22987 & ~n22988;
  assign n22990 = n22895 ^ n22841;
  assign n22991 = ~n22989 & n22990;
  assign n22992 = ~n22965 & ~n22991;
  assign n22993 = n22901 ^ n20410;
  assign n22994 = n22993 ^ n22835;
  assign n22995 = ~n22992 & n22994;
  assign n22996 = n22904 ^ n22834;
  assign n22997 = n22995 & ~n22996;
  assign n22998 = n22963 & n22997;
  assign n22999 = n22910 ^ n22830;
  assign n23000 = n22998 & n22999;
  assign n23001 = ~n22962 & ~n23000;
  assign n23002 = n22918 ^ n20338;
  assign n23003 = n23001 & ~n23002;
  assign n23004 = n22921 ^ n20335;
  assign n23005 = n23004 ^ n22824;
  assign n23006 = ~n23003 & ~n23005;
  assign n23007 = n22924 ^ n20334;
  assign n23008 = n23007 ^ n22822;
  assign n23009 = n23006 & ~n23008;
  assign n23010 = n22927 ^ n22821;
  assign n23011 = ~n23009 & n23010;
  assign n23012 = n22930 ^ n20540;
  assign n23013 = n23012 ^ n22818;
  assign n23014 = ~n23011 & ~n23013;
  assign n23015 = n22933 ^ n22816;
  assign n23016 = n23014 & ~n23015;
  assign n23017 = n22936 ^ n20767;
  assign n23018 = n23017 ^ n22813;
  assign n23019 = ~n23016 & n23018;
  assign n23020 = n22960 & ~n23019;
  assign n22812 = n22811 ^ n20121;
  assign n22940 = n22939 ^ n22811;
  assign n22941 = n22812 & ~n22940;
  assign n22942 = n22941 ^ n20121;
  assign n22796 = n22795 ^ n22548;
  assign n22797 = n22793 & n22796;
  assign n22798 = n22797 ^ n22795;
  assign n22543 = n21303 ^ n20718;
  assign n22545 = n22544 ^ n22543;
  assign n22808 = n22798 ^ n22545;
  assign n22542 = n22492 ^ n882;
  assign n22809 = n22808 ^ n22542;
  assign n22810 = n22809 ^ n20126;
  assign n23021 = n22942 ^ n22810;
  assign n23022 = n23020 & n23021;
  assign n22943 = n22942 ^ n22809;
  assign n22944 = n22810 & ~n22943;
  assign n22945 = n22944 ^ n20126;
  assign n22803 = n21329 ^ n20722;
  assign n22804 = n22803 ^ n21938;
  assign n22802 = n22495 ^ n22359;
  assign n22805 = n22804 ^ n22802;
  assign n22546 = n22545 ^ n22542;
  assign n22799 = n22798 ^ n22542;
  assign n22800 = ~n22546 & ~n22799;
  assign n22801 = n22800 ^ n22545;
  assign n22806 = n22805 ^ n22801;
  assign n22807 = n22806 ^ n20130;
  assign n23023 = n22945 ^ n22807;
  assign n23024 = n23022 & ~n23023;
  assign n22953 = n21358 ^ n20707;
  assign n22954 = n22953 ^ n21960;
  assign n22952 = n22498 ^ n22357;
  assign n22955 = n22954 ^ n22952;
  assign n22949 = n22802 ^ n22801;
  assign n22950 = ~n22805 & ~n22949;
  assign n22951 = n22950 ^ n22804;
  assign n22956 = n22955 ^ n22951;
  assign n22957 = n22956 ^ n20137;
  assign n22946 = n22945 ^ n22806;
  assign n22947 = ~n22807 & n22946;
  assign n22948 = n22947 ^ n20130;
  assign n22958 = n22957 ^ n22948;
  assign n23041 = n23024 ^ n22958;
  assign n23045 = n23044 ^ n23041;
  assign n23046 = n23021 ^ n23020;
  assign n23047 = n23046 ^ n1336;
  assign n23048 = n23019 ^ n22960;
  assign n1319 = n1309 ^ n1219;
  assign n1320 = n1319 ^ n1152;
  assign n1324 = n1323 ^ n1320;
  assign n23049 = n23048 ^ n1324;
  assign n23199 = n23018 ^ n23016;
  assign n23194 = n23015 ^ n23014;
  assign n23050 = n23013 ^ n23011;
  assign n23051 = n23050 ^ n1002;
  assign n23052 = n23010 ^ n23009;
  assign n23053 = n23052 ^ n990;
  assign n23054 = n23008 ^ n23006;
  assign n23058 = n23057 ^ n23054;
  assign n23059 = n23005 ^ n23003;
  assign n23063 = n23062 ^ n23059;
  assign n23177 = n23002 ^ n23001;
  assign n23065 = n21143 ^ n14192;
  assign n23066 = n23065 ^ n643;
  assign n23067 = n23066 ^ n547;
  assign n23064 = n23000 ^ n22962;
  assign n23068 = n23067 ^ n23064;
  assign n23069 = n22999 ^ n22998;
  assign n23070 = n23069 ^ n639;
  assign n23071 = n22997 ^ n22963;
  assign n23075 = n23074 ^ n23071;
  assign n23076 = n22994 ^ n22992;
  assign n23080 = n23079 ^ n23076;
  assign n23081 = n22991 ^ n22965;
  assign n23085 = n23084 ^ n23081;
  assign n23086 = n22990 ^ n22989;
  assign n23090 = n23089 ^ n23086;
  assign n23148 = n23147 ^ n23091;
  assign n23149 = n23092 & ~n23148;
  assign n23150 = n23149 ^ n2146;
  assign n23151 = n23150 ^ n23086;
  assign n23152 = n23090 & ~n23151;
  assign n23153 = n23152 ^ n23089;
  assign n23154 = n23153 ^ n23081;
  assign n23155 = n23085 & ~n23154;
  assign n23156 = n23155 ^ n23084;
  assign n23157 = n23156 ^ n23076;
  assign n23158 = n23080 & ~n23157;
  assign n23159 = n23158 ^ n23079;
  assign n23163 = n23162 ^ n23159;
  assign n23164 = n22996 ^ n22995;
  assign n23165 = n23164 ^ n23159;
  assign n23166 = n23163 & ~n23165;
  assign n23167 = n23166 ^ n23162;
  assign n23168 = n23167 ^ n23071;
  assign n23169 = ~n23075 & n23168;
  assign n23170 = n23169 ^ n23074;
  assign n23171 = n23170 ^ n23069;
  assign n23172 = ~n23070 & n23171;
  assign n23173 = n23172 ^ n639;
  assign n23174 = n23173 ^ n23064;
  assign n23175 = n23068 & ~n23174;
  assign n23176 = n23175 ^ n23067;
  assign n23178 = n23177 ^ n23176;
  assign n23179 = n23177 ^ n554;
  assign n23180 = n23178 & ~n23179;
  assign n23181 = n23180 ^ n554;
  assign n23182 = n23181 ^ n23059;
  assign n23183 = ~n23063 & n23182;
  assign n23184 = n23183 ^ n23062;
  assign n23185 = n23184 ^ n23054;
  assign n23186 = n23058 & ~n23185;
  assign n23187 = n23186 ^ n23057;
  assign n23188 = n23187 ^ n23052;
  assign n23189 = ~n23053 & n23188;
  assign n23190 = n23189 ^ n990;
  assign n23191 = n23190 ^ n23050;
  assign n23192 = ~n23051 & n23191;
  assign n23193 = n23192 ^ n1002;
  assign n23195 = n23194 ^ n23193;
  assign n1015 = n975 ^ n939;
  assign n1016 = n1015 ^ n1009;
  assign n1020 = n1019 ^ n1016;
  assign n23196 = n23194 ^ n1020;
  assign n23197 = ~n23195 & n23196;
  assign n23198 = n23197 ^ n1020;
  assign n23200 = n23199 ^ n23198;
  assign n23201 = n23199 ^ n1145;
  assign n23202 = n23200 & ~n23201;
  assign n23203 = n23202 ^ n1145;
  assign n23204 = n23203 ^ n23048;
  assign n23205 = n23049 & ~n23204;
  assign n23206 = n23205 ^ n1324;
  assign n23207 = n23206 ^ n23046;
  assign n23208 = ~n23047 & n23207;
  assign n23209 = n23208 ^ n1336;
  assign n2310 = n2309 ^ n2273;
  assign n2311 = n2310 ^ n2306;
  assign n2315 = n2314 ^ n2311;
  assign n23210 = n23209 ^ n2315;
  assign n23211 = n23023 ^ n23022;
  assign n23212 = n23211 ^ n2315;
  assign n23213 = ~n23210 & n23212;
  assign n23214 = n23213 ^ n23211;
  assign n23215 = n23214 ^ n23044;
  assign n23216 = n23045 & ~n23215;
  assign n23217 = n23216 ^ n23041;
  assign n23033 = n21388 ^ n20772;
  assign n23034 = n23033 ^ n21983;
  assign n23030 = n22952 ^ n22951;
  assign n23031 = ~n22955 & ~n23030;
  assign n23032 = n23031 ^ n22954;
  assign n23035 = n23034 ^ n23032;
  assign n23029 = n22501 ^ n22355;
  assign n23036 = n23035 ^ n23029;
  assign n23026 = n22956 ^ n22948;
  assign n23027 = n22957 & ~n23026;
  assign n23028 = n23027 ^ n20137;
  assign n23037 = n23036 ^ n23028;
  assign n23038 = n23037 ^ n20115;
  assign n23025 = ~n22958 & ~n23024;
  assign n23039 = n23038 ^ n23025;
  assign n2427 = n2426 ^ n2363;
  assign n2428 = n2427 ^ n2420;
  assign n2429 = n2428 ^ n1511;
  assign n23040 = n23039 ^ n2429;
  assign n23243 = n23217 ^ n23040;
  assign n23246 = n23245 ^ n23243;
  assign n23249 = n23211 ^ n23210;
  assign n23250 = n21674 ^ n20856;
  assign n23251 = n23250 ^ n22606;
  assign n23252 = n23249 & n23251;
  assign n23247 = n21670 ^ n20855;
  assign n23248 = n23247 ^ n22602;
  assign n23253 = n23252 ^ n23248;
  assign n23254 = n23214 ^ n23045;
  assign n23255 = n23254 ^ n23248;
  assign n23256 = n23253 & ~n23255;
  assign n23257 = n23256 ^ n23252;
  assign n23258 = n23257 ^ n23243;
  assign n23259 = ~n23246 & n23258;
  assign n23260 = n23259 ^ n23245;
  assign n23236 = n23036 ^ n20115;
  assign n23237 = n23037 & ~n23236;
  assign n23238 = n23237 ^ n20115;
  assign n23232 = n21395 ^ n20818;
  assign n23233 = n23232 ^ n22012;
  assign n23227 = n23034 ^ n23029;
  assign n23228 = n23032 ^ n23029;
  assign n23229 = ~n23227 & n23228;
  assign n23230 = n23229 ^ n23034;
  assign n23226 = n22504 ^ n22350;
  assign n23231 = n23230 ^ n23226;
  assign n23234 = n23233 ^ n23231;
  assign n23235 = n23234 ^ n20147;
  assign n23239 = n23238 ^ n23235;
  assign n23225 = ~n23025 & ~n23038;
  assign n23240 = n23239 ^ n23225;
  assign n23221 = n21328 ^ n2589;
  assign n23222 = n23221 ^ n1544;
  assign n23223 = n23222 ^ n2559;
  assign n23218 = n23217 ^ n23039;
  assign n23219 = ~n23040 & n23218;
  assign n23220 = n23219 ^ n2429;
  assign n23224 = n23223 ^ n23220;
  assign n23241 = n23240 ^ n23224;
  assign n22539 = n21668 ^ n20850;
  assign n22541 = n22540 ^ n22539;
  assign n23242 = n23241 ^ n22541;
  assign n23320 = n23260 ^ n23242;
  assign n23321 = n23320 ^ n20906;
  assign n23322 = n23251 ^ n23249;
  assign n23323 = n20889 & n23322;
  assign n23324 = n23323 ^ n20882;
  assign n23325 = n23254 ^ n23253;
  assign n23326 = n23325 ^ n23323;
  assign n23327 = n23324 & ~n23326;
  assign n23328 = n23327 ^ n20882;
  assign n23329 = n23328 ^ n20899;
  assign n23330 = n23257 ^ n23246;
  assign n23331 = n23330 ^ n23328;
  assign n23332 = n23329 & n23331;
  assign n23333 = n23332 ^ n20899;
  assign n23334 = n23333 ^ n23320;
  assign n23335 = n23321 & ~n23334;
  assign n23336 = n23335 ^ n20906;
  assign n23368 = n23336 ^ n20913;
  assign n23289 = n22067 ^ n20849;
  assign n23290 = n23289 ^ n22591;
  assign n23281 = n23280 ^ n22678;
  assign n23282 = n23281 ^ n20857;
  assign n23276 = n23225 & ~n23239;
  assign n23275 = n22507 ^ n22348;
  assign n23277 = n23276 ^ n23275;
  assign n23283 = n23282 ^ n23277;
  assign n23284 = n23283 ^ n22035;
  assign n23272 = n23233 ^ n23226;
  assign n23273 = n23231 & ~n23272;
  assign n23274 = n23273 ^ n23233;
  assign n23285 = n23284 ^ n23274;
  assign n23268 = n23240 ^ n23223;
  assign n23269 = n23240 ^ n23220;
  assign n23270 = n23268 & ~n23269;
  assign n23271 = n23270 ^ n23223;
  assign n23286 = n23285 ^ n23271;
  assign n23264 = n23238 ^ n20147;
  assign n23265 = n23238 ^ n23234;
  assign n23266 = n23264 & n23265;
  assign n23267 = n23266 ^ n20147;
  assign n23287 = n23286 ^ n23267;
  assign n23261 = n23260 ^ n22541;
  assign n23262 = n23242 & ~n23261;
  assign n23263 = n23262 ^ n23241;
  assign n23288 = n23287 ^ n23263;
  assign n23318 = n23290 ^ n23288;
  assign n23369 = n23368 ^ n23318;
  assign n23361 = n23330 ^ n23329;
  assign n23362 = n23325 ^ n23324;
  assign n23363 = n23322 ^ n20889;
  assign n23364 = n23362 & n23363;
  assign n23365 = ~n23361 & n23364;
  assign n23366 = n23333 ^ n23321;
  assign n23367 = n23365 & n23366;
  assign n23387 = n23369 ^ n23367;
  assign n23388 = n23387 ^ n23386;
  assign n23389 = n23366 ^ n23365;
  assign n23393 = n23392 ^ n23389;
  assign n1551 = n1550 ^ n1427;
  assign n1552 = n1551 ^ n1520;
  assign n1553 = n1552 ^ n1463;
  assign n23394 = n1553 & ~n23363;
  assign n23398 = n23397 ^ n23394;
  assign n23399 = n23363 ^ n23362;
  assign n23400 = n23399 ^ n23394;
  assign n23401 = n23398 & ~n23400;
  assign n23402 = n23401 ^ n23397;
  assign n23406 = n23405 ^ n23402;
  assign n23407 = n23364 ^ n23361;
  assign n23408 = n23407 ^ n23402;
  assign n23409 = n23406 & n23408;
  assign n23410 = n23409 ^ n23405;
  assign n23411 = n23410 ^ n23389;
  assign n23412 = n23393 & ~n23411;
  assign n23413 = n23412 ^ n23392;
  assign n23414 = n23413 ^ n23387;
  assign n23415 = n23388 & ~n23414;
  assign n23416 = n23415 ^ n23386;
  assign n23319 = n23318 ^ n20913;
  assign n23337 = n23336 ^ n23318;
  assign n23338 = n23319 & ~n23337;
  assign n23339 = n23338 ^ n20913;
  assign n23295 = n22729 ^ n21491;
  assign n23296 = n23295 ^ n21663;
  assign n23291 = n23290 ^ n23287;
  assign n23292 = ~n23288 & n23291;
  assign n23293 = n23292 ^ n23290;
  assign n22538 = n22537 ^ n22534;
  assign n23294 = n23293 ^ n22538;
  assign n23316 = n23296 ^ n23294;
  assign n23317 = n23316 ^ n20920;
  assign n23371 = n23339 ^ n23317;
  assign n23370 = n23367 & n23369;
  assign n23382 = n23371 ^ n23370;
  assign n23383 = n23382 ^ n1724;
  assign n23492 = n23416 ^ n23383;
  assign n23496 = n23495 ^ n23492;
  assign n23498 = n23144 ^ n23094;
  assign n23499 = n23498 ^ n22090;
  assign n23500 = n23499 ^ n22577;
  assign n23497 = n23413 ^ n23388;
  assign n23501 = n23500 ^ n23497;
  assign n23505 = n23410 ^ n23393;
  assign n23502 = n23141 ^ n23096;
  assign n23503 = n23502 ^ n21650;
  assign n23504 = n23503 ^ n22581;
  assign n23506 = n23505 ^ n23504;
  assign n23508 = n23138 ^ n1760;
  assign n23509 = n23508 ^ n22080;
  assign n23510 = n23509 ^ n22585;
  assign n23507 = n23407 ^ n23406;
  assign n23511 = n23510 ^ n23507;
  assign n23513 = n23133 ^ n23101;
  assign n23514 = n23513 ^ n21658;
  assign n23515 = n23514 ^ n22746;
  assign n23512 = n23399 ^ n23398;
  assign n23516 = n23515 ^ n23512;
  assign n23518 = n22589 ^ n21663;
  assign n23465 = n23130 ^ n23103;
  assign n23519 = n23518 ^ n23465;
  assign n23517 = n23363 ^ n1553;
  assign n23520 = n23519 ^ n23517;
  assign n23948 = n22736 ^ n22067;
  assign n23439 = n23127 ^ n1591;
  assign n23440 = n23439 ^ n23125;
  assign n23949 = n23948 ^ n23440;
  assign n23757 = n21679 ^ n21395;
  assign n23758 = n23757 ^ n22691;
  assign n23755 = n23203 ^ n23049;
  assign n23649 = n23200 ^ n1145;
  assign n23646 = n22035 ^ n21388;
  assign n23647 = n23646 ^ n22693;
  assign n23751 = n23649 ^ n23647;
  assign n23523 = n22701 ^ n22012;
  assign n23524 = n23523 ^ n21358;
  assign n23521 = n23193 ^ n1020;
  assign n23522 = n23521 ^ n23194;
  assign n23525 = n23524 ^ n23522;
  assign n23527 = n22530 ^ n21983;
  assign n23528 = n23527 ^ n21329;
  assign n23526 = n23190 ^ n23051;
  assign n23529 = n23528 ^ n23526;
  assign n23531 = n21960 ^ n21303;
  assign n23532 = n23531 ^ n23275;
  assign n23530 = n23187 ^ n23053;
  assign n23533 = n23532 ^ n23530;
  assign n23535 = n23226 ^ n21938;
  assign n23536 = n23535 ^ n21279;
  assign n23534 = n23184 ^ n23058;
  assign n23537 = n23536 ^ n23534;
  assign n23540 = n23029 ^ n22026;
  assign n23541 = n23540 ^ n22544;
  assign n23538 = n23181 ^ n23062;
  assign n23539 = n23538 ^ n23059;
  assign n23542 = n23541 ^ n23539;
  assign n23545 = n23178 ^ n554;
  assign n23543 = n22645 ^ n22001;
  assign n23544 = n23543 ^ n22952;
  assign n23546 = n23545 ^ n23544;
  assign n23549 = n23173 ^ n23067;
  assign n23550 = n23549 ^ n23064;
  assign n23547 = n22802 ^ n22551;
  assign n23548 = n23547 ^ n21973;
  assign n23551 = n23550 ^ n23548;
  assign n23554 = n23170 ^ n23070;
  assign n23552 = n22614 ^ n21949;
  assign n23553 = n23552 ^ n22542;
  assign n23555 = n23554 ^ n23553;
  assign n23556 = n22518 ^ n21931;
  assign n23557 = n23556 ^ n22548;
  assign n23470 = n23167 ^ n23075;
  assign n23558 = n23557 ^ n23470;
  assign n23561 = n22337 ^ n21911;
  assign n23562 = n23561 ^ n22549;
  assign n23559 = n23164 ^ n23162;
  assign n23560 = n23559 ^ n23159;
  assign n23563 = n23562 ^ n23560;
  assign n23564 = n22554 ^ n21808;
  assign n23565 = n23564 ^ n22323;
  assign n23475 = n23156 ^ n23080;
  assign n23566 = n23565 ^ n23475;
  assign n23567 = n22555 ^ n21748;
  assign n23568 = n23567 ^ n22309;
  assign n23482 = n23153 ^ n23085;
  assign n23569 = n23568 ^ n23482;
  assign n23570 = n22559 ^ n22294;
  assign n23571 = n23570 ^ n21741;
  assign n23488 = n23150 ^ n23089;
  assign n23489 = n23488 ^ n23086;
  assign n23572 = n23571 ^ n23489;
  assign n23573 = n22563 ^ n21646;
  assign n23574 = n23573 ^ n22279;
  assign n23575 = n23574 ^ n23493;
  assign n23576 = n22573 ^ n21694;
  assign n23577 = n23576 ^ n21644;
  assign n23578 = n23577 ^ n23508;
  assign n23462 = n22581 ^ n21661;
  assign n23463 = n23462 ^ n21648;
  assign n23579 = n23465 ^ n23463;
  assign n23437 = n22585 ^ n22090;
  assign n23438 = n23437 ^ n21701;
  assign n23441 = n23440 ^ n23438;
  assign n23355 = n22746 ^ n21650;
  assign n23356 = n23355 ^ n21666;
  assign n23353 = n23122 ^ n1579;
  assign n23354 = n23353 ^ n23104;
  assign n23357 = n23356 ^ n23354;
  assign n23309 = n22589 ^ n21631;
  assign n23310 = n23309 ^ n22080;
  assign n23307 = n23119 ^ n23114;
  assign n23308 = n23307 ^ n23115;
  assign n23311 = n23310 ^ n23308;
  assign n23300 = n23111 ^ n23110;
  assign n23297 = n23296 ^ n22538;
  assign n23298 = ~n23294 & ~n23297;
  assign n23299 = n23298 ^ n23296;
  assign n23301 = n23300 ^ n23299;
  assign n23302 = n22736 ^ n21527;
  assign n23303 = n23302 ^ n21658;
  assign n23304 = n23303 ^ n23300;
  assign n23305 = ~n23301 & ~n23304;
  assign n23306 = n23305 ^ n23303;
  assign n23350 = n23308 ^ n23306;
  assign n23351 = n23311 & ~n23350;
  assign n23352 = n23351 ^ n23310;
  assign n23434 = n23356 ^ n23352;
  assign n23435 = ~n23357 & n23434;
  assign n23436 = n23435 ^ n23354;
  assign n23459 = n23440 ^ n23436;
  assign n23460 = ~n23441 & n23459;
  assign n23461 = n23460 ^ n23438;
  assign n23580 = n23465 ^ n23461;
  assign n23581 = ~n23579 & n23580;
  assign n23582 = n23581 ^ n23463;
  assign n23583 = n23582 ^ n23513;
  assign n23584 = n22577 ^ n22100;
  assign n23585 = n23584 ^ n21656;
  assign n23586 = n23585 ^ n23513;
  assign n23587 = n23583 & ~n23586;
  assign n23588 = n23587 ^ n23585;
  assign n23589 = n23588 ^ n23508;
  assign n23590 = ~n23578 & n23589;
  assign n23591 = n23590 ^ n23577;
  assign n23592 = n23591 ^ n23502;
  assign n23593 = n22567 ^ n21652;
  assign n23594 = n23593 ^ n22113;
  assign n23595 = n23594 ^ n23502;
  assign n23596 = n23592 & ~n23595;
  assign n23597 = n23596 ^ n23594;
  assign n23598 = n23597 ^ n23498;
  assign n23599 = n22225 ^ n21692;
  assign n23600 = n23599 ^ n22768;
  assign n23601 = n23600 ^ n23498;
  assign n23602 = ~n23598 & ~n23601;
  assign n23603 = n23602 ^ n23600;
  assign n23604 = n23603 ^ n23493;
  assign n23605 = n23575 & n23604;
  assign n23606 = n23605 ^ n23574;
  assign n23607 = n23606 ^ n23489;
  assign n23608 = n23572 & ~n23607;
  assign n23609 = n23608 ^ n23571;
  assign n23610 = n23609 ^ n23482;
  assign n23611 = n23569 & ~n23610;
  assign n23612 = n23611 ^ n23568;
  assign n23613 = n23612 ^ n23475;
  assign n23614 = n23566 & ~n23613;
  assign n23615 = n23614 ^ n23565;
  assign n23616 = n23615 ^ n23560;
  assign n23617 = n23563 & ~n23616;
  assign n23618 = n23617 ^ n23562;
  assign n23619 = n23618 ^ n23470;
  assign n23620 = n23558 & n23619;
  assign n23621 = n23620 ^ n23557;
  assign n23622 = n23621 ^ n23554;
  assign n23623 = n23555 & ~n23622;
  assign n23624 = n23623 ^ n23553;
  assign n23625 = n23624 ^ n23548;
  assign n23626 = ~n23551 & ~n23625;
  assign n23627 = n23626 ^ n23550;
  assign n23628 = n23627 ^ n23545;
  assign n23629 = n23546 & n23628;
  assign n23630 = n23629 ^ n23544;
  assign n23631 = n23630 ^ n23541;
  assign n23632 = ~n23542 & n23631;
  assign n23633 = n23632 ^ n23539;
  assign n23634 = n23633 ^ n23534;
  assign n23635 = n23537 & n23634;
  assign n23636 = n23635 ^ n23536;
  assign n23637 = n23636 ^ n23530;
  assign n23638 = ~n23533 & n23637;
  assign n23639 = n23638 ^ n23532;
  assign n23640 = n23639 ^ n23528;
  assign n23641 = ~n23529 & ~n23640;
  assign n23642 = n23641 ^ n23526;
  assign n23643 = n23642 ^ n23522;
  assign n23644 = n23525 & n23643;
  assign n23645 = n23644 ^ n23524;
  assign n23752 = n23649 ^ n23645;
  assign n23753 = ~n23751 & n23752;
  assign n23754 = n23753 ^ n23647;
  assign n23756 = n23755 ^ n23754;
  assign n23759 = n23758 ^ n23756;
  assign n23648 = n23647 ^ n23645;
  assign n23650 = n23649 ^ n23648;
  assign n23651 = n23650 ^ n20772;
  assign n23652 = n23642 ^ n23525;
  assign n23653 = n23652 ^ n20707;
  assign n23654 = n23639 ^ n23529;
  assign n23655 = n23654 ^ n20722;
  assign n23656 = n23636 ^ n23533;
  assign n23657 = n23656 ^ n20718;
  assign n23658 = n23633 ^ n23537;
  assign n23659 = n23658 ^ n20715;
  assign n23660 = n23630 ^ n23542;
  assign n23661 = n23660 ^ n21383;
  assign n23662 = n23627 ^ n23546;
  assign n23663 = n23662 ^ n21346;
  assign n23664 = n23624 ^ n23551;
  assign n23665 = n23664 ^ n21318;
  assign n23721 = n23621 ^ n23555;
  assign n23666 = n23618 ^ n23557;
  assign n23667 = n23666 ^ n23470;
  assign n23668 = n23667 ^ n21268;
  assign n23713 = n23615 ^ n23563;
  assign n23669 = n23612 ^ n23566;
  assign n23670 = n23669 ^ n21120;
  assign n23705 = n23609 ^ n23569;
  assign n23700 = n23606 ^ n23572;
  assign n23671 = n23603 ^ n23575;
  assign n23672 = n23671 ^ n20862;
  assign n23692 = n23600 ^ n23598;
  assign n23673 = n23594 ^ n23592;
  assign n23674 = n23673 ^ n20962;
  assign n23675 = n23588 ^ n23578;
  assign n23676 = n23675 ^ n20870;
  assign n23681 = n23585 ^ n23583;
  assign n23464 = n23463 ^ n23461;
  assign n23466 = n23465 ^ n23464;
  assign n23677 = n23466 ^ n20877;
  assign n23442 = n23441 ^ n23436;
  assign n23358 = n23357 ^ n23352;
  assign n23430 = n23358 ^ n20852;
  assign n23312 = n23311 ^ n23306;
  assign n23313 = n23312 ^ n20934;
  assign n23314 = n23303 ^ n23301;
  assign n23315 = n23314 ^ n20927;
  assign n23340 = n23339 ^ n23316;
  assign n23341 = ~n23317 & n23340;
  assign n23342 = n23341 ^ n20920;
  assign n23343 = n23342 ^ n23314;
  assign n23344 = n23315 & ~n23343;
  assign n23345 = n23344 ^ n20927;
  assign n23346 = n23345 ^ n23312;
  assign n23347 = ~n23313 & ~n23346;
  assign n23348 = n23347 ^ n20934;
  assign n23431 = n23358 ^ n23348;
  assign n23432 = n23430 & ~n23431;
  assign n23433 = n23432 ^ n20852;
  assign n23443 = n23442 ^ n23433;
  assign n23455 = n23442 ^ n20330;
  assign n23456 = ~n23443 & n23455;
  assign n23457 = n23456 ^ n20330;
  assign n23678 = n23466 ^ n23457;
  assign n23679 = n23677 & ~n23678;
  assign n23680 = n23679 ^ n20877;
  assign n23682 = n23681 ^ n23680;
  assign n23683 = n23681 ^ n20874;
  assign n23684 = ~n23682 & ~n23683;
  assign n23685 = n23684 ^ n20874;
  assign n23686 = n23685 ^ n23675;
  assign n23687 = n23676 & n23686;
  assign n23688 = n23687 ^ n20870;
  assign n23689 = n23688 ^ n23673;
  assign n23690 = n23674 & ~n23689;
  assign n23691 = n23690 ^ n20962;
  assign n23693 = n23692 ^ n23691;
  assign n23694 = n23692 ^ n20866;
  assign n23695 = ~n23693 & ~n23694;
  assign n23696 = n23695 ^ n20866;
  assign n23697 = n23696 ^ n23671;
  assign n23698 = ~n23672 & n23697;
  assign n23699 = n23698 ^ n20862;
  assign n23701 = n23700 ^ n23699;
  assign n23702 = n23700 ^ n20975;
  assign n23703 = ~n23701 & ~n23702;
  assign n23704 = n23703 ^ n20975;
  assign n23706 = n23705 ^ n23704;
  assign n23707 = n23705 ^ n21070;
  assign n23708 = n23706 & n23707;
  assign n23709 = n23708 ^ n21070;
  assign n23710 = n23709 ^ n23669;
  assign n23711 = n23670 & ~n23710;
  assign n23712 = n23711 ^ n21120;
  assign n23714 = n23713 ^ n23712;
  assign n23715 = n23713 ^ n21249;
  assign n23716 = ~n23714 & n23715;
  assign n23717 = n23716 ^ n21249;
  assign n23718 = n23717 ^ n23667;
  assign n23719 = ~n23668 & ~n23718;
  assign n23720 = n23719 ^ n21268;
  assign n23722 = n23721 ^ n23720;
  assign n23723 = n23721 ^ n21292;
  assign n23724 = ~n23722 & n23723;
  assign n23725 = n23724 ^ n21292;
  assign n23726 = n23725 ^ n23664;
  assign n23727 = n23665 & n23726;
  assign n23728 = n23727 ^ n21318;
  assign n23729 = n23728 ^ n23662;
  assign n23730 = n23663 & ~n23729;
  assign n23731 = n23730 ^ n21346;
  assign n23732 = n23731 ^ n23660;
  assign n23733 = ~n23661 & ~n23732;
  assign n23734 = n23733 ^ n21383;
  assign n23735 = n23734 ^ n23658;
  assign n23736 = n23659 & ~n23735;
  assign n23737 = n23736 ^ n20715;
  assign n23738 = n23737 ^ n23656;
  assign n23739 = ~n23657 & ~n23738;
  assign n23740 = n23739 ^ n20718;
  assign n23741 = n23740 ^ n23654;
  assign n23742 = ~n23655 & n23741;
  assign n23743 = n23742 ^ n20722;
  assign n23744 = n23743 ^ n23652;
  assign n23745 = n23653 & n23744;
  assign n23746 = n23745 ^ n20707;
  assign n23747 = n23746 ^ n23650;
  assign n23748 = ~n23651 & ~n23747;
  assign n23749 = n23748 ^ n20772;
  assign n23750 = n23749 ^ n20818;
  assign n23760 = n23759 ^ n23750;
  assign n23761 = n23737 ^ n23657;
  assign n23762 = n23731 ^ n21383;
  assign n23763 = n23762 ^ n23660;
  assign n23764 = n23717 ^ n23668;
  assign n23765 = n23709 ^ n23670;
  assign n23766 = n23696 ^ n23672;
  assign n23767 = n23693 ^ n20866;
  assign n23768 = n23685 ^ n23676;
  assign n23769 = n23682 ^ n20874;
  assign n23349 = n23348 ^ n20852;
  assign n23359 = n23358 ^ n23349;
  assign n23360 = n23345 ^ n23313;
  assign n23372 = ~n23370 & n23371;
  assign n23373 = n23342 ^ n23315;
  assign n23374 = ~n23372 & n23373;
  assign n23375 = n23360 & ~n23374;
  assign n23429 = n23359 & n23375;
  assign n23444 = n23443 ^ n20330;
  assign n23454 = n23429 & n23444;
  assign n23458 = n23457 ^ n20877;
  assign n23467 = n23466 ^ n23458;
  assign n23770 = ~n23454 & ~n23467;
  assign n23771 = ~n23769 & ~n23770;
  assign n23772 = n23768 & ~n23771;
  assign n23773 = n23688 ^ n23674;
  assign n23774 = ~n23772 & n23773;
  assign n23775 = ~n23767 & n23774;
  assign n23776 = n23766 & n23775;
  assign n23777 = n23701 ^ n20975;
  assign n23778 = n23776 & n23777;
  assign n23779 = n23706 ^ n21070;
  assign n23780 = ~n23778 & ~n23779;
  assign n23781 = n23765 & n23780;
  assign n23782 = n23714 ^ n21249;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = n23764 & n23783;
  assign n23785 = n23722 ^ n21292;
  assign n23786 = ~n23784 & ~n23785;
  assign n23787 = n23725 ^ n23665;
  assign n23788 = ~n23786 & n23787;
  assign n23789 = n23728 ^ n23663;
  assign n23790 = n23788 & ~n23789;
  assign n23791 = ~n23763 & ~n23790;
  assign n23792 = n23734 ^ n23659;
  assign n23793 = ~n23791 & n23792;
  assign n23794 = ~n23761 & n23793;
  assign n23795 = n23740 ^ n23655;
  assign n23796 = n23794 & n23795;
  assign n23797 = n23743 ^ n23653;
  assign n23798 = ~n23796 & n23797;
  assign n23799 = n23746 ^ n23651;
  assign n23800 = ~n23798 & ~n23799;
  assign n23945 = n23760 & n23800;
  assign n23940 = n22685 ^ n20857;
  assign n23941 = n23940 ^ n21675;
  assign n23937 = n23206 ^ n1336;
  assign n23938 = n23937 ^ n23046;
  assign n23934 = n23758 ^ n23755;
  assign n23935 = ~n23756 & ~n23934;
  assign n23936 = n23935 ^ n23758;
  assign n23939 = n23938 ^ n23936;
  assign n23942 = n23941 ^ n23939;
  assign n23943 = n23942 ^ n20839;
  assign n23930 = n23759 ^ n20818;
  assign n23931 = n23759 ^ n23749;
  assign n23932 = ~n23930 & n23931;
  assign n23933 = n23932 ^ n20818;
  assign n23944 = n23943 ^ n23933;
  assign n23946 = n23945 ^ n23944;
  assign n23801 = n23800 ^ n23760;
  assign n23802 = n23801 ^ n2480;
  assign n23803 = n23799 ^ n23798;
  assign n2495 = n2484 ^ n2417;
  assign n2496 = n2495 ^ n2401;
  assign n2497 = n2496 ^ n2476;
  assign n23804 = n23803 ^ n2497;
  assign n23805 = n23797 ^ n23796;
  assign n23806 = n23805 ^ n2396;
  assign n23915 = n23795 ^ n23794;
  assign n23808 = n2286 ^ n1344;
  assign n23809 = n23808 ^ n1298;
  assign n23810 = n23809 ^ n2376;
  assign n23807 = n23793 ^ n23761;
  assign n23811 = n23810 ^ n23807;
  assign n23812 = n23792 ^ n23791;
  assign n1286 = n1243 ^ n1186;
  assign n1287 = n1286 ^ n1280;
  assign n1288 = n1287 ^ n1202;
  assign n23813 = n23812 ^ n1288;
  assign n23814 = n23790 ^ n23763;
  assign n23815 = n23814 ^ n1273;
  assign n23816 = n23787 ^ n23786;
  assign n23817 = n23816 ^ n904;
  assign n23818 = n23785 ^ n23784;
  assign n23822 = n23821 ^ n23818;
  assign n23823 = n23783 ^ n23764;
  assign n23824 = n23823 ^ n768;
  assign n23825 = n23782 ^ n23781;
  assign n701 = n679 ^ n568;
  assign n702 = n701 ^ n698;
  assign n706 = n705 ^ n702;
  assign n23826 = n23825 ^ n706;
  assign n23827 = n23780 ^ n23765;
  assign n683 = n670 ^ n562;
  assign n690 = n689 ^ n683;
  assign n694 = n693 ^ n690;
  assign n23828 = n23827 ^ n694;
  assign n23829 = n23779 ^ n23778;
  assign n23833 = n23832 ^ n23829;
  assign n23834 = n23777 ^ n23776;
  assign n23838 = n23837 ^ n23834;
  assign n23872 = n23775 ^ n23766;
  assign n23839 = n23774 ^ n23767;
  assign n23843 = n23842 ^ n23839;
  assign n23861 = n23773 ^ n23772;
  assign n23844 = n23771 ^ n23768;
  assign n23848 = n23847 ^ n23844;
  assign n23849 = n23770 ^ n23769;
  assign n23850 = n23849 ^ n2183;
  assign n23468 = n23467 ^ n23454;
  assign n23851 = n23468 ^ n23452;
  assign n23445 = n23444 ^ n23429;
  assign n23376 = n23375 ^ n23359;
  assign n23377 = n23376 ^ n1846;
  assign n23378 = n23374 ^ n23360;
  assign n23379 = n23378 ^ n1834;
  assign n23380 = n23373 ^ n23372;
  assign n23381 = n23380 ^ n1736;
  assign n23417 = n23416 ^ n23382;
  assign n23418 = n23383 & ~n23417;
  assign n23419 = n23418 ^ n1724;
  assign n23420 = n23419 ^ n23380;
  assign n23421 = ~n23381 & n23420;
  assign n23422 = n23421 ^ n1736;
  assign n23423 = n23422 ^ n23378;
  assign n23424 = n23379 & ~n23423;
  assign n23425 = n23424 ^ n1834;
  assign n23426 = n23425 ^ n23376;
  assign n23427 = ~n23377 & n23426;
  assign n23428 = n23427 ^ n1846;
  assign n23446 = n23445 ^ n23428;
  assign n23447 = n23445 ^ n1995;
  assign n23448 = n23446 & ~n23447;
  assign n23449 = n23448 ^ n1995;
  assign n23852 = n23468 ^ n23449;
  assign n23853 = n23851 & ~n23852;
  assign n23854 = n23853 ^ n23452;
  assign n23855 = n23854 ^ n23849;
  assign n23856 = ~n23850 & n23855;
  assign n23857 = n23856 ^ n2183;
  assign n23858 = n23857 ^ n23844;
  assign n23859 = ~n23848 & n23858;
  assign n23860 = n23859 ^ n23847;
  assign n23862 = n23861 ^ n23860;
  assign n23866 = n23865 ^ n23861;
  assign n23867 = ~n23862 & n23866;
  assign n23868 = n23867 ^ n23865;
  assign n23869 = n23868 ^ n23839;
  assign n23870 = n23843 & ~n23869;
  assign n23871 = n23870 ^ n23842;
  assign n23873 = n23872 ^ n23871;
  assign n23877 = n23876 ^ n23872;
  assign n23878 = n23873 & ~n23877;
  assign n23879 = n23878 ^ n23876;
  assign n23880 = n23879 ^ n23834;
  assign n23881 = ~n23838 & n23880;
  assign n23882 = n23881 ^ n23837;
  assign n23883 = n23882 ^ n23829;
  assign n23884 = n23833 & ~n23883;
  assign n23885 = n23884 ^ n23832;
  assign n23886 = n23885 ^ n23827;
  assign n23887 = n23828 & ~n23886;
  assign n23888 = n23887 ^ n694;
  assign n23889 = n23888 ^ n23825;
  assign n23890 = ~n23826 & n23889;
  assign n23891 = n23890 ^ n706;
  assign n23892 = n23891 ^ n23823;
  assign n23893 = ~n23824 & n23892;
  assign n23894 = n23893 ^ n768;
  assign n23895 = n23894 ^ n23818;
  assign n23896 = n23822 & ~n23895;
  assign n23897 = n23896 ^ n23821;
  assign n23898 = n23897 ^ n23816;
  assign n23899 = n23817 & ~n23898;
  assign n23900 = n23899 ^ n904;
  assign n23901 = n23900 ^ n1264;
  assign n23902 = n23789 ^ n23788;
  assign n23903 = n23902 ^ n23900;
  assign n23904 = n23901 & ~n23903;
  assign n23905 = n23904 ^ n1264;
  assign n23906 = n23905 ^ n23814;
  assign n23907 = n23815 & ~n23906;
  assign n23908 = n23907 ^ n1273;
  assign n23909 = n23908 ^ n23812;
  assign n23910 = n23813 & ~n23909;
  assign n23911 = n23910 ^ n1288;
  assign n23912 = n23911 ^ n23807;
  assign n23913 = n23811 & ~n23912;
  assign n23914 = n23913 ^ n23810;
  assign n23916 = n23915 ^ n23914;
  assign n2373 = n2294 ^ n1359;
  assign n2380 = n2379 ^ n2373;
  assign n2384 = n2383 ^ n2380;
  assign n23917 = n23915 ^ n2384;
  assign n23918 = n23916 & ~n23917;
  assign n23919 = n23918 ^ n2384;
  assign n23920 = n23919 ^ n23805;
  assign n23921 = ~n23806 & n23920;
  assign n23922 = n23921 ^ n2396;
  assign n23923 = n23922 ^ n23803;
  assign n23924 = ~n23804 & n23923;
  assign n23925 = n23924 ^ n2497;
  assign n23926 = n23925 ^ n23801;
  assign n23927 = ~n23802 & n23926;
  assign n23928 = n23927 ^ n2480;
  assign n2643 = n2639 ^ n2568;
  assign n2647 = n2646 ^ n2643;
  assign n2648 = n2647 ^ n1497;
  assign n23929 = n23928 ^ n2648;
  assign n23947 = n23946 ^ n23929;
  assign n23950 = n23949 ^ n23947;
  assign n23969 = n23925 ^ n23802;
  assign n23962 = n23922 ^ n23804;
  assign n23953 = n22538 ^ n21674;
  assign n23954 = n23953 ^ n22598;
  assign n23955 = n23916 ^ n2384;
  assign n23956 = ~n23954 & ~n23955;
  assign n23951 = n23300 ^ n21670;
  assign n23952 = n23951 ^ n22540;
  assign n23957 = n23956 ^ n23952;
  assign n23958 = n23919 ^ n23806;
  assign n23959 = n23958 ^ n23952;
  assign n23960 = n23957 & n23959;
  assign n23961 = n23960 ^ n23956;
  assign n23963 = n23962 ^ n23961;
  assign n23964 = n23308 ^ n22591;
  assign n23965 = n23964 ^ n22057;
  assign n23966 = n23965 ^ n23962;
  assign n23967 = n23963 & ~n23966;
  assign n23968 = n23967 ^ n23965;
  assign n23970 = n23969 ^ n23968;
  assign n23971 = n23354 ^ n21668;
  assign n23972 = n23971 ^ n22729;
  assign n23973 = n23972 ^ n23969;
  assign n23974 = n23970 & ~n23973;
  assign n23975 = n23974 ^ n23972;
  assign n23976 = n23975 ^ n23947;
  assign n23977 = n23950 & ~n23976;
  assign n23978 = n23977 ^ n23949;
  assign n23979 = n23978 ^ n23517;
  assign n23980 = n23520 & n23979;
  assign n23981 = n23980 ^ n23519;
  assign n23982 = n23981 ^ n23512;
  assign n23983 = ~n23516 & n23982;
  assign n23984 = n23983 ^ n23515;
  assign n23985 = n23984 ^ n23510;
  assign n23986 = n23511 & ~n23985;
  assign n23987 = n23986 ^ n23507;
  assign n23988 = n23987 ^ n23504;
  assign n23989 = ~n23506 & ~n23988;
  assign n23990 = n23989 ^ n23505;
  assign n23991 = n23990 ^ n23497;
  assign n23992 = ~n23501 & ~n23991;
  assign n23993 = n23992 ^ n23500;
  assign n23994 = n23993 ^ n23492;
  assign n23995 = ~n23496 & n23994;
  assign n23996 = n23995 ^ n23495;
  assign n23487 = n22567 ^ n22100;
  assign n23490 = n23489 ^ n23487;
  assign n23486 = n23419 ^ n23381;
  assign n23491 = n23490 ^ n23486;
  assign n24030 = n23996 ^ n23491;
  assign n24031 = n24030 ^ n21656;
  assign n24032 = n23993 ^ n23495;
  assign n24033 = n24032 ^ n23492;
  assign n24034 = n24033 ^ n21661;
  assign n24035 = n23990 ^ n23501;
  assign n24036 = n24035 ^ n21701;
  assign n24037 = n23987 ^ n23506;
  assign n24038 = n24037 ^ n21666;
  assign n24072 = n23984 ^ n23511;
  assign n24061 = n23978 ^ n23520;
  assign n24039 = n23975 ^ n23950;
  assign n24040 = n24039 ^ n20849;
  assign n24041 = n23972 ^ n23970;
  assign n24042 = n24041 ^ n20850;
  assign n24043 = n23965 ^ n23963;
  assign n24044 = n24043 ^ n21420;
  assign n24045 = n23955 ^ n23954;
  assign n24046 = n20856 & n24045;
  assign n24047 = n24046 ^ n20855;
  assign n24048 = n23958 ^ n23957;
  assign n24049 = n24048 ^ n24046;
  assign n24050 = ~n24047 & n24049;
  assign n24051 = n24050 ^ n20855;
  assign n24052 = n24051 ^ n24043;
  assign n24053 = n24044 & ~n24052;
  assign n24054 = n24053 ^ n21420;
  assign n24055 = n24054 ^ n24041;
  assign n24056 = ~n24042 & ~n24055;
  assign n24057 = n24056 ^ n20850;
  assign n24058 = n24057 ^ n24039;
  assign n24059 = ~n24040 & ~n24058;
  assign n24060 = n24059 ^ n20849;
  assign n24062 = n24061 ^ n24060;
  assign n24063 = n24060 ^ n21491;
  assign n24064 = n24062 & ~n24063;
  assign n24065 = n24064 ^ n21491;
  assign n24066 = n24065 ^ n21527;
  assign n24067 = n23981 ^ n23515;
  assign n24068 = n24067 ^ n23512;
  assign n24069 = n24068 ^ n24065;
  assign n24070 = n24066 & ~n24069;
  assign n24071 = n24070 ^ n21527;
  assign n24073 = n24072 ^ n24071;
  assign n24074 = n24072 ^ n21631;
  assign n24075 = n24073 & n24074;
  assign n24076 = n24075 ^ n21631;
  assign n24077 = n24076 ^ n24037;
  assign n24078 = n24038 & n24077;
  assign n24079 = n24078 ^ n21666;
  assign n24080 = n24079 ^ n24035;
  assign n24081 = n24036 & n24080;
  assign n24082 = n24081 ^ n21701;
  assign n24083 = n24082 ^ n24033;
  assign n24084 = ~n24034 & n24083;
  assign n24085 = n24084 ^ n21661;
  assign n24086 = n24085 ^ n24030;
  assign n24087 = ~n24031 & ~n24086;
  assign n24088 = n24087 ^ n21656;
  assign n24146 = n24088 ^ n21694;
  assign n23997 = n23996 ^ n23490;
  assign n23998 = n23491 & ~n23997;
  assign n23999 = n23998 ^ n23486;
  assign n23483 = n23482 ^ n21644;
  assign n23484 = n23483 ^ n22768;
  assign n23480 = n23422 ^ n1834;
  assign n23481 = n23480 ^ n23378;
  assign n23485 = n23484 ^ n23481;
  assign n24028 = n23999 ^ n23485;
  assign n24147 = n24146 ^ n24028;
  assign n24119 = n24079 ^ n21701;
  assign n24120 = n24119 ^ n24035;
  assign n24121 = n24076 ^ n24038;
  assign n24122 = n24057 ^ n24040;
  assign n24123 = n24054 ^ n20850;
  assign n24124 = n24123 ^ n24041;
  assign n24125 = n24051 ^ n24044;
  assign n24126 = n24045 ^ n20856;
  assign n24127 = n24048 ^ n24047;
  assign n24128 = n24126 & n24127;
  assign n24129 = ~n24125 & n24128;
  assign n24130 = n24124 & n24129;
  assign n24131 = ~n24122 & n24130;
  assign n24132 = n24062 ^ n21491;
  assign n24133 = ~n24131 & n24132;
  assign n24134 = n24068 ^ n21527;
  assign n24135 = n24134 ^ n24065;
  assign n24136 = ~n24133 & n24135;
  assign n24137 = n24073 ^ n21631;
  assign n24138 = ~n24136 & ~n24137;
  assign n24139 = n24121 & n24138;
  assign n24140 = ~n24120 & n24139;
  assign n24141 = n24082 ^ n21661;
  assign n24142 = n24141 ^ n24033;
  assign n24143 = ~n24140 & n24142;
  assign n24144 = n24085 ^ n24031;
  assign n24145 = ~n24143 & ~n24144;
  assign n24245 = n24147 ^ n24145;
  assign n24171 = n24144 ^ n24143;
  assign n24175 = n24174 ^ n24171;
  assign n24176 = n24142 ^ n24140;
  assign n24177 = n24176 ^ n2102;
  assign n24178 = n24139 ^ n24120;
  assign n24179 = n24178 ^ n1974;
  assign n24231 = n24138 ^ n24121;
  assign n24226 = n24137 ^ n24136;
  assign n24183 = n24135 ^ n24133;
  assign n24180 = n22412 ^ n1789;
  assign n24181 = n24180 ^ n1643;
  assign n24182 = n24181 ^ n1939;
  assign n24184 = n24183 ^ n24182;
  assign n24185 = n24132 ^ n24131;
  assign n24189 = n24188 ^ n24185;
  assign n24190 = n24130 ^ n24122;
  assign n24191 = n24190 ^ n1460;
  assign n24192 = n24129 ^ n24124;
  assign n24196 = n24195 ^ n24192;
  assign n24209 = n24128 ^ n24125;
  assign n24203 = ~n24126 & n24202;
  assign n24197 = n22392 ^ n1466;
  assign n24198 = n24197 ^ n18851;
  assign n24199 = n24198 ^ n1490;
  assign n24204 = n24203 ^ n24199;
  assign n24205 = n24127 ^ n24126;
  assign n24206 = n24205 ^ n24203;
  assign n24207 = n24204 & ~n24206;
  assign n24208 = n24207 ^ n24199;
  assign n24210 = n24209 ^ n24208;
  assign n24211 = n24208 ^ n1529;
  assign n24212 = n24210 & n24211;
  assign n24213 = n24212 ^ n1529;
  assign n24214 = n24213 ^ n24192;
  assign n24215 = n24196 & ~n24214;
  assign n24216 = n24215 ^ n24195;
  assign n24217 = n24216 ^ n24190;
  assign n24218 = ~n24191 & n24217;
  assign n24219 = n24218 ^ n1460;
  assign n24220 = n24219 ^ n24185;
  assign n24221 = n24189 & ~n24220;
  assign n24222 = n24221 ^ n24188;
  assign n24223 = n24222 ^ n24183;
  assign n24224 = ~n24184 & n24223;
  assign n24225 = n24224 ^ n24182;
  assign n24227 = n24226 ^ n24225;
  assign n24228 = n24226 ^ n1944;
  assign n24229 = n24227 & ~n24228;
  assign n24230 = n24229 ^ n1944;
  assign n24232 = n24231 ^ n24230;
  assign n24233 = n24231 ^ n1956;
  assign n24234 = n24232 & ~n24233;
  assign n24235 = n24234 ^ n1956;
  assign n24236 = n24235 ^ n24178;
  assign n24237 = n24179 & ~n24236;
  assign n24238 = n24237 ^ n1974;
  assign n24239 = n24238 ^ n24176;
  assign n24240 = ~n24177 & n24239;
  assign n24241 = n24240 ^ n2102;
  assign n24242 = n24241 ^ n24171;
  assign n24243 = ~n24175 & n24242;
  assign n24244 = n24243 ^ n24174;
  assign n24246 = n24245 ^ n24244;
  assign n24707 = n24249 ^ n24246;
  assign n24700 = n24241 ^ n24175;
  assign n24323 = n23876 ^ n23871;
  assign n24324 = n24323 ^ n23872;
  assign n24325 = n24324 ^ n23550;
  assign n24326 = n24325 ^ n22555;
  assign n24322 = n24238 ^ n24177;
  assign n24327 = n24326 ^ n24322;
  assign n24331 = n23470 ^ n22563;
  assign n24282 = n23865 ^ n23862;
  assign n24332 = n24331 ^ n24282;
  assign n24330 = n24232 ^ n1956;
  assign n24333 = n24332 ^ n24330;
  assign n24336 = n24227 ^ n1944;
  assign n24110 = n23857 ^ n23847;
  assign n24111 = n24110 ^ n23844;
  assign n24334 = n24111 ^ n22768;
  assign n24335 = n24334 ^ n23560;
  assign n24337 = n24336 ^ n24335;
  assign n24340 = n24222 ^ n24184;
  assign n24338 = n23475 ^ n22567;
  assign n24018 = n23854 ^ n23850;
  assign n24339 = n24338 ^ n24018;
  assign n24341 = n24340 ^ n24339;
  assign n24674 = n24219 ^ n24188;
  assign n24675 = n24674 ^ n24185;
  assign n24343 = n23489 ^ n22577;
  assign n23474 = n23446 ^ n1995;
  assign n24344 = n24343 ^ n23474;
  assign n24342 = n24216 ^ n24191;
  assign n24345 = n24344 ^ n24342;
  assign n24347 = n23493 ^ n22581;
  assign n23478 = n23425 ^ n23377;
  assign n24348 = n24347 ^ n23478;
  assign n24346 = n24213 ^ n24196;
  assign n24349 = n24348 ^ n24346;
  assign n24352 = n23486 ^ n22746;
  assign n24353 = n24352 ^ n23502;
  assign n24351 = n24205 ^ n24204;
  assign n24354 = n24353 ^ n24351;
  assign n24356 = n23508 ^ n23492;
  assign n24357 = n24356 ^ n22589;
  assign n24355 = n24202 ^ n24126;
  assign n24358 = n24357 ^ n24355;
  assign n24499 = n23241 ^ n22606;
  assign n24500 = n24499 ^ n21679;
  assign n24496 = n23908 ^ n1288;
  assign n24497 = n24496 ^ n23812;
  assign n24432 = n23905 ^ n23815;
  assign n24430 = n23243 ^ n22685;
  assign n24431 = n24430 ^ n22035;
  assign n24433 = n24432 ^ n24431;
  assign n24361 = n22691 ^ n22012;
  assign n24362 = n24361 ^ n23254;
  assign n24293 = n23902 ^ n1264;
  assign n24294 = n24293 ^ n23900;
  assign n24363 = n24362 ^ n24294;
  assign n24364 = n23938 ^ n22701;
  assign n24365 = n24364 ^ n21960;
  assign n24304 = n23894 ^ n23822;
  assign n24366 = n24365 ^ n24304;
  assign n24369 = n23891 ^ n23824;
  assign n24367 = n23755 ^ n21938;
  assign n24368 = n24367 ^ n22530;
  assign n24370 = n24369 ^ n24368;
  assign n24373 = n23882 ^ n23832;
  assign n24374 = n24373 ^ n23829;
  assign n24371 = n23029 ^ n22551;
  assign n24372 = n24371 ^ n23526;
  assign n24375 = n24374 ^ n24372;
  assign n24378 = n23879 ^ n23838;
  assign n24376 = n22952 ^ n22614;
  assign n24377 = n24376 ^ n23530;
  assign n24379 = n24378 ^ n24377;
  assign n24382 = n23539 ^ n22542;
  assign n24383 = n24382 ^ n22337;
  assign n24380 = n23868 ^ n23842;
  assign n24381 = n24380 ^ n23839;
  assign n24384 = n24383 ^ n24381;
  assign n24280 = n23545 ^ n22323;
  assign n24281 = n24280 ^ n22548;
  assign n24283 = n24282 ^ n24281;
  assign n24108 = n23550 ^ n22549;
  assign n24109 = n24108 ^ n22309;
  assign n24112 = n24111 ^ n24109;
  assign n24015 = n23554 ^ n22554;
  assign n24016 = n24015 ^ n22294;
  assign n24104 = n24018 ^ n24016;
  assign n23471 = n23470 ^ n22279;
  assign n23472 = n23471 ^ n22555;
  assign n23453 = n23452 ^ n23449;
  assign n23469 = n23468 ^ n23453;
  assign n23473 = n23472 ^ n23469;
  assign n23476 = n23475 ^ n22113;
  assign n23477 = n23476 ^ n22563;
  assign n23479 = n23478 ^ n23477;
  assign n24000 = n23999 ^ n23481;
  assign n24001 = n23485 & n24000;
  assign n24002 = n24001 ^ n23484;
  assign n24003 = n24002 ^ n23478;
  assign n24004 = n23479 & n24003;
  assign n24005 = n24004 ^ n23477;
  assign n24006 = n24005 ^ n23474;
  assign n24007 = n23560 ^ n22559;
  assign n24008 = n24007 ^ n22225;
  assign n24009 = n24008 ^ n23474;
  assign n24010 = ~n24006 & ~n24009;
  assign n24011 = n24010 ^ n24008;
  assign n24012 = n24011 ^ n23469;
  assign n24013 = ~n23473 & ~n24012;
  assign n24014 = n24013 ^ n23472;
  assign n24105 = n24018 ^ n24014;
  assign n24106 = ~n24104 & ~n24105;
  assign n24107 = n24106 ^ n24016;
  assign n24277 = n24111 ^ n24107;
  assign n24278 = n24112 & n24277;
  assign n24279 = n24278 ^ n24109;
  assign n24385 = n24282 ^ n24279;
  assign n24386 = ~n24283 & n24385;
  assign n24387 = n24386 ^ n24281;
  assign n24388 = n24387 ^ n24381;
  assign n24389 = ~n24384 & n24388;
  assign n24390 = n24389 ^ n24383;
  assign n24391 = n24390 ^ n24324;
  assign n24392 = n23534 ^ n22802;
  assign n24393 = n24392 ^ n22518;
  assign n24394 = n24393 ^ n24324;
  assign n24395 = ~n24391 & ~n24394;
  assign n24396 = n24395 ^ n24393;
  assign n24397 = n24396 ^ n24378;
  assign n24398 = n24379 & n24397;
  assign n24399 = n24398 ^ n24377;
  assign n24400 = n24399 ^ n24374;
  assign n24401 = n24375 & n24400;
  assign n24402 = n24401 ^ n24372;
  assign n24317 = n23885 ^ n694;
  assign n24318 = n24317 ^ n23827;
  assign n24403 = n24402 ^ n24318;
  assign n24404 = n23226 ^ n22645;
  assign n24405 = n24404 ^ n23522;
  assign n24406 = n24405 ^ n24318;
  assign n24407 = ~n24403 & ~n24406;
  assign n24408 = n24407 ^ n24405;
  assign n24311 = n23888 ^ n23826;
  assign n24409 = n24408 ^ n24311;
  assign n24410 = n23649 ^ n22544;
  assign n24411 = n24410 ^ n23275;
  assign n24412 = n24411 ^ n24311;
  assign n24413 = ~n24409 & n24412;
  assign n24414 = n24413 ^ n24411;
  assign n24415 = n24414 ^ n24369;
  assign n24416 = n24370 & ~n24415;
  assign n24417 = n24416 ^ n24368;
  assign n24418 = n24417 ^ n24304;
  assign n24419 = n24366 & n24418;
  assign n24420 = n24419 ^ n24365;
  assign n24298 = n23897 ^ n23817;
  assign n24421 = n24420 ^ n24298;
  assign n24422 = n23249 ^ n22693;
  assign n24423 = n24422 ^ n21983;
  assign n24424 = n24423 ^ n24298;
  assign n24425 = ~n24421 & ~n24424;
  assign n24426 = n24425 ^ n24423;
  assign n24427 = n24426 ^ n24294;
  assign n24428 = n24363 & n24427;
  assign n24429 = n24428 ^ n24362;
  assign n24493 = n24431 ^ n24429;
  assign n24494 = n24433 & ~n24493;
  assign n24495 = n24494 ^ n24432;
  assign n24498 = n24497 ^ n24495;
  assign n24501 = n24500 ^ n24498;
  assign n24502 = n24501 ^ n21395;
  assign n24434 = n24433 ^ n24429;
  assign n24435 = n24434 ^ n21388;
  assign n24436 = n24426 ^ n24363;
  assign n24437 = n24436 ^ n21358;
  assign n24438 = n24423 ^ n24421;
  assign n24439 = n24438 ^ n21329;
  assign n24440 = n24417 ^ n24366;
  assign n24441 = n24440 ^ n21303;
  assign n24442 = n24414 ^ n24370;
  assign n24443 = n24442 ^ n21279;
  assign n24444 = n24411 ^ n24409;
  assign n24445 = n24444 ^ n22026;
  assign n24446 = n24405 ^ n24403;
  assign n24447 = n24446 ^ n22001;
  assign n24466 = n24399 ^ n24372;
  assign n24467 = n24466 ^ n24374;
  assign n24461 = n24396 ^ n24379;
  assign n24456 = n24393 ^ n24391;
  assign n24448 = n24387 ^ n24384;
  assign n24449 = n24448 ^ n21911;
  assign n24284 = n24283 ^ n24279;
  assign n24113 = n24112 ^ n24107;
  assign n24017 = n24016 ^ n24014;
  assign n24019 = n24018 ^ n24017;
  assign n24020 = n24019 ^ n21741;
  assign n24021 = n24011 ^ n23473;
  assign n24022 = n24021 ^ n21646;
  assign n24023 = n24008 ^ n24006;
  assign n24024 = n24023 ^ n21692;
  assign n24025 = n24002 ^ n23477;
  assign n24026 = n24025 ^ n23478;
  assign n24027 = n24026 ^ n21652;
  assign n24029 = n24028 ^ n21694;
  assign n24089 = n24088 ^ n24028;
  assign n24090 = n24029 & n24089;
  assign n24091 = n24090 ^ n21694;
  assign n24092 = n24091 ^ n24026;
  assign n24093 = n24027 & n24092;
  assign n24094 = n24093 ^ n21652;
  assign n24095 = n24094 ^ n24023;
  assign n24096 = n24024 & ~n24095;
  assign n24097 = n24096 ^ n21692;
  assign n24098 = n24097 ^ n24021;
  assign n24099 = n24022 & n24098;
  assign n24100 = n24099 ^ n21646;
  assign n24101 = n24100 ^ n24019;
  assign n24102 = ~n24020 & n24101;
  assign n24103 = n24102 ^ n21741;
  assign n24114 = n24113 ^ n24103;
  assign n24274 = n24113 ^ n21748;
  assign n24275 = n24114 & ~n24274;
  assign n24276 = n24275 ^ n21748;
  assign n24285 = n24284 ^ n24276;
  assign n24450 = n24284 ^ n21808;
  assign n24451 = n24285 & n24450;
  assign n24452 = n24451 ^ n21808;
  assign n24453 = n24452 ^ n24448;
  assign n24454 = ~n24449 & ~n24453;
  assign n24455 = n24454 ^ n21911;
  assign n24457 = n24456 ^ n24455;
  assign n24458 = n24456 ^ n21931;
  assign n24459 = n24457 & n24458;
  assign n24460 = n24459 ^ n21931;
  assign n24462 = n24461 ^ n24460;
  assign n24463 = n24461 ^ n21949;
  assign n24464 = ~n24462 & ~n24463;
  assign n24465 = n24464 ^ n21949;
  assign n24468 = n24467 ^ n24465;
  assign n24469 = n24467 ^ n21973;
  assign n24470 = ~n24468 & n24469;
  assign n24471 = n24470 ^ n21973;
  assign n24472 = n24471 ^ n24446;
  assign n24473 = ~n24447 & ~n24472;
  assign n24474 = n24473 ^ n22001;
  assign n24475 = n24474 ^ n24444;
  assign n24476 = n24445 & n24475;
  assign n24477 = n24476 ^ n22026;
  assign n24478 = n24477 ^ n24442;
  assign n24479 = ~n24443 & ~n24478;
  assign n24480 = n24479 ^ n21279;
  assign n24481 = n24480 ^ n24440;
  assign n24482 = ~n24441 & n24481;
  assign n24483 = n24482 ^ n21303;
  assign n24484 = n24483 ^ n24438;
  assign n24485 = ~n24439 & n24484;
  assign n24486 = n24485 ^ n21329;
  assign n24487 = n24486 ^ n24436;
  assign n24488 = n24437 & n24487;
  assign n24489 = n24488 ^ n21358;
  assign n24490 = n24489 ^ n24434;
  assign n24491 = n24435 & n24490;
  assign n24492 = n24491 ^ n21388;
  assign n24503 = n24502 ^ n24492;
  assign n24504 = n24489 ^ n21388;
  assign n24505 = n24504 ^ n24434;
  assign n24506 = n24483 ^ n21329;
  assign n24507 = n24506 ^ n24438;
  assign n24508 = n24480 ^ n21303;
  assign n24509 = n24508 ^ n24440;
  assign n24510 = n24471 ^ n24447;
  assign n24511 = n24468 ^ n21973;
  assign n24512 = n24462 ^ n21949;
  assign n24513 = n24457 ^ n21931;
  assign n24115 = n24114 ^ n21748;
  assign n24116 = n24100 ^ n24020;
  assign n24117 = n24094 ^ n24024;
  assign n24118 = n24091 ^ n24027;
  assign n24148 = ~n24145 & n24147;
  assign n24149 = n24118 & ~n24148;
  assign n24150 = ~n24117 & n24149;
  assign n24151 = n24097 ^ n24022;
  assign n24152 = n24150 & ~n24151;
  assign n24153 = ~n24116 & n24152;
  assign n24273 = n24115 & ~n24153;
  assign n24286 = n24285 ^ n21808;
  assign n24514 = n24273 & ~n24286;
  assign n24515 = n24452 ^ n21911;
  assign n24516 = n24515 ^ n24448;
  assign n24517 = ~n24514 & n24516;
  assign n24518 = n24513 & n24517;
  assign n24519 = ~n24512 & ~n24518;
  assign n24520 = n24511 & ~n24519;
  assign n24521 = ~n24510 & n24520;
  assign n24522 = n24474 ^ n24445;
  assign n24523 = ~n24521 & n24522;
  assign n24524 = n24477 ^ n24443;
  assign n24525 = ~n24523 & ~n24524;
  assign n24526 = n24509 & n24525;
  assign n24527 = n24507 & n24526;
  assign n24528 = n24486 ^ n24437;
  assign n24529 = ~n24527 & n24528;
  assign n24530 = n24505 & ~n24529;
  assign n24621 = n24503 & n24530;
  assign n24615 = n23911 ^ n23810;
  assign n24616 = n24615 ^ n23807;
  assign n24613 = n23287 ^ n22602;
  assign n24614 = n24613 ^ n21675;
  assign n24617 = n24616 ^ n24614;
  assign n24610 = n24500 ^ n24497;
  assign n24611 = ~n24498 & ~n24610;
  assign n24612 = n24611 ^ n24500;
  assign n24618 = n24617 ^ n24612;
  assign n24607 = n24501 ^ n24492;
  assign n24608 = ~n24502 & n24607;
  assign n24609 = n24608 ^ n21395;
  assign n24619 = n24618 ^ n24609;
  assign n24620 = n24619 ^ n20857;
  assign n24622 = n24621 ^ n24620;
  assign n24531 = n24530 ^ n24503;
  assign n24532 = n24531 ^ n2590;
  assign n24533 = n24529 ^ n24505;
  assign n2596 = n2511 ^ n2445;
  assign n2597 = n2596 ^ n2595;
  assign n2598 = n2597 ^ n2426;
  assign n24534 = n24533 ^ n2598;
  assign n24536 = n22528 ^ n2437;
  assign n24537 = n24536 ^ n2318;
  assign n24538 = n24537 ^ n1538;
  assign n24535 = n24528 ^ n24527;
  assign n24539 = n24538 ^ n24535;
  assign n24541 = n22347 ^ n2452;
  assign n24542 = n24541 ^ n19442;
  assign n24543 = n24542 ^ n2309;
  assign n24540 = n24526 ^ n24507;
  assign n24544 = n24543 ^ n24540;
  assign n24545 = n24525 ^ n24509;
  assign n1305 = n1304 ^ n1214;
  assign n1312 = n1311 ^ n1305;
  assign n1316 = n1315 ^ n1312;
  assign n24546 = n24545 ^ n1316;
  assign n24547 = n24524 ^ n24523;
  assign n24551 = n24550 ^ n24547;
  assign n24552 = n24522 ^ n24521;
  assign n24553 = n24552 ^ n1125;
  assign n24580 = n24520 ^ n24510;
  assign n24554 = n24519 ^ n24511;
  assign n24555 = n24554 ^ n964;
  assign n24556 = n24518 ^ n24512;
  assign n24557 = n24556 ^ n860;
  assign n24558 = n24517 ^ n24513;
  assign n837 = n788 ^ n737;
  assign n844 = n843 ^ n837;
  assign n848 = n847 ^ n844;
  assign n24559 = n24558 ^ n848;
  assign n24560 = n24516 ^ n24514;
  assign n24564 = n24563 ^ n24560;
  assign n24287 = n24286 ^ n24273;
  assign n24291 = n24290 ^ n24287;
  assign n24154 = n24153 ^ n24115;
  assign n24158 = n24157 ^ n24154;
  assign n24262 = n24152 ^ n24116;
  assign n24159 = n24151 ^ n24150;
  assign n24160 = n24159 ^ n614;
  assign n24161 = n24149 ^ n24117;
  assign n24165 = n24164 ^ n24161;
  assign n24166 = n24148 ^ n24118;
  assign n24170 = n24169 ^ n24166;
  assign n24250 = n24249 ^ n24245;
  assign n24251 = n24246 & ~n24250;
  assign n24252 = n24251 ^ n24249;
  assign n24253 = n24252 ^ n24166;
  assign n24254 = n24170 & ~n24253;
  assign n24255 = n24254 ^ n24169;
  assign n24256 = n24255 ^ n24161;
  assign n24257 = n24165 & ~n24256;
  assign n24258 = n24257 ^ n24164;
  assign n24259 = n24258 ^ n24159;
  assign n24260 = n24160 & ~n24259;
  assign n24261 = n24260 ^ n614;
  assign n24263 = n24262 ^ n24261;
  assign n24264 = n22463 ^ n15587;
  assign n24265 = n24264 ^ n19321;
  assign n24266 = n24265 ^ n528;
  assign n24267 = n24266 ^ n24262;
  assign n24268 = ~n24263 & n24267;
  assign n24269 = n24268 ^ n24266;
  assign n24270 = n24269 ^ n24154;
  assign n24271 = ~n24158 & n24270;
  assign n24272 = n24271 ^ n24157;
  assign n24565 = n24287 ^ n24272;
  assign n24566 = ~n24291 & n24565;
  assign n24567 = n24566 ^ n24290;
  assign n24568 = n24567 ^ n24560;
  assign n24569 = n24564 & ~n24568;
  assign n24570 = n24569 ^ n24563;
  assign n24571 = n24570 ^ n24558;
  assign n24572 = ~n24559 & n24571;
  assign n24573 = n24572 ^ n848;
  assign n24574 = n24573 ^ n24556;
  assign n24575 = n24557 & ~n24574;
  assign n24576 = n24575 ^ n860;
  assign n24577 = n24576 ^ n24554;
  assign n24578 = n24555 & ~n24577;
  assign n24579 = n24578 ^ n964;
  assign n24581 = n24580 ^ n24579;
  assign n24582 = n24580 ^ n976;
  assign n24583 = ~n24581 & n24582;
  assign n24584 = n24583 ^ n976;
  assign n24585 = n24584 ^ n24552;
  assign n24586 = ~n24553 & n24585;
  assign n24587 = n24586 ^ n1125;
  assign n24588 = n24587 ^ n24547;
  assign n24589 = ~n24551 & n24588;
  assign n24590 = n24589 ^ n24550;
  assign n24591 = n24590 ^ n24545;
  assign n24592 = ~n24546 & n24591;
  assign n24593 = n24592 ^ n1316;
  assign n24594 = n24593 ^ n24543;
  assign n24595 = ~n24544 & ~n24594;
  assign n24596 = n24595 ^ n24540;
  assign n24597 = n24596 ^ n24535;
  assign n24598 = ~n24539 & ~n24597;
  assign n24599 = n24598 ^ n24538;
  assign n24600 = n24599 ^ n24533;
  assign n24601 = n24534 & ~n24600;
  assign n24602 = n24601 ^ n2598;
  assign n24603 = n24602 ^ n24531;
  assign n24604 = ~n24532 & n24603;
  assign n24605 = n24604 ^ n2590;
  assign n24606 = n24605 ^ n2617;
  assign n24623 = n24622 ^ n24606;
  assign n24359 = n23497 ^ n22736;
  assign n24360 = n24359 ^ n23513;
  assign n24624 = n24623 ^ n24360;
  assign n24627 = n24602 ^ n2590;
  assign n24628 = n24627 ^ n24531;
  assign n24625 = n23505 ^ n23465;
  assign n24626 = n24625 ^ n22729;
  assign n24629 = n24628 ^ n24626;
  assign n24632 = n23440 ^ n22591;
  assign n24633 = n24632 ^ n23507;
  assign n24630 = n24599 ^ n2598;
  assign n24631 = n24630 ^ n24533;
  assign n24634 = n24633 ^ n24631;
  assign n24637 = n24593 ^ n24544;
  assign n24638 = n23517 ^ n23308;
  assign n24639 = n24638 ^ n22598;
  assign n24640 = ~n24637 & ~n24639;
  assign n24635 = n23512 ^ n22540;
  assign n24636 = n24635 ^ n23354;
  assign n24641 = n24640 ^ n24636;
  assign n24642 = n24596 ^ n24538;
  assign n24643 = n24642 ^ n24535;
  assign n24644 = n24643 ^ n24636;
  assign n24645 = n24641 & ~n24644;
  assign n24646 = n24645 ^ n24640;
  assign n24647 = n24646 ^ n24631;
  assign n24648 = ~n24634 & ~n24647;
  assign n24649 = n24648 ^ n24633;
  assign n24650 = n24649 ^ n24628;
  assign n24651 = n24629 & ~n24650;
  assign n24652 = n24651 ^ n24626;
  assign n24653 = n24652 ^ n24360;
  assign n24654 = n24624 & n24653;
  assign n24655 = n24654 ^ n24623;
  assign n24656 = n24655 ^ n24357;
  assign n24657 = ~n24358 & ~n24656;
  assign n24658 = n24657 ^ n24355;
  assign n24659 = n24658 ^ n24351;
  assign n24660 = ~n24354 & n24659;
  assign n24661 = n24660 ^ n24353;
  assign n24350 = n24210 ^ n1529;
  assign n24662 = n24661 ^ n24350;
  assign n24663 = n23481 ^ n22585;
  assign n24664 = n24663 ^ n23498;
  assign n24665 = n24664 ^ n24350;
  assign n24666 = ~n24662 & ~n24665;
  assign n24667 = n24666 ^ n24664;
  assign n24668 = n24667 ^ n24346;
  assign n24669 = ~n24349 & ~n24668;
  assign n24670 = n24669 ^ n24348;
  assign n24671 = n24670 ^ n24342;
  assign n24672 = n24345 & ~n24671;
  assign n24673 = n24672 ^ n24344;
  assign n24676 = n24675 ^ n24673;
  assign n24677 = n23469 ^ n22573;
  assign n24678 = n24677 ^ n23482;
  assign n24679 = n24678 ^ n24675;
  assign n24680 = n24676 & n24679;
  assign n24681 = n24680 ^ n24678;
  assign n24682 = n24681 ^ n24340;
  assign n24683 = ~n24341 & n24682;
  assign n24684 = n24683 ^ n24339;
  assign n24685 = n24684 ^ n24336;
  assign n24686 = ~n24337 & n24685;
  assign n24687 = n24686 ^ n24335;
  assign n24688 = n24687 ^ n24330;
  assign n24689 = n24333 & n24688;
  assign n24690 = n24689 ^ n24332;
  assign n24328 = n24235 ^ n1974;
  assign n24329 = n24328 ^ n24178;
  assign n24691 = n24690 ^ n24329;
  assign n24692 = n24381 ^ n22559;
  assign n24693 = n24692 ^ n23554;
  assign n24694 = n24693 ^ n24690;
  assign n24695 = ~n24691 & ~n24694;
  assign n24696 = n24695 ^ n24329;
  assign n24697 = n24696 ^ n24322;
  assign n24698 = ~n24327 & n24697;
  assign n24699 = n24698 ^ n24326;
  assign n24701 = n24700 ^ n24699;
  assign n24702 = n24378 ^ n22554;
  assign n24703 = n24702 ^ n23545;
  assign n24704 = n24703 ^ n24700;
  assign n24705 = n24701 & ~n24704;
  assign n24706 = n24705 ^ n24703;
  assign n24708 = n24707 ^ n24706;
  assign n24709 = n24374 ^ n22549;
  assign n24710 = n24709 ^ n23539;
  assign n24711 = n24710 ^ n24707;
  assign n24712 = n24708 & ~n24711;
  assign n24713 = n24712 ^ n24710;
  assign n24319 = n24318 ^ n23534;
  assign n24320 = n24319 ^ n22548;
  assign n24749 = n24713 ^ n24320;
  assign n24315 = n24252 ^ n24169;
  assign n24316 = n24315 ^ n24166;
  assign n24750 = n24749 ^ n24316;
  assign n24751 = n24750 ^ n22323;
  assign n24752 = n24710 ^ n24708;
  assign n24753 = n24752 ^ n22309;
  assign n24834 = n24703 ^ n24701;
  assign n24754 = n24696 ^ n24327;
  assign n24755 = n24754 ^ n22279;
  assign n24756 = n24693 ^ n24329;
  assign n24757 = n24756 ^ n24690;
  assign n24758 = n24757 ^ n22225;
  assign n24759 = n24687 ^ n24333;
  assign n24760 = n24759 ^ n22113;
  assign n24761 = n24684 ^ n24335;
  assign n24762 = n24761 ^ n24336;
  assign n24763 = n24762 ^ n21644;
  assign n24817 = n24681 ^ n24341;
  assign n24764 = n24678 ^ n24676;
  assign n24765 = n24764 ^ n21648;
  assign n24809 = n24670 ^ n24345;
  assign n24804 = n24667 ^ n24349;
  assign n24766 = n24664 ^ n24662;
  assign n24767 = n24766 ^ n22080;
  assign n24796 = n24658 ^ n24354;
  assign n24768 = n24652 ^ n24624;
  assign n24769 = n24768 ^ n22067;
  assign n24782 = n24649 ^ n24626;
  assign n24783 = n24782 ^ n24628;
  assign n24770 = n24646 ^ n24634;
  assign n24771 = n24770 ^ n22057;
  assign n24772 = n24639 ^ n24637;
  assign n24773 = ~n21674 & n24772;
  assign n24774 = n24773 ^ n21670;
  assign n24775 = n24643 ^ n24641;
  assign n24776 = n24775 ^ n24773;
  assign n24777 = ~n24774 & ~n24776;
  assign n24778 = n24777 ^ n21670;
  assign n24779 = n24778 ^ n24770;
  assign n24780 = n24771 & ~n24779;
  assign n24781 = n24780 ^ n22057;
  assign n24784 = n24783 ^ n24781;
  assign n24785 = n24783 ^ n21668;
  assign n24786 = ~n24784 & ~n24785;
  assign n24787 = n24786 ^ n21668;
  assign n24788 = n24787 ^ n24768;
  assign n24789 = ~n24769 & n24788;
  assign n24790 = n24789 ^ n22067;
  assign n24791 = n24790 ^ n21663;
  assign n24792 = n24655 ^ n24358;
  assign n24793 = n24792 ^ n24790;
  assign n24794 = ~n24791 & n24793;
  assign n24795 = n24794 ^ n21663;
  assign n24797 = n24796 ^ n24795;
  assign n24798 = n24796 ^ n21658;
  assign n24799 = n24797 & ~n24798;
  assign n24800 = n24799 ^ n21658;
  assign n24801 = n24800 ^ n24766;
  assign n24802 = n24767 & n24801;
  assign n24803 = n24802 ^ n22080;
  assign n24805 = n24804 ^ n24803;
  assign n24806 = n24804 ^ n21650;
  assign n24807 = n24805 & ~n24806;
  assign n24808 = n24807 ^ n21650;
  assign n24810 = n24809 ^ n24808;
  assign n24811 = n24809 ^ n22090;
  assign n24812 = n24810 & n24811;
  assign n24813 = n24812 ^ n22090;
  assign n24814 = n24813 ^ n24764;
  assign n24815 = n24765 & ~n24814;
  assign n24816 = n24815 ^ n21648;
  assign n24818 = n24817 ^ n24816;
  assign n24819 = n24817 ^ n22100;
  assign n24820 = ~n24818 & ~n24819;
  assign n24821 = n24820 ^ n22100;
  assign n24822 = n24821 ^ n24762;
  assign n24823 = n24763 & n24822;
  assign n24824 = n24823 ^ n21644;
  assign n24825 = n24824 ^ n24759;
  assign n24826 = ~n24760 & n24825;
  assign n24827 = n24826 ^ n22113;
  assign n24828 = n24827 ^ n24757;
  assign n24829 = n24758 & n24828;
  assign n24830 = n24829 ^ n22225;
  assign n24831 = n24830 ^ n24754;
  assign n24832 = n24755 & n24831;
  assign n24833 = n24832 ^ n22279;
  assign n24835 = n24834 ^ n24833;
  assign n24836 = n24834 ^ n22294;
  assign n24837 = ~n24835 & n24836;
  assign n24838 = n24837 ^ n22294;
  assign n24839 = n24838 ^ n24752;
  assign n24840 = ~n24753 & ~n24839;
  assign n24841 = n24840 ^ n22309;
  assign n24842 = n24841 ^ n24750;
  assign n24843 = n24751 & ~n24842;
  assign n24844 = n24843 ^ n22323;
  assign n24321 = n24320 ^ n24316;
  assign n24714 = n24713 ^ n24316;
  assign n24715 = n24321 & ~n24714;
  assign n24716 = n24715 ^ n24320;
  assign n24312 = n24311 ^ n23530;
  assign n24313 = n24312 ^ n22542;
  assign n24746 = n24716 ^ n24313;
  assign n24310 = n24255 ^ n24165;
  assign n24747 = n24746 ^ n24310;
  assign n24748 = n24747 ^ n22337;
  assign n24925 = n24844 ^ n24748;
  assign n24880 = n24838 ^ n22309;
  assign n24881 = n24880 ^ n24752;
  assign n24882 = n24824 ^ n22113;
  assign n24883 = n24882 ^ n24759;
  assign n24884 = n24821 ^ n21644;
  assign n24885 = n24884 ^ n24762;
  assign n24886 = n24818 ^ n22100;
  assign n24887 = n24810 ^ n22090;
  assign n24888 = n24805 ^ n21650;
  assign n24889 = n24792 ^ n24791;
  assign n24890 = n24787 ^ n22067;
  assign n24891 = n24890 ^ n24768;
  assign n24892 = n24784 ^ n21668;
  assign n24893 = n24775 ^ n24774;
  assign n24894 = n24772 ^ n21674;
  assign n24895 = ~n24893 & ~n24894;
  assign n24896 = n24778 ^ n24771;
  assign n24897 = n24895 & ~n24896;
  assign n24898 = n24892 & n24897;
  assign n24899 = ~n24891 & n24898;
  assign n24900 = ~n24889 & ~n24899;
  assign n24901 = n24797 ^ n21658;
  assign n24902 = ~n24900 & n24901;
  assign n24903 = n24800 ^ n22080;
  assign n24904 = n24903 ^ n24766;
  assign n24905 = ~n24902 & n24904;
  assign n24906 = n24888 & n24905;
  assign n24907 = ~n24887 & n24906;
  assign n24908 = n24813 ^ n24765;
  assign n24909 = ~n24907 & ~n24908;
  assign n24910 = ~n24886 & ~n24909;
  assign n24911 = n24885 & ~n24910;
  assign n24912 = ~n24883 & ~n24911;
  assign n24913 = n24827 ^ n22225;
  assign n24914 = n24913 ^ n24757;
  assign n24915 = n24912 & n24914;
  assign n24916 = n24830 ^ n22279;
  assign n24917 = n24916 ^ n24754;
  assign n24918 = n24915 & ~n24917;
  assign n24919 = n24835 ^ n22294;
  assign n24920 = n24918 & n24919;
  assign n24921 = n24881 & ~n24920;
  assign n24922 = n24841 ^ n22323;
  assign n24923 = n24922 ^ n24750;
  assign n24924 = n24921 & n24923;
  assign n25084 = n24925 ^ n24924;
  assign n25076 = n24923 ^ n24921;
  assign n24960 = n24920 ^ n24881;
  assign n646 = n639 ^ n537;
  assign n653 = n652 ^ n646;
  assign n657 = n656 ^ n653;
  assign n24961 = n24960 ^ n657;
  assign n24962 = n24919 ^ n24918;
  assign n24966 = n24965 ^ n24962;
  assign n24967 = n24917 ^ n24915;
  assign n24971 = n24970 ^ n24967;
  assign n24972 = n24914 ^ n24912;
  assign n24976 = n24975 ^ n24972;
  assign n24977 = n24911 ^ n24883;
  assign n24981 = n24980 ^ n24977;
  assign n24982 = n24910 ^ n24885;
  assign n24986 = n24985 ^ n24982;
  assign n25053 = n24909 ^ n24886;
  assign n25048 = n24908 ^ n24907;
  assign n24987 = n24906 ^ n24887;
  assign n24988 = n24987 ^ n2226;
  assign n24989 = n24905 ^ n24888;
  assign n24990 = n24989 ^ n1826;
  assign n24991 = n24904 ^ n24902;
  assign n24995 = n24994 ^ n24991;
  assign n25034 = n24901 ^ n24900;
  assign n24996 = n24899 ^ n24889;
  assign n24997 = n24996 ^ n1636;
  assign n25026 = n24898 ^ n24891;
  assign n25001 = n24897 ^ n24892;
  assign n25002 = n25001 ^ n25000;
  assign n25006 = n24896 ^ n24895;
  assign n25007 = n25006 ^ n25005;
  assign n25011 = n24894 & n25010;
  assign n25015 = n25014 ^ n25011;
  assign n25016 = n24894 ^ n24893;
  assign n25017 = n25016 ^ n25014;
  assign n25018 = n25015 & ~n25017;
  assign n25019 = n25018 ^ n25011;
  assign n25020 = n25019 ^ n25006;
  assign n25021 = ~n25007 & n25020;
  assign n25022 = n25021 ^ n25005;
  assign n25023 = n25022 ^ n25001;
  assign n25024 = n25002 & ~n25023;
  assign n25025 = n25024 ^ n25000;
  assign n25027 = n25026 ^ n25025;
  assign n25028 = n25025 ^ n1614;
  assign n25029 = n25027 & n25028;
  assign n25030 = n25029 ^ n1614;
  assign n25031 = n25030 ^ n24996;
  assign n25032 = ~n24997 & n25031;
  assign n25033 = n25032 ^ n1636;
  assign n25035 = n25034 ^ n25033;
  assign n25036 = n25033 ^ n1704;
  assign n25037 = n25035 & n25036;
  assign n25038 = n25037 ^ n1704;
  assign n25039 = n25038 ^ n24991;
  assign n25040 = n24995 & ~n25039;
  assign n25041 = n25040 ^ n24994;
  assign n25042 = n25041 ^ n24989;
  assign n25043 = ~n24990 & n25042;
  assign n25044 = n25043 ^ n1826;
  assign n25045 = n25044 ^ n24987;
  assign n25046 = n24988 & ~n25045;
  assign n25047 = n25046 ^ n2226;
  assign n25049 = n25048 ^ n25047;
  assign n25050 = n25048 ^ n2236;
  assign n25051 = ~n25049 & n25050;
  assign n25052 = n25051 ^ n2236;
  assign n25054 = n25053 ^ n25052;
  assign n25055 = n25053 ^ n2250;
  assign n25056 = n25054 & ~n25055;
  assign n25057 = n25056 ^ n2250;
  assign n25058 = n25057 ^ n24982;
  assign n25059 = ~n24986 & n25058;
  assign n25060 = n25059 ^ n24985;
  assign n25061 = n25060 ^ n24977;
  assign n25062 = ~n24981 & n25061;
  assign n25063 = n25062 ^ n24980;
  assign n25064 = n25063 ^ n24972;
  assign n25065 = ~n24976 & n25064;
  assign n25066 = n25065 ^ n24975;
  assign n25067 = n25066 ^ n24967;
  assign n25068 = n24971 & ~n25067;
  assign n25069 = n25068 ^ n24970;
  assign n25070 = n25069 ^ n24962;
  assign n25071 = ~n24966 & n25070;
  assign n25072 = n25071 ^ n24965;
  assign n25073 = n25072 ^ n24960;
  assign n25074 = ~n24961 & n25073;
  assign n25075 = n25074 ^ n657;
  assign n25077 = n25076 ^ n25075;
  assign n25078 = n23067 ^ n15963;
  assign n25079 = n25078 ^ n661;
  assign n25080 = n25079 ^ n562;
  assign n25081 = n25080 ^ n25076;
  assign n25082 = ~n25077 & n25081;
  assign n25083 = n25082 ^ n25080;
  assign n25085 = n25084 ^ n25083;
  assign n25529 = n25085 ^ n569;
  assign n26340 = n25529 ^ n24304;
  assign n24944 = n24573 ^ n24557;
  assign n26341 = n26340 ^ n24944;
  assign n25270 = n24381 ^ n23560;
  assign n25271 = n25270 ^ n24707;
  assign n25269 = n25038 ^ n24995;
  assign n25272 = n25271 ^ n25269;
  assign n25274 = n24282 ^ n23475;
  assign n25275 = n25274 ^ n24700;
  assign n25273 = n25035 ^ n1704;
  assign n25276 = n25275 ^ n25273;
  assign n25279 = n24018 ^ n23489;
  assign n25280 = n25279 ^ n24329;
  assign n25278 = n25027 ^ n1614;
  assign n25281 = n25280 ^ n25278;
  assign n25284 = n23493 ^ n23469;
  assign n25285 = n25284 ^ n24330;
  assign n25282 = n25022 ^ n25000;
  assign n25283 = n25282 ^ n25001;
  assign n25286 = n25285 ^ n25283;
  assign n25287 = n24336 ^ n23474;
  assign n25288 = n25287 ^ n23498;
  assign n25221 = n25019 ^ n25005;
  assign n25222 = n25221 ^ n25006;
  assign n25289 = n25288 ^ n25222;
  assign n25355 = n25016 ^ n25015;
  assign n25290 = n24675 ^ n23508;
  assign n25291 = n25290 ^ n23481;
  assign n25224 = n25010 ^ n24894;
  assign n25292 = n25291 ^ n25224;
  assign n25334 = n23223 ^ n16339;
  assign n25335 = n25334 ^ n1547;
  assign n25336 = n25335 ^ n2639;
  assign n25131 = n24576 ^ n964;
  assign n25132 = n25131 ^ n24554;
  assign n25129 = n23243 ^ n22693;
  assign n25130 = n25129 ^ n23955;
  assign n25133 = n25132 ^ n25130;
  assign n24941 = n24616 ^ n23254;
  assign n24942 = n24941 ^ n22701;
  assign n25125 = n24944 ^ n24942;
  assign n24875 = n24570 ^ n24559;
  assign n24872 = n23249 ^ n22530;
  assign n24873 = n24872 ^ n24497;
  assign n24937 = n24875 ^ n24873;
  assign n24738 = n24567 ^ n24563;
  assign n24739 = n24738 ^ n24560;
  assign n24735 = n24432 ^ n23275;
  assign n24736 = n24735 ^ n23938;
  assign n24868 = n24739 ^ n24736;
  assign n24295 = n24294 ^ n23755;
  assign n24296 = n24295 ^ n23226;
  assign n24292 = n24291 ^ n24272;
  assign n24297 = n24296 ^ n24292;
  assign n24301 = n24269 ^ n24157;
  assign n24302 = n24301 ^ n24154;
  assign n24299 = n24298 ^ n23029;
  assign n24300 = n24299 ^ n23649;
  assign n24303 = n24302 ^ n24300;
  assign n24307 = n24266 ^ n24263;
  assign n24305 = n24304 ^ n22952;
  assign n24306 = n24305 ^ n23522;
  assign n24308 = n24307 ^ n24306;
  assign n24314 = n24313 ^ n24310;
  assign n24717 = n24716 ^ n24310;
  assign n24718 = n24314 & ~n24717;
  assign n24719 = n24718 ^ n24313;
  assign n24309 = n24258 ^ n24160;
  assign n24720 = n24719 ^ n24309;
  assign n24721 = n24369 ^ n23526;
  assign n24722 = n24721 ^ n22802;
  assign n24723 = n24722 ^ n24309;
  assign n24724 = ~n24720 & ~n24723;
  assign n24725 = n24724 ^ n24722;
  assign n24726 = n24725 ^ n24307;
  assign n24727 = n24308 & n24726;
  assign n24728 = n24727 ^ n24306;
  assign n24729 = n24728 ^ n24300;
  assign n24730 = n24303 & n24729;
  assign n24731 = n24730 ^ n24302;
  assign n24732 = n24731 ^ n24292;
  assign n24733 = ~n24297 & ~n24732;
  assign n24734 = n24733 ^ n24296;
  assign n24869 = n24739 ^ n24734;
  assign n24870 = n24868 & ~n24869;
  assign n24871 = n24870 ^ n24736;
  assign n24938 = n24875 ^ n24871;
  assign n24939 = n24937 & n24938;
  assign n24940 = n24939 ^ n24873;
  assign n25126 = n24944 ^ n24940;
  assign n25127 = n25125 & n25126;
  assign n25128 = n25127 ^ n24942;
  assign n25157 = n25130 ^ n25128;
  assign n25158 = n25133 & ~n25157;
  assign n25159 = n25158 ^ n25132;
  assign n25156 = n24581 ^ n976;
  assign n25160 = n25159 ^ n25156;
  assign n25154 = n23241 ^ n22691;
  assign n25155 = n25154 ^ n23958;
  assign n25201 = n25156 ^ n25155;
  assign n25202 = ~n25160 & n25201;
  assign n25203 = n25202 ^ n25155;
  assign n25198 = n23287 ^ n22685;
  assign n25199 = n25198 ^ n23962;
  assign n25197 = n24584 ^ n24553;
  assign n25200 = n25199 ^ n25197;
  assign n25204 = n25203 ^ n25200;
  assign n25205 = n25204 ^ n22035;
  assign n25161 = n25160 ^ n25155;
  assign n25162 = n25161 ^ n22012;
  assign n25134 = n25133 ^ n25128;
  assign n25135 = n25134 ^ n21983;
  assign n24874 = n24873 ^ n24871;
  assign n24876 = n24875 ^ n24874;
  assign n24737 = n24736 ^ n24734;
  assign n24740 = n24739 ^ n24737;
  assign n24741 = n24740 ^ n22544;
  assign n24859 = n24731 ^ n24296;
  assign n24860 = n24859 ^ n24292;
  assign n24854 = n24728 ^ n24303;
  assign n24742 = n24725 ^ n24308;
  assign n24743 = n24742 ^ n22614;
  assign n24744 = n24722 ^ n24720;
  assign n24745 = n24744 ^ n22518;
  assign n24845 = n24844 ^ n24747;
  assign n24846 = n24748 & ~n24845;
  assign n24847 = n24846 ^ n22337;
  assign n24848 = n24847 ^ n24744;
  assign n24849 = n24745 & n24848;
  assign n24850 = n24849 ^ n22518;
  assign n24851 = n24850 ^ n24742;
  assign n24852 = ~n24743 & ~n24851;
  assign n24853 = n24852 ^ n22614;
  assign n24855 = n24854 ^ n24853;
  assign n24856 = n24854 ^ n22551;
  assign n24857 = ~n24855 & ~n24856;
  assign n24858 = n24857 ^ n22551;
  assign n24861 = n24860 ^ n24858;
  assign n24862 = n24860 ^ n22645;
  assign n24863 = n24861 & ~n24862;
  assign n24864 = n24863 ^ n22645;
  assign n24865 = n24864 ^ n24740;
  assign n24866 = ~n24741 & n24865;
  assign n24867 = n24866 ^ n22544;
  assign n24877 = n24876 ^ n24867;
  assign n24946 = n24876 ^ n21938;
  assign n24947 = n24877 & n24946;
  assign n24948 = n24947 ^ n21938;
  assign n24943 = n24942 ^ n24940;
  assign n24945 = n24944 ^ n24943;
  assign n24949 = n24948 ^ n24945;
  assign n25122 = n24945 ^ n21960;
  assign n25123 = n24949 & n25122;
  assign n25124 = n25123 ^ n21960;
  assign n25151 = n25134 ^ n25124;
  assign n25152 = ~n25135 & n25151;
  assign n25153 = n25152 ^ n21983;
  assign n25194 = n25161 ^ n25153;
  assign n25195 = ~n25162 & n25194;
  assign n25196 = n25195 ^ n22012;
  assign n25206 = n25205 ^ n25196;
  assign n25136 = n25135 ^ n25124;
  assign n24878 = n24877 ^ n21938;
  assign n24879 = n24855 ^ n22551;
  assign n24926 = ~n24924 & ~n24925;
  assign n24927 = n24847 ^ n24745;
  assign n24928 = n24926 & ~n24927;
  assign n24929 = n24850 ^ n24743;
  assign n24930 = ~n24928 & n24929;
  assign n24931 = n24879 & ~n24930;
  assign n24932 = n24861 ^ n22645;
  assign n24933 = n24931 & ~n24932;
  assign n24934 = n24864 ^ n24741;
  assign n24935 = ~n24933 & n24934;
  assign n24936 = n24878 & ~n24935;
  assign n24950 = n24949 ^ n21960;
  assign n25137 = n24936 & ~n24950;
  assign n25150 = ~n25136 & n25137;
  assign n25163 = n25162 ^ n25153;
  assign n25207 = ~n25150 & n25163;
  assign n25298 = ~n25206 & ~n25207;
  assign n25307 = n25204 ^ n25196;
  assign n25308 = ~n25205 & ~n25307;
  assign n25309 = n25308 ^ n22035;
  assign n25310 = n25309 ^ n21679;
  assign n25303 = n22606 ^ n22538;
  assign n25304 = n25303 ^ n23969;
  assign n25302 = n24587 ^ n24551;
  assign n25305 = n25304 ^ n25302;
  assign n25299 = n25203 ^ n25199;
  assign n25300 = ~n25200 & ~n25299;
  assign n25301 = n25300 ^ n25197;
  assign n25306 = n25305 ^ n25301;
  assign n25311 = n25310 ^ n25306;
  assign n25331 = n25298 & ~n25311;
  assign n25327 = n23947 ^ n23300;
  assign n25328 = n25327 ^ n22602;
  assign n25325 = n24590 ^ n24546;
  assign n25322 = n25302 ^ n25301;
  assign n25323 = ~n25305 & ~n25322;
  assign n25324 = n25323 ^ n25304;
  assign n25326 = n25325 ^ n25324;
  assign n25329 = n25328 ^ n25326;
  assign n25317 = n25306 ^ n21679;
  assign n25318 = n25309 ^ n25306;
  assign n25319 = n25317 & ~n25318;
  assign n25320 = n25319 ^ n21679;
  assign n25321 = n25320 ^ n21675;
  assign n25330 = n25329 ^ n25321;
  assign n25332 = n25331 ^ n25330;
  assign n25312 = n25311 ^ n25298;
  assign n25209 = n23044 ^ n1541;
  assign n25210 = n25209 ^ n2368;
  assign n25211 = n25210 ^ n2484;
  assign n25208 = n25207 ^ n25206;
  assign n25212 = n25211 ^ n25208;
  assign n25164 = n25163 ^ n25150;
  assign n2352 = n2351 ^ n2315;
  assign n2353 = n2352 ^ n2348;
  assign n2357 = n2356 ^ n2353;
  assign n25165 = n25164 ^ n2357;
  assign n25138 = n25137 ^ n25136;
  assign n25146 = n25138 ^ n2295;
  assign n24951 = n24950 ^ n24936;
  assign n2298 = n2271 ^ n1324;
  assign n2299 = n2298 ^ n1251;
  assign n2300 = n2299 ^ n2286;
  assign n24952 = n24951 ^ n2300;
  assign n24953 = n24935 ^ n24878;
  assign n1239 = n1223 ^ n1145;
  assign n1240 = n1239 ^ n1236;
  assign n1244 = n1243 ^ n1240;
  assign n24954 = n24953 ^ n1244;
  assign n25110 = n24934 ^ n24933;
  assign n25105 = n24932 ^ n24931;
  assign n25100 = n24930 ^ n24879;
  assign n24955 = n24927 ^ n24926;
  assign n24959 = n24958 ^ n24955;
  assign n25086 = n25084 ^ n569;
  assign n25087 = n25085 & ~n25086;
  assign n25088 = n25087 ^ n569;
  assign n25089 = n25088 ^ n24955;
  assign n25090 = n24959 & ~n25089;
  assign n25091 = n25090 ^ n24958;
  assign n25095 = n25094 ^ n25091;
  assign n25096 = n24929 ^ n24928;
  assign n25097 = n25096 ^ n25091;
  assign n25098 = n25095 & n25097;
  assign n25099 = n25098 ^ n25094;
  assign n25101 = n25100 ^ n25099;
  assign n25102 = n25100 ^ n1087;
  assign n25103 = ~n25101 & n25102;
  assign n25104 = n25103 ^ n1087;
  assign n25106 = n25105 ^ n25104;
  assign n25107 = n25105 ^ n1076;
  assign n25108 = ~n25106 & n25107;
  assign n25109 = n25108 ^ n1076;
  assign n25111 = n25110 ^ n25109;
  assign n1101 = n1055 ^ n1020;
  assign n1102 = n1101 ^ n1096;
  assign n1106 = n1105 ^ n1102;
  assign n25112 = n25110 ^ n1106;
  assign n25113 = n25111 & ~n25112;
  assign n25114 = n25113 ^ n1106;
  assign n25115 = n25114 ^ n24953;
  assign n25116 = n24954 & ~n25115;
  assign n25117 = n25116 ^ n1244;
  assign n25118 = n25117 ^ n24951;
  assign n25119 = n24952 & ~n25118;
  assign n25120 = n25119 ^ n2300;
  assign n25147 = n25138 ^ n25120;
  assign n25148 = n25146 & ~n25147;
  assign n25149 = n25148 ^ n2295;
  assign n25191 = n25164 ^ n25149;
  assign n25192 = ~n25165 & n25191;
  assign n25193 = n25192 ^ n2357;
  assign n25295 = n25208 ^ n25193;
  assign n25296 = ~n25212 & n25295;
  assign n25297 = n25296 ^ n25211;
  assign n25313 = n25312 ^ n25297;
  assign n2490 = n2489 ^ n2429;
  assign n2491 = n2490 ^ n2486;
  assign n2492 = n2491 ^ n1514;
  assign n25314 = n25312 ^ n2492;
  assign n25315 = ~n25313 & n25314;
  assign n25316 = n25315 ^ n2492;
  assign n25333 = n25332 ^ n25316;
  assign n25337 = n25336 ^ n25333;
  assign n25293 = n24342 ^ n23486;
  assign n25294 = n25293 ^ n23513;
  assign n25338 = n25337 ^ n25294;
  assign n25342 = n24346 ^ n23465;
  assign n25343 = n25342 ^ n23492;
  assign n25213 = n25212 ^ n25193;
  assign n25189 = n24350 ^ n23497;
  assign n25190 = n25189 ^ n23440;
  assign n25214 = n25213 ^ n25190;
  assign n25121 = n25120 ^ n2295;
  assign n25139 = n25138 ^ n25121;
  assign n25140 = n24355 ^ n23507;
  assign n25141 = n25140 ^ n23308;
  assign n25169 = n25139 & n25141;
  assign n25167 = n23505 ^ n23354;
  assign n25168 = n25167 ^ n24351;
  assign n25170 = n25169 ^ n25168;
  assign n25166 = n25165 ^ n25149;
  assign n25186 = n25168 ^ n25166;
  assign n25187 = n25170 & n25186;
  assign n25188 = n25187 ^ n25169;
  assign n25339 = n25213 ^ n25188;
  assign n25340 = ~n25214 & n25339;
  assign n25341 = n25340 ^ n25190;
  assign n25344 = n25343 ^ n25341;
  assign n25345 = n25313 ^ n2492;
  assign n25346 = n25345 ^ n25341;
  assign n25347 = ~n25344 & ~n25346;
  assign n25348 = n25347 ^ n25343;
  assign n25349 = n25348 ^ n25337;
  assign n25350 = n25338 & ~n25349;
  assign n25351 = n25350 ^ n25294;
  assign n25352 = n25351 ^ n25291;
  assign n25353 = ~n25292 & ~n25352;
  assign n25354 = n25353 ^ n25224;
  assign n25356 = n25355 ^ n25354;
  assign n25357 = n23502 ^ n23478;
  assign n25358 = n25357 ^ n24340;
  assign n25359 = n25358 ^ n25355;
  assign n25360 = ~n25356 & ~n25359;
  assign n25361 = n25360 ^ n25358;
  assign n25362 = n25361 ^ n25222;
  assign n25363 = ~n25289 & ~n25362;
  assign n25364 = n25363 ^ n25288;
  assign n25365 = n25364 ^ n25283;
  assign n25366 = ~n25286 & ~n25365;
  assign n25367 = n25366 ^ n25285;
  assign n25368 = n25367 ^ n25278;
  assign n25369 = n25281 & ~n25368;
  assign n25370 = n25369 ^ n25280;
  assign n25277 = n25030 ^ n24997;
  assign n25371 = n25370 ^ n25277;
  assign n25372 = n24322 ^ n23482;
  assign n25373 = n25372 ^ n24111;
  assign n25374 = n25373 ^ n25277;
  assign n25375 = ~n25371 & ~n25374;
  assign n25376 = n25375 ^ n25373;
  assign n25377 = n25376 ^ n25273;
  assign n25378 = n25276 & n25377;
  assign n25379 = n25378 ^ n25275;
  assign n25380 = n25379 ^ n25269;
  assign n25381 = ~n25272 & n25380;
  assign n25382 = n25381 ^ n25271;
  assign n25266 = n24324 ^ n24316;
  assign n25267 = n25266 ^ n23470;
  assign n25264 = n25041 ^ n1826;
  assign n25265 = n25264 ^ n24989;
  assign n25268 = n25267 ^ n25265;
  assign n25434 = n25382 ^ n25268;
  assign n25435 = n25434 ^ n22563;
  assign n25436 = n25379 ^ n25272;
  assign n25437 = n25436 ^ n22768;
  assign n25438 = n25376 ^ n25276;
  assign n25439 = n25438 ^ n22567;
  assign n25478 = n25373 ^ n25371;
  assign n25440 = n25367 ^ n25281;
  assign n25441 = n25440 ^ n22577;
  assign n25442 = n25361 ^ n25289;
  assign n25443 = n25442 ^ n22585;
  assign n25444 = n25358 ^ n25356;
  assign n25445 = n25444 ^ n22746;
  assign n25446 = n25351 ^ n25292;
  assign n25447 = n25446 ^ n22589;
  assign n25448 = n25348 ^ n25338;
  assign n25449 = n25448 ^ n22736;
  assign n25450 = n25345 ^ n25344;
  assign n25451 = n25450 ^ n22729;
  assign n25215 = n25214 ^ n25188;
  assign n25216 = n25215 ^ n22591;
  assign n25142 = n25141 ^ n25139;
  assign n25172 = n22598 & n25142;
  assign n25173 = n25172 ^ n22540;
  assign n25171 = n25170 ^ n25166;
  assign n25183 = n25172 ^ n25171;
  assign n25184 = n25173 & n25183;
  assign n25185 = n25184 ^ n22540;
  assign n25452 = n25215 ^ n25185;
  assign n25453 = n25216 & n25452;
  assign n25454 = n25453 ^ n22591;
  assign n25455 = n25454 ^ n25450;
  assign n25456 = ~n25451 & ~n25455;
  assign n25457 = n25456 ^ n22729;
  assign n25458 = n25457 ^ n25448;
  assign n25459 = n25449 & n25458;
  assign n25460 = n25459 ^ n22736;
  assign n25461 = n25460 ^ n25446;
  assign n25462 = ~n25447 & n25461;
  assign n25463 = n25462 ^ n22589;
  assign n25464 = n25463 ^ n25444;
  assign n25465 = n25445 & ~n25464;
  assign n25466 = n25465 ^ n22746;
  assign n25467 = n25466 ^ n25442;
  assign n25468 = n25443 & n25467;
  assign n25469 = n25468 ^ n22585;
  assign n25470 = n25469 ^ n22581;
  assign n25471 = n25364 ^ n25286;
  assign n25472 = n25471 ^ n25469;
  assign n25473 = n25470 & n25472;
  assign n25474 = n25473 ^ n22581;
  assign n25475 = n25474 ^ n25440;
  assign n25476 = ~n25441 & n25475;
  assign n25477 = n25476 ^ n22577;
  assign n25479 = n25478 ^ n25477;
  assign n25480 = n25478 ^ n22573;
  assign n25481 = ~n25479 & n25480;
  assign n25482 = n25481 ^ n22573;
  assign n25483 = n25482 ^ n25438;
  assign n25484 = ~n25439 & ~n25483;
  assign n25485 = n25484 ^ n22567;
  assign n25486 = n25485 ^ n25436;
  assign n25487 = ~n25437 & n25486;
  assign n25488 = n25487 ^ n22768;
  assign n25489 = n25488 ^ n25434;
  assign n25490 = n25435 & n25489;
  assign n25491 = n25490 ^ n22563;
  assign n25593 = n25491 ^ n22559;
  assign n25383 = n25382 ^ n25265;
  assign n25384 = ~n25268 & ~n25383;
  assign n25385 = n25384 ^ n25267;
  assign n25262 = n25044 ^ n24988;
  assign n25260 = n24378 ^ n23554;
  assign n25261 = n25260 ^ n24310;
  assign n25263 = n25262 ^ n25261;
  assign n25432 = n25385 ^ n25263;
  assign n25594 = n25593 ^ n25432;
  assign n25566 = n25488 ^ n25435;
  assign n25567 = n25485 ^ n25437;
  assign n25568 = n25482 ^ n22567;
  assign n25569 = n25568 ^ n25438;
  assign n25570 = n25479 ^ n22573;
  assign n25571 = n25474 ^ n25441;
  assign n25572 = n25466 ^ n25443;
  assign n25573 = n25460 ^ n22589;
  assign n25574 = n25573 ^ n25446;
  assign n25575 = n25457 ^ n25449;
  assign n25143 = n25142 ^ n22598;
  assign n25174 = n25173 ^ n25171;
  assign n25182 = n25143 & ~n25174;
  assign n25217 = n25216 ^ n25185;
  assign n25576 = n25182 & n25217;
  assign n25577 = n25454 ^ n22729;
  assign n25578 = n25577 ^ n25450;
  assign n25579 = n25576 & n25578;
  assign n25580 = n25575 & n25579;
  assign n25581 = ~n25574 & ~n25580;
  assign n25582 = n25463 ^ n22746;
  assign n25583 = n25582 ^ n25444;
  assign n25584 = ~n25581 & ~n25583;
  assign n25585 = n25572 & ~n25584;
  assign n25586 = n25471 ^ n25470;
  assign n25587 = n25585 & n25586;
  assign n25588 = n25571 & n25587;
  assign n25589 = n25570 & ~n25588;
  assign n25590 = n25569 & ~n25589;
  assign n25591 = n25567 & ~n25590;
  assign n25592 = n25566 & ~n25591;
  assign n25715 = n25594 ^ n25592;
  assign n25691 = n25589 ^ n25569;
  assign n25639 = n25587 ^ n25571;
  assign n25640 = n25639 ^ n1930;
  assign n25641 = n25584 ^ n25572;
  assign n25642 = n25641 ^ n1802;
  assign n25670 = n25583 ^ n25581;
  assign n25662 = n25580 ^ n25574;
  assign n25643 = n25579 ^ n25575;
  assign n25647 = n25646 ^ n25643;
  assign n25648 = n25578 ^ n25576;
  assign n25652 = n25651 ^ n25648;
  assign n25218 = n25217 ^ n25182;
  assign n25219 = n25218 ^ n25181;
  assign n2649 = n2648 ^ n2642;
  assign n2653 = n2652 ^ n2649;
  assign n2654 = n2653 ^ n1499;
  assign n25144 = n2654 & ~n25143;
  assign n1554 = n1553 ^ n1430;
  assign n1555 = n1554 ^ n1523;
  assign n1556 = n1555 ^ n1466;
  assign n25145 = n25144 ^ n1556;
  assign n25175 = n25174 ^ n25143;
  assign n25176 = n25175 ^ n1556;
  assign n25177 = n25145 & n25176;
  assign n25178 = n25177 ^ n25144;
  assign n25653 = n25218 ^ n25178;
  assign n25654 = n25219 & ~n25653;
  assign n25655 = n25654 ^ n25181;
  assign n25656 = n25655 ^ n25648;
  assign n25657 = n25652 & ~n25656;
  assign n25658 = n25657 ^ n25651;
  assign n25659 = n25658 ^ n25643;
  assign n25660 = n25647 & ~n25659;
  assign n25661 = n25660 ^ n25646;
  assign n25663 = n25662 ^ n25661;
  assign n25667 = n25666 ^ n25662;
  assign n25668 = n25663 & ~n25667;
  assign n25669 = n25668 ^ n25666;
  assign n25671 = n25670 ^ n25669;
  assign n1779 = n1724 ^ n1683;
  assign n1786 = n1785 ^ n1779;
  assign n1790 = n1789 ^ n1786;
  assign n25672 = n25670 ^ n1790;
  assign n25673 = ~n25671 & n25672;
  assign n25674 = n25673 ^ n1790;
  assign n25675 = n25674 ^ n25641;
  assign n25676 = n25642 & ~n25675;
  assign n25677 = n25676 ^ n1802;
  assign n25678 = n25677 ^ n1918;
  assign n25679 = n25586 ^ n25585;
  assign n25680 = n25679 ^ n25677;
  assign n25681 = n25678 & n25680;
  assign n25682 = n25681 ^ n1918;
  assign n25683 = n25682 ^ n25639;
  assign n25684 = ~n25640 & n25683;
  assign n25685 = n25684 ^ n1930;
  assign n25686 = n25685 ^ n2085;
  assign n25687 = n25588 ^ n25570;
  assign n25688 = n25687 ^ n25685;
  assign n25689 = n25686 & n25688;
  assign n25690 = n25689 ^ n2085;
  assign n25692 = n25691 ^ n25690;
  assign n25696 = n25695 ^ n25691;
  assign n25697 = ~n25692 & n25696;
  assign n25698 = n25697 ^ n25695;
  assign n25702 = n25701 ^ n25698;
  assign n25703 = n25590 ^ n25567;
  assign n25704 = n25703 ^ n25698;
  assign n25705 = n25702 & n25704;
  assign n25706 = n25705 ^ n25701;
  assign n25710 = n25709 ^ n25706;
  assign n25711 = n25591 ^ n25566;
  assign n25712 = n25711 ^ n25706;
  assign n25713 = n25710 & ~n25712;
  assign n25714 = n25713 ^ n25709;
  assign n25716 = n25715 ^ n25714;
  assign n26339 = n25719 ^ n25716;
  assign n26342 = n26341 ^ n26339;
  assign n26258 = n25711 ^ n25710;
  assign n25413 = n25080 ^ n25077;
  assign n26255 = n25413 ^ n24369;
  assign n26256 = n26255 ^ n24875;
  assign n26343 = n26258 ^ n26256;
  assign n26234 = n25703 ^ n25702;
  assign n25227 = n25072 ^ n24961;
  assign n26231 = n25227 ^ n24739;
  assign n26232 = n26231 ^ n24311;
  assign n26251 = n26234 ^ n26232;
  assign n26077 = n25695 ^ n25692;
  assign n26063 = n25687 ^ n2085;
  assign n26064 = n26063 ^ n25685;
  assign n26051 = n25682 ^ n25640;
  assign n25975 = n25679 ^ n25678;
  assign n25243 = n25060 ^ n24980;
  assign n25244 = n25243 ^ n24977;
  assign n25973 = n25244 ^ n24309;
  assign n25974 = n25973 ^ n24324;
  assign n25976 = n25975 ^ n25974;
  assign n25811 = n24381 ^ n24310;
  assign n25248 = n25057 ^ n24986;
  assign n25812 = n25811 ^ n25248;
  assign n25809 = n25674 ^ n1802;
  assign n25810 = n25809 ^ n25641;
  assign n25813 = n25812 ^ n25810;
  assign n25252 = n25054 ^ n2250;
  assign n25815 = n25252 ^ n24282;
  assign n25816 = n25815 ^ n24316;
  assign n25814 = n25671 ^ n1790;
  assign n25817 = n25816 ^ n25814;
  assign n25256 = n25049 ^ n2236;
  assign n25819 = n25256 ^ n24111;
  assign n25820 = n25819 ^ n24707;
  assign n25818 = n25666 ^ n25663;
  assign n25821 = n25820 ^ n25818;
  assign n25956 = n25658 ^ n25646;
  assign n25957 = n25956 ^ n25643;
  assign n25823 = n24322 ^ n23469;
  assign n25824 = n25823 ^ n25265;
  assign n25822 = n25655 ^ n25652;
  assign n25825 = n25824 ^ n25822;
  assign n25826 = n25269 ^ n23474;
  assign n25827 = n25826 ^ n24329;
  assign n25220 = n25219 ^ n25178;
  assign n25828 = n25827 ^ n25220;
  assign n25830 = n25273 ^ n24330;
  assign n25831 = n25830 ^ n23478;
  assign n25829 = n25175 ^ n25145;
  assign n25832 = n25831 ^ n25829;
  assign n25834 = n25277 ^ n23481;
  assign n25835 = n25834 ^ n24336;
  assign n25833 = n25143 ^ n2654;
  assign n25836 = n25835 ^ n25833;
  assign n25915 = n25278 ^ n23486;
  assign n25916 = n25915 ^ n24340;
  assign n25857 = n24631 ^ n23287;
  assign n25858 = n25857 ^ n23947;
  assign n25856 = n25111 ^ n1106;
  assign n25859 = n25858 ^ n25856;
  assign n25841 = n24643 ^ n23241;
  assign n25842 = n25841 ^ n23969;
  assign n25840 = n25106 ^ n1076;
  assign n25843 = n25842 ^ n25840;
  assign n25555 = n25096 ^ n25095;
  assign n25553 = n25325 ^ n23254;
  assign n25554 = n25553 ^ n23958;
  assign n25556 = n25555 ^ n25554;
  assign n25543 = n25088 ^ n24959;
  assign n25541 = n25302 ^ n23249;
  assign n25542 = n25541 ^ n23955;
  assign n25544 = n25543 ^ n25542;
  assign n25530 = n25197 ^ n24616;
  assign n25531 = n25530 ^ n23938;
  assign n25532 = n25531 ^ n25529;
  assign n25414 = n25156 ^ n24497;
  assign n25415 = n25414 ^ n23755;
  assign n25416 = n25415 ^ n25413;
  assign n25228 = n25132 ^ n23649;
  assign n25229 = n25228 ^ n24432;
  assign n25230 = n25229 ^ n25227;
  assign n25233 = n25069 ^ n24966;
  assign n25231 = n24944 ^ n23522;
  assign n25232 = n25231 ^ n24294;
  assign n25234 = n25233 ^ n25232;
  assign n25237 = n25066 ^ n24971;
  assign n25235 = n24298 ^ n23526;
  assign n25236 = n25235 ^ n24875;
  assign n25238 = n25237 ^ n25236;
  assign n25241 = n25063 ^ n24976;
  assign n25239 = n24739 ^ n23530;
  assign n25240 = n25239 ^ n24304;
  assign n25242 = n25241 ^ n25240;
  assign n25245 = n24369 ^ n23534;
  assign n25246 = n25245 ^ n24292;
  assign n25247 = n25246 ^ n25244;
  assign n25249 = n24311 ^ n23539;
  assign n25250 = n25249 ^ n24302;
  assign n25251 = n25250 ^ n25248;
  assign n25253 = n24307 ^ n23545;
  assign n25254 = n25253 ^ n24318;
  assign n25255 = n25254 ^ n25252;
  assign n25257 = n24374 ^ n24309;
  assign n25258 = n25257 ^ n23550;
  assign n25259 = n25258 ^ n25256;
  assign n25386 = n25385 ^ n25262;
  assign n25387 = n25263 & ~n25386;
  assign n25388 = n25387 ^ n25261;
  assign n25389 = n25388 ^ n25256;
  assign n25390 = n25259 & ~n25389;
  assign n25391 = n25390 ^ n25258;
  assign n25392 = n25391 ^ n25252;
  assign n25393 = n25255 & n25392;
  assign n25394 = n25393 ^ n25254;
  assign n25395 = n25394 ^ n25248;
  assign n25396 = n25251 & ~n25395;
  assign n25397 = n25396 ^ n25250;
  assign n25398 = n25397 ^ n25244;
  assign n25399 = ~n25247 & ~n25398;
  assign n25400 = n25399 ^ n25246;
  assign n25401 = n25400 ^ n25241;
  assign n25402 = n25242 & n25401;
  assign n25403 = n25402 ^ n25240;
  assign n25404 = n25403 ^ n25236;
  assign n25405 = n25238 & n25404;
  assign n25406 = n25405 ^ n25237;
  assign n25407 = n25406 ^ n25233;
  assign n25408 = ~n25234 & n25407;
  assign n25409 = n25408 ^ n25232;
  assign n25410 = n25409 ^ n25227;
  assign n25411 = n25230 & n25410;
  assign n25412 = n25411 ^ n25229;
  assign n25526 = n25413 ^ n25412;
  assign n25527 = n25416 & n25526;
  assign n25528 = n25527 ^ n25415;
  assign n25538 = n25531 ^ n25528;
  assign n25539 = ~n25532 & ~n25538;
  assign n25540 = n25539 ^ n25529;
  assign n25550 = n25542 ^ n25540;
  assign n25551 = n25544 & n25550;
  assign n25552 = n25551 ^ n25543;
  assign n25783 = n25555 ^ n25552;
  assign n25784 = ~n25556 & n25783;
  assign n25785 = n25784 ^ n25554;
  assign n25782 = n25101 ^ n1087;
  assign n25786 = n25785 ^ n25782;
  assign n25780 = n24637 ^ n23962;
  assign n25781 = n25780 ^ n23243;
  assign n25844 = n25782 ^ n25781;
  assign n25845 = ~n25786 & ~n25844;
  assign n25846 = n25845 ^ n25781;
  assign n25853 = n25846 ^ n25840;
  assign n25854 = ~n25843 & n25853;
  assign n25855 = n25854 ^ n25842;
  assign n25867 = n25856 ^ n25855;
  assign n25868 = ~n25859 & ~n25867;
  assign n25869 = n25868 ^ n25858;
  assign n25864 = n24628 ^ n22538;
  assign n25865 = n25864 ^ n23517;
  assign n25802 = n25114 ^ n24954;
  assign n25866 = n25865 ^ n25802;
  assign n25870 = n25869 ^ n25866;
  assign n25871 = n25870 ^ n22606;
  assign n25847 = n25846 ^ n25843;
  assign n25787 = n25786 ^ n25781;
  assign n25557 = n25556 ^ n25552;
  assign n25545 = n25544 ^ n25540;
  assign n25533 = n25532 ^ n25528;
  assign n25417 = n25416 ^ n25412;
  assign n25418 = n25417 ^ n23226;
  assign n25518 = n25410 ^ n25229;
  assign n25419 = n25406 ^ n25234;
  assign n25420 = n25419 ^ n22952;
  assign n25421 = n25403 ^ n25238;
  assign n25422 = n25421 ^ n22802;
  assign n25423 = n25400 ^ n25242;
  assign n25424 = n25423 ^ n22542;
  assign n25425 = n25394 ^ n25251;
  assign n25426 = n25425 ^ n22549;
  assign n25427 = n25391 ^ n25255;
  assign n25428 = n25427 ^ n22554;
  assign n25429 = n25388 ^ n25258;
  assign n25430 = n25429 ^ n25256;
  assign n25431 = n25430 ^ n22555;
  assign n25433 = n25432 ^ n22559;
  assign n25492 = n25491 ^ n25432;
  assign n25493 = n25433 & ~n25492;
  assign n25494 = n25493 ^ n22559;
  assign n25495 = n25494 ^ n25430;
  assign n25496 = ~n25431 & ~n25495;
  assign n25497 = n25496 ^ n22555;
  assign n25498 = n25497 ^ n25427;
  assign n25499 = n25428 & n25498;
  assign n25500 = n25499 ^ n22554;
  assign n25501 = n25500 ^ n25425;
  assign n25502 = n25426 & n25501;
  assign n25503 = n25502 ^ n22549;
  assign n25504 = n25503 ^ n22548;
  assign n25505 = n25397 ^ n25247;
  assign n25506 = n25505 ^ n25503;
  assign n25507 = ~n25504 & n25506;
  assign n25508 = n25507 ^ n22548;
  assign n25509 = n25508 ^ n25423;
  assign n25510 = n25424 & ~n25509;
  assign n25511 = n25510 ^ n22542;
  assign n25512 = n25511 ^ n25421;
  assign n25513 = n25422 & n25512;
  assign n25514 = n25513 ^ n22802;
  assign n25515 = n25514 ^ n25419;
  assign n25516 = ~n25420 & ~n25515;
  assign n25517 = n25516 ^ n22952;
  assign n25519 = n25518 ^ n25517;
  assign n25520 = n25518 ^ n23029;
  assign n25521 = ~n25519 & n25520;
  assign n25522 = n25521 ^ n23029;
  assign n25523 = n25522 ^ n25417;
  assign n25524 = ~n25418 & n25523;
  assign n25525 = n25524 ^ n23226;
  assign n25534 = n25533 ^ n25525;
  assign n25535 = n25525 ^ n23275;
  assign n25536 = n25534 & ~n25535;
  assign n25537 = n25536 ^ n23275;
  assign n25546 = n25545 ^ n25537;
  assign n25547 = n25545 ^ n22530;
  assign n25548 = ~n25546 & n25547;
  assign n25549 = n25548 ^ n22530;
  assign n25558 = n25557 ^ n25549;
  assign n25777 = n25557 ^ n22701;
  assign n25778 = ~n25558 & ~n25777;
  assign n25779 = n25778 ^ n22701;
  assign n25788 = n25787 ^ n25779;
  assign n25837 = n25787 ^ n22693;
  assign n25838 = n25788 & ~n25837;
  assign n25839 = n25838 ^ n22693;
  assign n25848 = n25847 ^ n25839;
  assign n25849 = n25847 ^ n22691;
  assign n25850 = ~n25848 & ~n25849;
  assign n25851 = n25850 ^ n22691;
  assign n25852 = n25851 ^ n22685;
  assign n25860 = n25859 ^ n25855;
  assign n25861 = n25860 ^ n25851;
  assign n25862 = n25852 & n25861;
  assign n25863 = n25862 ^ n22685;
  assign n25872 = n25871 ^ n25863;
  assign n25873 = n25860 ^ n22685;
  assign n25874 = n25873 ^ n25851;
  assign n25875 = n25848 ^ n22691;
  assign n25789 = n25788 ^ n22693;
  assign n25559 = n25558 ^ n22701;
  assign n25560 = n25546 ^ n22530;
  assign n25561 = n25533 ^ n23275;
  assign n25562 = n25561 ^ n25525;
  assign n25563 = n25508 ^ n25424;
  assign n25564 = n25500 ^ n25426;
  assign n25565 = n25497 ^ n25428;
  assign n25595 = n25592 & ~n25594;
  assign n25596 = n25494 ^ n25431;
  assign n25597 = n25595 & n25596;
  assign n25598 = n25565 & n25597;
  assign n25599 = n25564 & ~n25598;
  assign n25600 = n25505 ^ n22548;
  assign n25601 = n25600 ^ n25503;
  assign n25602 = n25599 & ~n25601;
  assign n25603 = ~n25563 & ~n25602;
  assign n25604 = n25511 ^ n25422;
  assign n25605 = n25603 & ~n25604;
  assign n25606 = n25514 ^ n25420;
  assign n25607 = ~n25605 & n25606;
  assign n25608 = n25519 ^ n23029;
  assign n25609 = ~n25607 & ~n25608;
  assign n25610 = n25522 ^ n25418;
  assign n25611 = n25609 & n25610;
  assign n25612 = n25562 & ~n25611;
  assign n25613 = n25560 & ~n25612;
  assign n25790 = ~n25559 & n25613;
  assign n25876 = n25789 & n25790;
  assign n25877 = ~n25875 & ~n25876;
  assign n25878 = ~n25874 & ~n25877;
  assign n25911 = ~n25872 & n25878;
  assign n25907 = n25117 ^ n24952;
  assign n25905 = n24623 ^ n23512;
  assign n25906 = n25905 ^ n23300;
  assign n25908 = n25907 ^ n25906;
  assign n25902 = n25869 ^ n25865;
  assign n25903 = ~n25866 & n25902;
  assign n25904 = n25903 ^ n25869;
  assign n25909 = n25908 ^ n25904;
  assign n25898 = n25870 ^ n25863;
  assign n25899 = ~n25871 & n25898;
  assign n25900 = n25899 ^ n22606;
  assign n25901 = n25900 ^ n22602;
  assign n25910 = n25909 ^ n25901;
  assign n25912 = n25911 ^ n25910;
  assign n25913 = n25912 ^ n2555;
  assign n25879 = n25878 ^ n25872;
  assign n2574 = n2566 ^ n2497;
  assign n2575 = n2574 ^ n2466;
  assign n2576 = n2575 ^ n2551;
  assign n25880 = n25879 ^ n2576;
  assign n25881 = n25877 ^ n25874;
  assign n25882 = n25881 ^ n2446;
  assign n25883 = n25876 ^ n25875;
  assign n2449 = n2384 ^ n2343;
  assign n2456 = n2455 ^ n2449;
  assign n2457 = n2456 ^ n2437;
  assign n25884 = n25883 ^ n2457;
  assign n25791 = n25790 ^ n25789;
  assign n25773 = n23810 ^ n2331;
  assign n25774 = n25773 ^ n1406;
  assign n25775 = n25774 ^ n2452;
  assign n25885 = n25791 ^ n25775;
  assign n25614 = n25613 ^ n25559;
  assign n1394 = n1351 ^ n1288;
  assign n1395 = n1394 ^ n1388;
  assign n1396 = n1395 ^ n1304;
  assign n25615 = n25614 ^ n1396;
  assign n25616 = n25612 ^ n25560;
  assign n25617 = n25616 ^ n1381;
  assign n25762 = n25611 ^ n25562;
  assign n25757 = n25610 ^ n25609;
  assign n25618 = n25608 ^ n25607;
  assign n25622 = n25621 ^ n25618;
  assign n25623 = n25606 ^ n25605;
  assign n25624 = n25623 ^ n828;
  assign n25625 = n25604 ^ n25603;
  assign n727 = n724 ^ n706;
  assign n734 = n733 ^ n727;
  assign n738 = n737 ^ n734;
  assign n25626 = n25625 ^ n738;
  assign n25627 = n25602 ^ n25563;
  assign n741 = n717 ^ n694;
  assign n748 = n747 ^ n741;
  assign n749 = n748 ^ n731;
  assign n25628 = n25627 ^ n749;
  assign n25629 = n25601 ^ n25599;
  assign n25633 = n25632 ^ n25629;
  assign n25734 = n25598 ^ n25564;
  assign n25634 = n25597 ^ n25565;
  assign n25638 = n25637 ^ n25634;
  assign n25723 = n25596 ^ n25595;
  assign n25720 = n25719 ^ n25715;
  assign n25721 = ~n25716 & n25720;
  assign n25722 = n25721 ^ n25719;
  assign n25724 = n25723 ^ n25722;
  assign n25728 = n25727 ^ n25722;
  assign n25729 = n25724 & n25728;
  assign n25730 = n25729 ^ n25727;
  assign n25731 = n25730 ^ n25634;
  assign n25732 = ~n25638 & n25731;
  assign n25733 = n25732 ^ n25637;
  assign n25735 = n25734 ^ n25733;
  assign n25739 = n25738 ^ n25734;
  assign n25740 = n25735 & ~n25739;
  assign n25741 = n25740 ^ n25738;
  assign n25742 = n25741 ^ n25629;
  assign n25743 = ~n25633 & n25742;
  assign n25744 = n25743 ^ n25632;
  assign n25745 = n25744 ^ n25627;
  assign n25746 = ~n25628 & n25745;
  assign n25747 = n25746 ^ n749;
  assign n25748 = n25747 ^ n25625;
  assign n25749 = n25626 & ~n25748;
  assign n25750 = n25749 ^ n738;
  assign n25751 = n25750 ^ n25623;
  assign n25752 = ~n25624 & n25751;
  assign n25753 = n25752 ^ n828;
  assign n25754 = n25753 ^ n25618;
  assign n25755 = ~n25622 & n25754;
  assign n25756 = n25755 ^ n25621;
  assign n25758 = n25757 ^ n25756;
  assign n25759 = n25757 ^ n956;
  assign n25760 = n25758 & ~n25759;
  assign n25761 = n25760 ^ n956;
  assign n25763 = n25762 ^ n25761;
  assign n25764 = n25762 ^ n1372;
  assign n25765 = n25763 & ~n25764;
  assign n25766 = n25765 ^ n1372;
  assign n25767 = n25766 ^ n1381;
  assign n25768 = n25617 & ~n25767;
  assign n25769 = n25768 ^ n25616;
  assign n25770 = n25769 ^ n25614;
  assign n25771 = n25615 & ~n25770;
  assign n25772 = n25771 ^ n1396;
  assign n25886 = n25791 ^ n25772;
  assign n25887 = ~n25885 & n25886;
  assign n25888 = n25887 ^ n25775;
  assign n25889 = n25888 ^ n25883;
  assign n25890 = n25884 & ~n25889;
  assign n25891 = n25890 ^ n2457;
  assign n25892 = n25891 ^ n2446;
  assign n25893 = ~n25882 & ~n25892;
  assign n25894 = n25893 ^ n25881;
  assign n25895 = n25894 ^ n25879;
  assign n25896 = n25880 & n25895;
  assign n25897 = n25896 ^ n2576;
  assign n25914 = n25913 ^ n25897;
  assign n25917 = n25916 ^ n25914;
  assign n25919 = n25283 ^ n23492;
  assign n25920 = n25919 ^ n24675;
  assign n25918 = n25894 ^ n25880;
  assign n25921 = n25920 ^ n25918;
  assign n25931 = n24342 ^ n23497;
  assign n25932 = n25931 ^ n25222;
  assign n25923 = n25355 ^ n24346;
  assign n25924 = n25923 ^ n23505;
  assign n25225 = n25224 ^ n23507;
  assign n25226 = n25225 ^ n24350;
  assign n25776 = n25775 ^ n25772;
  assign n25792 = n25791 ^ n25776;
  assign n25922 = n25226 & ~n25792;
  assign n25925 = n25924 ^ n25922;
  assign n25926 = n25888 ^ n2457;
  assign n25927 = n25926 ^ n25883;
  assign n25928 = n25927 ^ n25922;
  assign n25929 = n25925 & ~n25928;
  assign n25930 = n25929 ^ n25924;
  assign n25933 = n25932 ^ n25930;
  assign n25934 = n25891 ^ n25882;
  assign n25935 = n25934 ^ n25930;
  assign n25936 = n25933 & n25935;
  assign n25937 = n25936 ^ n25932;
  assign n25938 = n25937 ^ n25918;
  assign n25939 = ~n25921 & n25938;
  assign n25940 = n25939 ^ n25920;
  assign n25941 = n25940 ^ n25914;
  assign n25942 = n25917 & n25941;
  assign n25943 = n25942 ^ n25916;
  assign n25944 = n25943 ^ n25833;
  assign n25945 = ~n25836 & ~n25944;
  assign n25946 = n25945 ^ n25835;
  assign n25947 = n25946 ^ n25829;
  assign n25948 = n25832 & n25947;
  assign n25949 = n25948 ^ n25831;
  assign n25950 = n25949 ^ n25827;
  assign n25951 = ~n25828 & ~n25950;
  assign n25952 = n25951 ^ n25220;
  assign n25953 = n25952 ^ n25822;
  assign n25954 = n25825 & ~n25953;
  assign n25955 = n25954 ^ n25824;
  assign n25958 = n25957 ^ n25955;
  assign n25959 = n25262 ^ n24700;
  assign n25960 = n25959 ^ n24018;
  assign n25961 = n25960 ^ n25957;
  assign n25962 = ~n25958 & n25961;
  assign n25963 = n25962 ^ n25960;
  assign n25964 = n25963 ^ n25818;
  assign n25965 = ~n25821 & n25964;
  assign n25966 = n25965 ^ n25820;
  assign n25967 = n25966 ^ n25814;
  assign n25968 = ~n25817 & ~n25967;
  assign n25969 = n25968 ^ n25816;
  assign n25970 = n25969 ^ n25812;
  assign n25971 = ~n25813 & ~n25970;
  assign n25972 = n25971 ^ n25810;
  assign n26048 = n25975 ^ n25972;
  assign n26049 = ~n25976 & n26048;
  assign n26050 = n26049 ^ n25974;
  assign n26052 = n26051 ^ n26050;
  assign n26046 = n25241 ^ n24378;
  assign n26047 = n26046 ^ n24307;
  assign n26060 = n26051 ^ n26047;
  assign n26061 = n26052 & ~n26060;
  assign n26062 = n26061 ^ n26047;
  assign n26065 = n26064 ^ n26062;
  assign n26058 = n25237 ^ n24302;
  assign n26059 = n26058 ^ n24374;
  assign n26074 = n26064 ^ n26059;
  assign n26075 = n26065 & n26074;
  assign n26076 = n26075 ^ n26059;
  assign n26078 = n26077 ^ n26076;
  assign n26072 = n24318 ^ n24292;
  assign n26073 = n26072 ^ n25233;
  assign n26228 = n26077 ^ n26073;
  assign n26229 = n26078 & n26228;
  assign n26230 = n26229 ^ n26073;
  assign n26252 = n26234 ^ n26230;
  assign n26253 = ~n26251 & n26252;
  assign n26254 = n26253 ^ n26232;
  assign n26344 = n26258 ^ n26254;
  assign n26345 = n26343 & ~n26344;
  assign n26346 = n26345 ^ n26256;
  assign n26347 = n26346 ^ n26339;
  assign n26348 = ~n26342 & ~n26347;
  assign n26349 = n26348 ^ n26341;
  assign n26289 = n25727 ^ n25724;
  assign n26350 = n26349 ^ n26289;
  assign n26351 = n25543 ^ n25132;
  assign n26352 = n26351 ^ n24298;
  assign n26353 = n26352 ^ n26289;
  assign n26354 = ~n26350 & ~n26353;
  assign n26355 = n26354 ^ n26352;
  assign n26336 = n25156 ^ n24294;
  assign n26337 = n26336 ^ n25555;
  assign n26283 = n25730 ^ n25637;
  assign n26284 = n26283 ^ n25634;
  assign n26338 = n26337 ^ n26284;
  assign n26389 = n26355 ^ n26338;
  assign n26390 = n26389 ^ n23522;
  assign n26391 = n26352 ^ n26350;
  assign n26392 = n26391 ^ n23526;
  assign n26393 = n26346 ^ n26341;
  assign n26394 = n26393 ^ n26339;
  assign n26395 = n26394 ^ n23530;
  assign n26257 = n26256 ^ n26254;
  assign n26259 = n26258 ^ n26257;
  assign n26233 = n26232 ^ n26230;
  assign n26235 = n26234 ^ n26233;
  assign n26236 = n26235 ^ n23539;
  assign n26079 = n26078 ^ n26073;
  assign n26224 = n26079 ^ n23545;
  assign n26066 = n26065 ^ n26059;
  assign n26053 = n26052 ^ n26047;
  assign n25977 = n25976 ^ n25972;
  assign n25978 = n25977 ^ n23470;
  assign n25979 = n25969 ^ n25813;
  assign n25980 = n25979 ^ n23560;
  assign n25981 = n25966 ^ n25817;
  assign n25982 = n25981 ^ n23475;
  assign n26032 = n25963 ^ n25821;
  assign n25983 = n25960 ^ n25958;
  assign n25984 = n25983 ^ n23489;
  assign n25985 = n25952 ^ n25825;
  assign n25986 = n25985 ^ n23493;
  assign n26021 = n25949 ^ n25828;
  assign n25987 = n25946 ^ n25831;
  assign n25988 = n25987 ^ n25829;
  assign n25989 = n25988 ^ n23502;
  assign n25990 = n25943 ^ n25836;
  assign n25991 = n25990 ^ n23508;
  assign n25992 = n25940 ^ n25916;
  assign n25993 = n25992 ^ n25914;
  assign n25994 = n25993 ^ n23513;
  assign n25995 = n25937 ^ n25920;
  assign n25996 = n25995 ^ n25918;
  assign n25997 = n25996 ^ n23465;
  assign n25793 = n25792 ^ n25226;
  assign n25998 = n23308 & ~n25793;
  assign n25999 = n25998 ^ n23354;
  assign n26000 = n25927 ^ n25925;
  assign n26001 = n26000 ^ n25998;
  assign n26002 = n25999 & ~n26001;
  assign n26003 = n26002 ^ n23354;
  assign n26004 = n26003 ^ n23440;
  assign n26005 = n25934 ^ n25933;
  assign n26006 = n26005 ^ n26003;
  assign n26007 = ~n26004 & n26006;
  assign n26008 = n26007 ^ n23440;
  assign n26009 = n26008 ^ n25996;
  assign n26010 = n25997 & ~n26009;
  assign n26011 = n26010 ^ n23465;
  assign n26012 = n26011 ^ n25993;
  assign n26013 = ~n25994 & n26012;
  assign n26014 = n26013 ^ n23513;
  assign n26015 = n26014 ^ n25990;
  assign n26016 = ~n25991 & n26015;
  assign n26017 = n26016 ^ n23508;
  assign n26018 = n26017 ^ n25988;
  assign n26019 = ~n25989 & n26018;
  assign n26020 = n26019 ^ n23502;
  assign n26022 = n26021 ^ n26020;
  assign n26023 = n26021 ^ n23498;
  assign n26024 = n26022 & n26023;
  assign n26025 = n26024 ^ n23498;
  assign n26026 = n26025 ^ n25985;
  assign n26027 = n25986 & ~n26026;
  assign n26028 = n26027 ^ n23493;
  assign n26029 = n26028 ^ n25983;
  assign n26030 = n25984 & ~n26029;
  assign n26031 = n26030 ^ n23489;
  assign n26033 = n26032 ^ n26031;
  assign n26034 = n26032 ^ n23482;
  assign n26035 = n26033 & ~n26034;
  assign n26036 = n26035 ^ n23482;
  assign n26037 = n26036 ^ n25981;
  assign n26038 = ~n25982 & n26037;
  assign n26039 = n26038 ^ n23475;
  assign n26040 = n26039 ^ n25979;
  assign n26041 = n25980 & ~n26040;
  assign n26042 = n26041 ^ n23560;
  assign n26043 = n26042 ^ n25977;
  assign n26044 = n25978 & n26043;
  assign n26045 = n26044 ^ n23470;
  assign n26054 = n26053 ^ n26045;
  assign n26055 = n26053 ^ n23554;
  assign n26056 = ~n26054 & n26055;
  assign n26057 = n26056 ^ n23554;
  assign n26067 = n26066 ^ n26057;
  assign n26068 = n26066 ^ n23550;
  assign n26069 = n26067 & n26068;
  assign n26070 = n26069 ^ n23550;
  assign n26225 = n26079 ^ n26070;
  assign n26226 = n26224 & n26225;
  assign n26227 = n26226 ^ n23545;
  assign n26248 = n26235 ^ n26227;
  assign n26249 = n26236 & ~n26248;
  assign n26250 = n26249 ^ n23539;
  assign n26260 = n26259 ^ n26250;
  assign n26396 = n26259 ^ n23534;
  assign n26397 = n26260 & n26396;
  assign n26398 = n26397 ^ n23534;
  assign n26399 = n26398 ^ n26394;
  assign n26400 = n26395 & n26399;
  assign n26401 = n26400 ^ n23530;
  assign n26402 = n26401 ^ n26391;
  assign n26403 = ~n26392 & n26402;
  assign n26404 = n26403 ^ n23526;
  assign n26405 = n26404 ^ n26389;
  assign n26406 = n26390 & n26405;
  assign n26407 = n26406 ^ n23522;
  assign n26356 = n26355 ^ n26284;
  assign n26357 = n26338 & n26356;
  assign n26358 = n26357 ^ n26337;
  assign n26334 = n25738 ^ n25735;
  assign n26332 = n25197 ^ n24432;
  assign n26333 = n26332 ^ n25782;
  assign n26335 = n26334 ^ n26333;
  assign n26387 = n26358 ^ n26335;
  assign n26388 = n26387 ^ n23649;
  assign n26440 = n26407 ^ n26388;
  assign n26432 = n26401 ^ n23526;
  assign n26433 = n26432 ^ n26391;
  assign n26434 = n26398 ^ n26395;
  assign n26237 = n26236 ^ n26227;
  assign n26071 = n26070 ^ n23545;
  assign n26080 = n26079 ^ n26071;
  assign n26081 = n26067 ^ n23550;
  assign n26082 = n26054 ^ n23554;
  assign n26083 = n26042 ^ n23470;
  assign n26084 = n26083 ^ n25977;
  assign n26085 = n26039 ^ n23560;
  assign n26086 = n26085 ^ n25979;
  assign n26087 = n26036 ^ n25982;
  assign n26088 = n26033 ^ n23482;
  assign n26089 = n26022 ^ n23498;
  assign n26090 = n26017 ^ n23502;
  assign n26091 = n26090 ^ n25988;
  assign n26092 = n26014 ^ n23508;
  assign n26093 = n26092 ^ n25990;
  assign n25794 = n25793 ^ n23308;
  assign n26094 = n26000 ^ n25999;
  assign n26095 = ~n25794 & n26094;
  assign n26096 = n26005 ^ n26004;
  assign n26097 = n26095 & n26096;
  assign n26098 = n26008 ^ n25997;
  assign n26099 = n26097 & ~n26098;
  assign n26100 = n26011 ^ n23513;
  assign n26101 = n26100 ^ n25993;
  assign n26102 = n26099 & n26101;
  assign n26103 = ~n26093 & ~n26102;
  assign n26104 = n26091 & ~n26103;
  assign n26105 = n26089 & ~n26104;
  assign n26106 = n26025 ^ n25986;
  assign n26107 = n26105 & ~n26106;
  assign n26108 = n26028 ^ n25984;
  assign n26109 = n26107 & ~n26108;
  assign n26110 = ~n26088 & ~n26109;
  assign n26111 = n26087 & ~n26110;
  assign n26112 = n26086 & ~n26111;
  assign n26113 = ~n26084 & ~n26112;
  assign n26114 = n26082 & n26113;
  assign n26115 = n26081 & n26114;
  assign n26238 = ~n26080 & n26115;
  assign n26247 = ~n26237 & ~n26238;
  assign n26261 = n26260 ^ n23534;
  assign n26435 = n26247 & ~n26261;
  assign n26436 = ~n26434 & ~n26435;
  assign n26437 = ~n26433 & n26436;
  assign n26438 = n26404 ^ n26390;
  assign n26439 = ~n26437 & ~n26438;
  assign n26517 = n26440 ^ n26439;
  assign n26493 = n26438 ^ n26437;
  assign n922 = n848 ^ n807;
  assign n929 = n928 ^ n922;
  assign n930 = n929 ^ n912;
  assign n26494 = n26493 ^ n930;
  assign n26495 = n26436 ^ n26433;
  assign n26499 = n26498 ^ n26495;
  assign n26262 = n26261 ^ n26247;
  assign n26239 = n26238 ^ n26237;
  assign n26116 = n26115 ^ n26080;
  assign n26117 = n26116 ^ n626;
  assign n26213 = n26114 ^ n26081;
  assign n26118 = n26113 ^ n26082;
  assign n26122 = n26121 ^ n26118;
  assign n26123 = n26112 ^ n26084;
  assign n26127 = n26126 ^ n26123;
  assign n26199 = n26111 ^ n26086;
  assign n26128 = n26110 ^ n26087;
  assign n26129 = n26128 ^ n2207;
  assign n26130 = n26109 ^ n26088;
  assign n26131 = n26130 ^ n2064;
  assign n26132 = n26108 ^ n26107;
  assign n26133 = n26132 ^ n2046;
  assign n26185 = n26106 ^ n26105;
  assign n26135 = n24182 ^ n1864;
  assign n26136 = n26135 ^ n1694;
  assign n26137 = n26136 ^ n2029;
  assign n26134 = n26104 ^ n26089;
  assign n26138 = n26137 ^ n26134;
  assign n26139 = n26103 ^ n26091;
  assign n26143 = n26142 ^ n26139;
  assign n26144 = n26102 ^ n26093;
  assign n26145 = n26144 ^ n1629;
  assign n26146 = n26101 ^ n26099;
  assign n26150 = n26149 ^ n26146;
  assign n26160 = n26096 ^ n26095;
  assign n26151 = n25794 & n25797;
  assign n26155 = n26154 ^ n26151;
  assign n26156 = n26094 ^ n25794;
  assign n26157 = n26156 ^ n26154;
  assign n26158 = n26155 & n26157;
  assign n26159 = n26158 ^ n26151;
  assign n26161 = n26160 ^ n26159;
  assign n26162 = n24199 ^ n1472;
  assign n26163 = n26162 ^ n20796;
  assign n26164 = n26163 ^ n1493;
  assign n26165 = n26164 ^ n26159;
  assign n26166 = ~n26161 & n26165;
  assign n26167 = n26166 ^ n26164;
  assign n26168 = n26167 ^ n1532;
  assign n26169 = n26098 ^ n26097;
  assign n26170 = n26169 ^ n26167;
  assign n26171 = n26168 & n26170;
  assign n26172 = n26171 ^ n1532;
  assign n26173 = n26172 ^ n26146;
  assign n26174 = n26150 & ~n26173;
  assign n26175 = n26174 ^ n26149;
  assign n26176 = n26175 ^ n26144;
  assign n26177 = ~n26145 & n26176;
  assign n26178 = n26177 ^ n1629;
  assign n26179 = n26178 ^ n26139;
  assign n26180 = ~n26143 & n26179;
  assign n26181 = n26180 ^ n26142;
  assign n26182 = n26181 ^ n26134;
  assign n26183 = n26138 & ~n26182;
  assign n26184 = n26183 ^ n26137;
  assign n26186 = n26185 ^ n26184;
  assign n26187 = n26185 ^ n2034;
  assign n26188 = ~n26186 & n26187;
  assign n26189 = n26188 ^ n2034;
  assign n26190 = n26189 ^ n26132;
  assign n26191 = n26133 & ~n26190;
  assign n26192 = n26191 ^ n2046;
  assign n26193 = n26192 ^ n26130;
  assign n26194 = n26131 & ~n26193;
  assign n26195 = n26194 ^ n2064;
  assign n26196 = n26195 ^ n26128;
  assign n26197 = n26129 & ~n26196;
  assign n26198 = n26197 ^ n2207;
  assign n26200 = n26199 ^ n26198;
  assign n26204 = n26203 ^ n26199;
  assign n26205 = n26200 & ~n26204;
  assign n26206 = n26205 ^ n26203;
  assign n26207 = n26206 ^ n26123;
  assign n26208 = ~n26127 & n26207;
  assign n26209 = n26208 ^ n26126;
  assign n26210 = n26209 ^ n26118;
  assign n26211 = ~n26122 & n26210;
  assign n26212 = n26211 ^ n26121;
  assign n26214 = n26213 ^ n26212;
  assign n26215 = n24164 ^ n17451;
  assign n26216 = n26215 ^ n21195;
  assign n26217 = n26216 ^ n619;
  assign n26218 = n26217 ^ n26213;
  assign n26219 = n26214 & ~n26218;
  assign n26220 = n26219 ^ n26217;
  assign n26221 = n26220 ^ n26116;
  assign n26222 = n26117 & ~n26221;
  assign n26223 = n26222 ^ n626;
  assign n26240 = n26239 ^ n26223;
  assign n26241 = n24266 ^ n17444;
  assign n26242 = n26241 ^ n21143;
  assign n26243 = n26242 ^ n537;
  assign n26244 = n26243 ^ n26239;
  assign n26245 = ~n26240 & n26244;
  assign n26246 = n26245 ^ n26243;
  assign n26263 = n26262 ^ n26246;
  assign n26500 = n26262 ^ n25808;
  assign n26501 = n26263 & ~n26500;
  assign n26502 = n26501 ^ n25808;
  assign n26506 = n26505 ^ n26502;
  assign n26507 = n26435 ^ n26434;
  assign n26508 = n26507 ^ n26502;
  assign n26509 = n26506 & n26508;
  assign n26510 = n26509 ^ n26505;
  assign n26511 = n26510 ^ n26495;
  assign n26512 = n26499 & ~n26511;
  assign n26513 = n26512 ^ n26498;
  assign n26514 = n26513 ^ n26493;
  assign n26515 = n26494 & ~n26514;
  assign n26516 = n26515 ^ n930;
  assign n26518 = n26517 ^ n26516;
  assign n26519 = n26516 ^ n919;
  assign n26520 = n26518 & n26519;
  assign n26521 = n26520 ^ n919;
  assign n26359 = n26358 ^ n26334;
  assign n26360 = n26335 & ~n26359;
  assign n26361 = n26360 ^ n26333;
  assign n26329 = n25840 ^ n24497;
  assign n26330 = n26329 ^ n25302;
  assign n26411 = n26361 ^ n26330;
  assign n26278 = n25741 ^ n25633;
  assign n26412 = n26411 ^ n26278;
  assign n26408 = n26407 ^ n26387;
  assign n26409 = n26388 & n26408;
  assign n26410 = n26409 ^ n23649;
  assign n26413 = n26412 ^ n26410;
  assign n26442 = n26413 ^ n23755;
  assign n26441 = ~n26439 & ~n26440;
  assign n26491 = n26442 ^ n26441;
  assign n1059 = n1033 ^ n964;
  assign n1060 = n1059 ^ n939;
  assign n1061 = n1060 ^ n1049;
  assign n26492 = n26491 ^ n1061;
  assign n27135 = n26521 ^ n26492;
  assign n27132 = n25927 ^ n24628;
  assign n27133 = n27132 ^ n25345;
  assign n27106 = n26518 ^ n919;
  assign n27103 = n25213 ^ n24631;
  assign n27104 = n27103 ^ n25792;
  assign n27128 = n27106 ^ n27104;
  assign n26856 = n26513 ^ n930;
  assign n26857 = n26856 ^ n26493;
  assign n26582 = n25769 ^ n25615;
  assign n26853 = n26582 ^ n25166;
  assign n26854 = n26853 ^ n24643;
  assign n27099 = n26857 ^ n26854;
  assign n26717 = n26510 ^ n26498;
  assign n26718 = n26717 ^ n26495;
  assign n26715 = n25139 ^ n24637;
  assign n26559 = n25766 ^ n25617;
  assign n26716 = n26715 ^ n26559;
  assign n26719 = n26718 ^ n26716;
  assign n26707 = n26507 ^ n26505;
  assign n26708 = n26707 ^ n26502;
  assign n26264 = n26263 ^ n25808;
  assign n25804 = n25758 ^ n956;
  assign n25803 = n25802 ^ n25302;
  assign n25805 = n25804 ^ n25803;
  assign n26265 = n26264 ^ n25805;
  assign n26696 = n26243 ^ n26223;
  assign n26697 = n26696 ^ n26239;
  assign n26267 = n25750 ^ n25624;
  assign n26268 = n26267 ^ n25840;
  assign n26269 = n26268 ^ n25156;
  assign n26266 = n26220 ^ n26117;
  assign n26270 = n26269 ^ n26266;
  assign n26274 = n25744 ^ n25628;
  assign n26273 = n25555 ^ n24944;
  assign n26275 = n26274 ^ n26273;
  assign n26272 = n26209 ^ n26122;
  assign n26276 = n26275 ^ n26272;
  assign n26279 = n26278 ^ n25543;
  assign n26280 = n26279 ^ n24875;
  assign n26277 = n26206 ^ n26127;
  assign n26281 = n26280 ^ n26277;
  assign n26674 = n26203 ^ n26200;
  assign n26286 = n26195 ^ n26129;
  assign n26282 = n25413 ^ n24292;
  assign n26285 = n26284 ^ n26282;
  assign n26287 = n26286 ^ n26285;
  assign n26290 = n26289 ^ n25227;
  assign n26291 = n26290 ^ n24302;
  assign n26288 = n26192 ^ n26131;
  assign n26292 = n26291 ^ n26288;
  assign n26660 = n26189 ^ n2046;
  assign n26661 = n26660 ^ n26132;
  assign n26652 = n26184 ^ n2034;
  assign n26653 = n26652 ^ n26185;
  assign n26295 = n26181 ^ n26138;
  assign n26293 = n26234 ^ n24310;
  assign n26294 = n26293 ^ n25241;
  assign n26296 = n26295 ^ n26294;
  assign n26642 = n26178 ^ n26143;
  assign n26299 = n26175 ^ n1629;
  assign n26300 = n26299 ^ n26144;
  assign n26297 = n26064 ^ n24707;
  assign n26298 = n26297 ^ n25248;
  assign n26301 = n26300 ^ n26298;
  assign n26303 = n26051 ^ n25252;
  assign n26304 = n26303 ^ n24700;
  assign n26302 = n26172 ^ n26150;
  assign n26305 = n26304 ^ n26302;
  assign n26308 = n25975 ^ n25256;
  assign n26309 = n26308 ^ n24322;
  assign n26306 = n26169 ^ n1532;
  assign n26307 = n26306 ^ n26167;
  assign n26310 = n26309 ^ n26307;
  assign n26312 = n25262 ^ n24329;
  assign n26313 = n26312 ^ n25810;
  assign n26311 = n26164 ^ n26161;
  assign n26314 = n26313 ^ n26311;
  assign n26316 = n25814 ^ n25265;
  assign n26317 = n26316 ^ n24330;
  assign n26315 = n26156 ^ n26155;
  assign n26318 = n26317 ^ n26315;
  assign n26319 = n25818 ^ n24336;
  assign n26320 = n26319 ^ n25269;
  assign n25798 = n25797 ^ n25794;
  assign n26321 = n26320 ^ n25798;
  assign n26593 = n25957 ^ n24340;
  assign n26594 = n26593 ^ n25273;
  assign n26580 = n24351 ^ n23512;
  assign n26581 = n26580 ^ n25337;
  assign n26583 = n26582 ^ n26581;
  assign n26557 = n24355 ^ n23517;
  assign n26558 = n26557 ^ n25345;
  assign n26560 = n26559 ^ n26558;
  assign n26473 = n25763 ^ n1372;
  assign n26471 = n24623 ^ n23947;
  assign n26472 = n26471 ^ n25213;
  assign n26474 = n26473 ^ n26472;
  assign n26457 = n25166 ^ n24628;
  assign n26458 = n26457 ^ n23969;
  assign n26459 = n26458 ^ n25804;
  assign n26380 = n25753 ^ n25622;
  assign n26377 = n24631 ^ n23962;
  assign n26378 = n26377 ^ n25139;
  assign n26453 = n26380 ^ n26378;
  assign n26322 = n24643 ^ n23958;
  assign n26323 = n26322 ^ n25907;
  assign n26324 = n26323 ^ n26267;
  assign n26327 = n25747 ^ n25626;
  assign n26325 = n24637 ^ n23955;
  assign n26326 = n26325 ^ n25802;
  assign n26328 = n26327 ^ n26326;
  assign n26331 = n26330 ^ n26278;
  assign n26362 = n26361 ^ n26278;
  assign n26363 = n26331 & ~n26362;
  assign n26364 = n26363 ^ n26330;
  assign n26365 = n26364 ^ n26274;
  assign n26366 = n25856 ^ n24616;
  assign n26367 = n26366 ^ n25325;
  assign n26368 = n26367 ^ n26274;
  assign n26369 = ~n26365 & ~n26368;
  assign n26370 = n26369 ^ n26367;
  assign n26371 = n26370 ^ n26326;
  assign n26372 = n26328 & ~n26371;
  assign n26373 = n26372 ^ n26327;
  assign n26374 = n26373 ^ n26323;
  assign n26375 = ~n26324 & ~n26374;
  assign n26376 = n26375 ^ n26373;
  assign n26454 = n26380 ^ n26376;
  assign n26455 = n26453 & n26454;
  assign n26456 = n26455 ^ n26378;
  assign n26468 = n26458 ^ n26456;
  assign n26469 = n26459 & ~n26468;
  assign n26470 = n26469 ^ n25804;
  assign n26554 = n26473 ^ n26470;
  assign n26555 = n26474 & ~n26554;
  assign n26556 = n26555 ^ n26472;
  assign n26577 = n26559 ^ n26556;
  assign n26578 = n26560 & n26577;
  assign n26579 = n26578 ^ n26558;
  assign n26584 = n26583 ^ n26579;
  assign n26561 = n26560 ^ n26556;
  assign n26562 = n26561 ^ n22538;
  assign n26475 = n26474 ^ n26470;
  assign n26550 = n26475 ^ n23287;
  assign n26460 = n26459 ^ n26456;
  assign n26463 = n26460 ^ n23241;
  assign n26379 = n26378 ^ n26376;
  assign n26381 = n26380 ^ n26379;
  assign n26382 = n26381 ^ n23243;
  assign n26383 = n26373 ^ n26324;
  assign n26384 = n26383 ^ n23254;
  assign n26385 = n26370 ^ n26328;
  assign n26386 = n26385 ^ n23249;
  assign n26417 = n26367 ^ n26365;
  assign n26414 = n26412 ^ n23755;
  assign n26415 = ~n26413 & ~n26414;
  assign n26416 = n26415 ^ n23755;
  assign n26418 = n26417 ^ n26416;
  assign n26419 = n26417 ^ n23938;
  assign n26420 = ~n26418 & ~n26419;
  assign n26421 = n26420 ^ n23938;
  assign n26422 = n26421 ^ n26385;
  assign n26423 = n26386 & n26422;
  assign n26424 = n26423 ^ n23249;
  assign n26425 = n26424 ^ n26383;
  assign n26426 = n26384 & ~n26425;
  assign n26427 = n26426 ^ n23254;
  assign n26449 = n26427 ^ n26381;
  assign n26450 = ~n26382 & ~n26449;
  assign n26451 = n26450 ^ n23243;
  assign n26464 = n26460 ^ n26451;
  assign n26465 = ~n26463 & ~n26464;
  assign n26466 = n26465 ^ n23241;
  assign n26551 = n26475 ^ n26466;
  assign n26552 = ~n26550 & n26551;
  assign n26553 = n26552 ^ n23287;
  assign n26574 = n26561 ^ n26553;
  assign n26575 = ~n26562 & n26574;
  assign n26576 = n26575 ^ n22538;
  assign n26585 = n26584 ^ n26576;
  assign n26586 = n26585 ^ n23300;
  assign n26563 = n26562 ^ n26553;
  assign n26428 = n26427 ^ n26382;
  assign n26429 = n26424 ^ n23254;
  assign n26430 = n26429 ^ n26383;
  assign n26431 = n26421 ^ n26386;
  assign n26443 = n26441 & ~n26442;
  assign n26444 = n26418 ^ n23938;
  assign n26445 = ~n26443 & ~n26444;
  assign n26446 = n26431 & ~n26445;
  assign n26447 = ~n26430 & n26446;
  assign n26448 = n26428 & n26447;
  assign n26452 = n26451 ^ n23241;
  assign n26461 = n26460 ^ n26452;
  assign n26462 = ~n26448 & n26461;
  assign n26467 = n26466 ^ n23287;
  assign n26476 = n26475 ^ n26467;
  assign n26564 = ~n26462 & n26476;
  assign n26573 = n26563 & n26564;
  assign n26587 = n26586 ^ n26573;
  assign n26591 = n26590 ^ n26587;
  assign n26565 = n26564 ^ n26563;
  assign n26478 = n24538 ^ n2515;
  assign n26479 = n26478 ^ n2363;
  assign n26480 = n26479 ^ n1541;
  assign n26477 = n26476 ^ n26462;
  assign n26481 = n26480 ^ n26477;
  assign n26539 = n26461 ^ n26448;
  assign n26482 = n26447 ^ n26428;
  assign n2277 = n2276 ^ n1316;
  assign n2278 = n2277 ^ n2273;
  assign n2282 = n2281 ^ n2278;
  assign n26483 = n26482 ^ n2282;
  assign n26485 = n24550 ^ n17431;
  assign n26486 = n26485 ^ n1228;
  assign n26487 = n26486 ^ n2271;
  assign n26484 = n26446 ^ n26430;
  assign n26488 = n26487 ^ n26484;
  assign n26489 = n26444 ^ n26443;
  assign n1045 = n1042 ^ n976;
  assign n1052 = n1051 ^ n1045;
  assign n1056 = n1055 ^ n1052;
  assign n26490 = n26489 ^ n1056;
  assign n26522 = n26521 ^ n26491;
  assign n26523 = n26492 & ~n26522;
  assign n26524 = n26523 ^ n1061;
  assign n26525 = n26524 ^ n26489;
  assign n26526 = n26490 & ~n26525;
  assign n26527 = n26526 ^ n1056;
  assign n1216 = n1209 ^ n1125;
  assign n1220 = n1219 ^ n1216;
  assign n1224 = n1223 ^ n1220;
  assign n26528 = n26527 ^ n1224;
  assign n26529 = n26445 ^ n26431;
  assign n26530 = n26529 ^ n26527;
  assign n26531 = n26528 & ~n26530;
  assign n26532 = n26531 ^ n1224;
  assign n26533 = n26532 ^ n26484;
  assign n26534 = n26488 & ~n26533;
  assign n26535 = n26534 ^ n26487;
  assign n26536 = n26535 ^ n26482;
  assign n26537 = ~n26483 & n26536;
  assign n26538 = n26537 ^ n2282;
  assign n26540 = n26539 ^ n26538;
  assign n26541 = n24543 ^ n2508;
  assign n26542 = n26541 ^ n21278;
  assign n26543 = n26542 ^ n2351;
  assign n26544 = n26543 ^ n26539;
  assign n26545 = n26540 & ~n26544;
  assign n26546 = n26545 ^ n26543;
  assign n26547 = n26546 ^ n26477;
  assign n26548 = n26481 & ~n26547;
  assign n26549 = n26548 ^ n26480;
  assign n26566 = n26565 ^ n26549;
  assign n26567 = n2598 ^ n2530;
  assign n26568 = n26567 ^ n21328;
  assign n26569 = n26568 ^ n2489;
  assign n26570 = n26569 ^ n26565;
  assign n26571 = n26566 & ~n26570;
  assign n26572 = n26571 ^ n26569;
  assign n26592 = n26591 ^ n26572;
  assign n26595 = n26594 ^ n26592;
  assign n26614 = n25822 ^ n24675;
  assign n26615 = n26614 ^ n25277;
  assign n26607 = n26546 ^ n26481;
  assign n26598 = n26535 ^ n26483;
  assign n26599 = n25833 ^ n25222;
  assign n26600 = n26599 ^ n24350;
  assign n26601 = ~n26598 & ~n26600;
  assign n26596 = n25829 ^ n24346;
  assign n26597 = n26596 ^ n25283;
  assign n26602 = n26601 ^ n26597;
  assign n26603 = n26543 ^ n26540;
  assign n26604 = n26603 ^ n26597;
  assign n26605 = ~n26602 & ~n26604;
  assign n26606 = n26605 ^ n26601;
  assign n26608 = n26607 ^ n26606;
  assign n26609 = n25220 ^ n24342;
  assign n26610 = n26609 ^ n25278;
  assign n26611 = n26610 ^ n26607;
  assign n26612 = ~n26608 & n26611;
  assign n26613 = n26612 ^ n26610;
  assign n26616 = n26615 ^ n26613;
  assign n26617 = n26569 ^ n26566;
  assign n26618 = n26617 ^ n26613;
  assign n26619 = ~n26616 & n26618;
  assign n26620 = n26619 ^ n26615;
  assign n26621 = n26620 ^ n26592;
  assign n26622 = ~n26595 & ~n26621;
  assign n26623 = n26622 ^ n26594;
  assign n26624 = n26623 ^ n25798;
  assign n26625 = n26321 & ~n26624;
  assign n26626 = n26625 ^ n26320;
  assign n26627 = n26626 ^ n26315;
  assign n26628 = ~n26318 & n26627;
  assign n26629 = n26628 ^ n26317;
  assign n26630 = n26629 ^ n26311;
  assign n26631 = n26314 & ~n26630;
  assign n26632 = n26631 ^ n26313;
  assign n26633 = n26632 ^ n26307;
  assign n26634 = ~n26310 & n26633;
  assign n26635 = n26634 ^ n26309;
  assign n26636 = n26635 ^ n26302;
  assign n26637 = ~n26305 & ~n26636;
  assign n26638 = n26637 ^ n26304;
  assign n26639 = n26638 ^ n26300;
  assign n26640 = n26301 & ~n26639;
  assign n26641 = n26640 ^ n26298;
  assign n26643 = n26642 ^ n26641;
  assign n26644 = n26077 ^ n25244;
  assign n26645 = n26644 ^ n24316;
  assign n26646 = n26645 ^ n26642;
  assign n26647 = ~n26643 & n26646;
  assign n26648 = n26647 ^ n26645;
  assign n26649 = n26648 ^ n26295;
  assign n26650 = n26296 & n26649;
  assign n26651 = n26650 ^ n26294;
  assign n26654 = n26653 ^ n26651;
  assign n26655 = n26258 ^ n25237;
  assign n26656 = n26655 ^ n24309;
  assign n26657 = n26656 ^ n26653;
  assign n26658 = ~n26654 & n26657;
  assign n26659 = n26658 ^ n26656;
  assign n26662 = n26661 ^ n26659;
  assign n26663 = n26339 ^ n25233;
  assign n26664 = n26663 ^ n24307;
  assign n26665 = n26664 ^ n26661;
  assign n26666 = ~n26662 & ~n26665;
  assign n26667 = n26666 ^ n26664;
  assign n26668 = n26667 ^ n26288;
  assign n26669 = ~n26292 & n26668;
  assign n26670 = n26669 ^ n26291;
  assign n26671 = n26670 ^ n26285;
  assign n26672 = n26287 & n26671;
  assign n26673 = n26672 ^ n26286;
  assign n26675 = n26674 ^ n26673;
  assign n26676 = n26334 ^ n25529;
  assign n26677 = n26676 ^ n24739;
  assign n26678 = n26677 ^ n26674;
  assign n26679 = n26675 & ~n26678;
  assign n26680 = n26679 ^ n26677;
  assign n26681 = n26680 ^ n26277;
  assign n26682 = ~n26281 & n26681;
  assign n26683 = n26682 ^ n26280;
  assign n26684 = n26683 ^ n26272;
  assign n26685 = ~n26276 & n26684;
  assign n26686 = n26685 ^ n26275;
  assign n26271 = n26217 ^ n26214;
  assign n26687 = n26686 ^ n26271;
  assign n26688 = n26327 ^ n25782;
  assign n26689 = n26688 ^ n25132;
  assign n26690 = n26689 ^ n26271;
  assign n26691 = n26687 & ~n26690;
  assign n26692 = n26691 ^ n26689;
  assign n26693 = n26692 ^ n26269;
  assign n26694 = ~n26270 & n26693;
  assign n26695 = n26694 ^ n26266;
  assign n26698 = n26697 ^ n26695;
  assign n26699 = n26380 ^ n25197;
  assign n26700 = n26699 ^ n25856;
  assign n26701 = n26700 ^ n26697;
  assign n26702 = ~n26698 & ~n26701;
  assign n26703 = n26702 ^ n26700;
  assign n26704 = n26703 ^ n26264;
  assign n26705 = ~n26265 & ~n26704;
  assign n26706 = n26705 ^ n25805;
  assign n26709 = n26708 ^ n26706;
  assign n26710 = n25907 ^ n25325;
  assign n26711 = n26710 ^ n26473;
  assign n26712 = n26711 ^ n26708;
  assign n26713 = n26709 & ~n26712;
  assign n26714 = n26713 ^ n26711;
  assign n26850 = n26716 ^ n26714;
  assign n26851 = ~n26719 & n26850;
  assign n26852 = n26851 ^ n26718;
  assign n27100 = n26857 ^ n26852;
  assign n27101 = ~n27099 & ~n27100;
  assign n27102 = n27101 ^ n26854;
  assign n27129 = n27106 ^ n27102;
  assign n27130 = ~n27128 & ~n27129;
  assign n27131 = n27130 ^ n27104;
  assign n27134 = n27133 ^ n27131;
  assign n27136 = n27135 ^ n27134;
  assign n27179 = n27136 ^ n23969;
  assign n27105 = n27104 ^ n27102;
  assign n27107 = n27106 ^ n27105;
  assign n27108 = n27107 ^ n23962;
  assign n26855 = n26854 ^ n26852;
  assign n26858 = n26857 ^ n26855;
  assign n26859 = n26858 ^ n23958;
  assign n26720 = n26719 ^ n26714;
  assign n26721 = n26720 ^ n23955;
  assign n26722 = n26711 ^ n26709;
  assign n26723 = n26722 ^ n24616;
  assign n26724 = n26703 ^ n26265;
  assign n26725 = n26724 ^ n24497;
  assign n26726 = n26700 ^ n26698;
  assign n26727 = n26726 ^ n24432;
  assign n26728 = n26692 ^ n26270;
  assign n26729 = n26728 ^ n24294;
  assign n26730 = n26689 ^ n26687;
  assign n26731 = n26730 ^ n24298;
  assign n26732 = n26683 ^ n26276;
  assign n26733 = n26732 ^ n24304;
  assign n26734 = n26680 ^ n26281;
  assign n26735 = n26734 ^ n24369;
  assign n26736 = n26677 ^ n26675;
  assign n26737 = n26736 ^ n24311;
  assign n26738 = n26670 ^ n26287;
  assign n26739 = n26738 ^ n24318;
  assign n26740 = n26667 ^ n26292;
  assign n26741 = n26740 ^ n24374;
  assign n26812 = n26664 ^ n26662;
  assign n26742 = n26656 ^ n26654;
  assign n26743 = n26742 ^ n24324;
  assign n26744 = n26648 ^ n26294;
  assign n26745 = n26744 ^ n26295;
  assign n26746 = n26745 ^ n24381;
  assign n26747 = n26645 ^ n26643;
  assign n26748 = n26747 ^ n24282;
  assign n26797 = n26638 ^ n26298;
  assign n26798 = n26797 ^ n26300;
  assign n26792 = n26635 ^ n26305;
  assign n26749 = n26632 ^ n26309;
  assign n26750 = n26749 ^ n26307;
  assign n26751 = n26750 ^ n23469;
  assign n26752 = n26629 ^ n26314;
  assign n26753 = n26752 ^ n23474;
  assign n26754 = n26626 ^ n26318;
  assign n26755 = n26754 ^ n23478;
  assign n26756 = n26623 ^ n26321;
  assign n26757 = n26756 ^ n23481;
  assign n26758 = n26620 ^ n26595;
  assign n26759 = n26758 ^ n23486;
  assign n26760 = n26617 ^ n26616;
  assign n26761 = n26760 ^ n23492;
  assign n26762 = n26610 ^ n26608;
  assign n26763 = n26762 ^ n23497;
  assign n26764 = n26600 ^ n26598;
  assign n26765 = ~n23507 & n26764;
  assign n26766 = n26765 ^ n23505;
  assign n26767 = n26603 ^ n26602;
  assign n26768 = n26767 ^ n26765;
  assign n26769 = n26766 & ~n26768;
  assign n26770 = n26769 ^ n23505;
  assign n26771 = n26770 ^ n26762;
  assign n26772 = n26763 & ~n26771;
  assign n26773 = n26772 ^ n23497;
  assign n26774 = n26773 ^ n26760;
  assign n26775 = n26761 & ~n26774;
  assign n26776 = n26775 ^ n23492;
  assign n26777 = n26776 ^ n26758;
  assign n26778 = ~n26759 & ~n26777;
  assign n26779 = n26778 ^ n23486;
  assign n26780 = n26779 ^ n26756;
  assign n26781 = n26757 & n26780;
  assign n26782 = n26781 ^ n23481;
  assign n26783 = n26782 ^ n26754;
  assign n26784 = n26755 & n26783;
  assign n26785 = n26784 ^ n23478;
  assign n26786 = n26785 ^ n26752;
  assign n26787 = ~n26753 & n26786;
  assign n26788 = n26787 ^ n23474;
  assign n26789 = n26788 ^ n26750;
  assign n26790 = ~n26751 & ~n26789;
  assign n26791 = n26790 ^ n23469;
  assign n26793 = n26792 ^ n26791;
  assign n26794 = n26792 ^ n24018;
  assign n26795 = n26793 & n26794;
  assign n26796 = n26795 ^ n24018;
  assign n26799 = n26798 ^ n26796;
  assign n26800 = n26798 ^ n24111;
  assign n26801 = ~n26799 & n26800;
  assign n26802 = n26801 ^ n24111;
  assign n26803 = n26802 ^ n26747;
  assign n26804 = ~n26748 & ~n26803;
  assign n26805 = n26804 ^ n24282;
  assign n26806 = n26805 ^ n26745;
  assign n26807 = ~n26746 & n26806;
  assign n26808 = n26807 ^ n24381;
  assign n26809 = n26808 ^ n26742;
  assign n26810 = ~n26743 & ~n26809;
  assign n26811 = n26810 ^ n24324;
  assign n26813 = n26812 ^ n26811;
  assign n26814 = n26812 ^ n24378;
  assign n26815 = ~n26813 & n26814;
  assign n26816 = n26815 ^ n24378;
  assign n26817 = n26816 ^ n26740;
  assign n26818 = n26741 & n26817;
  assign n26819 = n26818 ^ n24374;
  assign n26820 = n26819 ^ n26738;
  assign n26821 = ~n26739 & n26820;
  assign n26822 = n26821 ^ n24318;
  assign n26823 = n26822 ^ n26736;
  assign n26824 = n26737 & n26823;
  assign n26825 = n26824 ^ n24311;
  assign n26826 = n26825 ^ n26734;
  assign n26827 = n26735 & ~n26826;
  assign n26828 = n26827 ^ n24369;
  assign n26829 = n26828 ^ n26732;
  assign n26830 = ~n26733 & ~n26829;
  assign n26831 = n26830 ^ n24304;
  assign n26832 = n26831 ^ n26730;
  assign n26833 = ~n26731 & n26832;
  assign n26834 = n26833 ^ n24298;
  assign n26835 = n26834 ^ n26728;
  assign n26836 = ~n26729 & n26835;
  assign n26837 = n26836 ^ n24294;
  assign n26838 = n26837 ^ n26726;
  assign n26839 = ~n26727 & n26838;
  assign n26840 = n26839 ^ n24432;
  assign n26841 = n26840 ^ n26724;
  assign n26842 = n26725 & ~n26841;
  assign n26843 = n26842 ^ n24497;
  assign n26844 = n26843 ^ n26722;
  assign n26845 = ~n26723 & n26844;
  assign n26846 = n26845 ^ n24616;
  assign n26847 = n26846 ^ n26720;
  assign n26848 = n26721 & n26847;
  assign n26849 = n26848 ^ n23955;
  assign n27096 = n26858 ^ n26849;
  assign n27097 = n26859 & ~n27096;
  assign n27098 = n27097 ^ n23958;
  assign n27124 = n27107 ^ n27098;
  assign n27125 = ~n27108 & n27124;
  assign n27126 = n27125 ^ n23962;
  assign n27180 = n27136 ^ n27126;
  assign n27181 = n27179 & ~n27180;
  assign n27182 = n27181 ^ n23969;
  assign n27174 = n25337 ^ n24623;
  assign n27175 = n27174 ^ n25934;
  assign n27173 = n26524 ^ n26490;
  assign n27176 = n27175 ^ n27173;
  assign n27169 = n27135 ^ n27133;
  assign n27170 = n27135 ^ n27131;
  assign n27171 = ~n27169 & ~n27170;
  assign n27172 = n27171 ^ n27133;
  assign n27177 = n27176 ^ n27172;
  assign n27178 = n27177 ^ n23947;
  assign n27183 = n27182 ^ n27178;
  assign n27127 = n27126 ^ n23969;
  assign n27137 = n27136 ^ n27127;
  assign n27109 = n27108 ^ n27098;
  assign n26860 = n26859 ^ n26849;
  assign n26861 = n26846 ^ n26721;
  assign n26862 = n26843 ^ n26723;
  assign n26863 = n26840 ^ n26725;
  assign n26864 = n26831 ^ n26731;
  assign n26865 = n26825 ^ n26735;
  assign n26866 = n26813 ^ n24378;
  assign n26867 = n26808 ^ n26743;
  assign n26868 = n26793 ^ n24018;
  assign n26869 = n26776 ^ n26759;
  assign n26870 = n26773 ^ n26761;
  assign n26871 = n26764 ^ n23507;
  assign n26872 = n26767 ^ n26766;
  assign n26873 = ~n26871 & n26872;
  assign n26874 = n26770 ^ n26763;
  assign n26875 = n26873 & n26874;
  assign n26876 = n26870 & n26875;
  assign n26877 = ~n26869 & n26876;
  assign n26878 = n26779 ^ n23481;
  assign n26879 = n26878 ^ n26756;
  assign n26880 = ~n26877 & n26879;
  assign n26881 = n26782 ^ n26755;
  assign n26882 = ~n26880 & n26881;
  assign n26883 = n26785 ^ n26753;
  assign n26884 = ~n26882 & ~n26883;
  assign n26885 = n26788 ^ n26751;
  assign n26886 = n26884 & ~n26885;
  assign n26887 = ~n26868 & n26886;
  assign n26888 = n26799 ^ n24111;
  assign n26889 = ~n26887 & ~n26888;
  assign n26890 = n26802 ^ n24282;
  assign n26891 = n26890 ^ n26747;
  assign n26892 = ~n26889 & ~n26891;
  assign n26893 = n26805 ^ n26746;
  assign n26894 = ~n26892 & ~n26893;
  assign n26895 = n26867 & ~n26894;
  assign n26896 = n26866 & n26895;
  assign n26897 = n26816 ^ n26741;
  assign n26898 = n26896 & n26897;
  assign n26899 = n26819 ^ n26739;
  assign n26900 = n26898 & n26899;
  assign n26901 = n26822 ^ n26737;
  assign n26902 = ~n26900 & n26901;
  assign n26903 = ~n26865 & n26902;
  assign n26904 = n26828 ^ n26733;
  assign n26905 = ~n26903 & ~n26904;
  assign n26906 = n26864 & n26905;
  assign n26907 = n26834 ^ n26729;
  assign n26908 = ~n26906 & ~n26907;
  assign n26909 = n26837 ^ n26727;
  assign n26910 = ~n26908 & n26909;
  assign n26911 = ~n26863 & n26910;
  assign n26912 = ~n26862 & ~n26911;
  assign n26913 = ~n26861 & ~n26912;
  assign n27110 = n26860 & n26913;
  assign n27138 = ~n27109 & n27110;
  assign n27168 = ~n27137 & ~n27138;
  assign n27184 = n27183 ^ n27168;
  assign n27139 = n27138 ^ n27137;
  assign n27140 = n27139 ^ n2344;
  assign n27111 = n27110 ^ n27109;
  assign n26914 = n26913 ^ n26860;
  assign n1347 = n1328 ^ n1244;
  assign n1348 = n1347 ^ n1344;
  assign n1352 = n1351 ^ n1348;
  assign n26915 = n26914 ^ n1352;
  assign n27088 = n26912 ^ n26861;
  assign n26916 = n26911 ^ n26862;
  assign n26917 = n26916 ^ n1179;
  assign n27080 = n26910 ^ n26863;
  assign n27072 = n26909 ^ n26908;
  assign n27064 = n26907 ^ n26906;
  assign n26918 = n26905 ^ n26864;
  assign n26919 = n26918 ^ n725;
  assign n27053 = n25080 ^ n18107;
  assign n27054 = n27053 ^ n679;
  assign n27055 = n27054 ^ n717;
  assign n26920 = n26902 ^ n26865;
  assign n664 = n657 ^ n549;
  assign n671 = n670 ^ n664;
  assign n675 = n674 ^ n671;
  assign n26921 = n26920 ^ n675;
  assign n26922 = n26901 ^ n26900;
  assign n26926 = n26925 ^ n26922;
  assign n26927 = n26899 ^ n26898;
  assign n26931 = n26930 ^ n26927;
  assign n27036 = n26897 ^ n26896;
  assign n26932 = n26895 ^ n26866;
  assign n26936 = n26935 ^ n26932;
  assign n26937 = n26894 ^ n26867;
  assign n26941 = n26940 ^ n26937;
  assign n26942 = n26893 ^ n26892;
  assign n26946 = n26945 ^ n26942;
  assign n26947 = n26891 ^ n26889;
  assign n26951 = n26950 ^ n26947;
  assign n26952 = n26888 ^ n26887;
  assign n26956 = n26955 ^ n26952;
  assign n27016 = n26886 ^ n26868;
  assign n27008 = n26885 ^ n26884;
  assign n26998 = n26881 ^ n26880;
  assign n26993 = n26879 ^ n26877;
  assign n26985 = n26876 ^ n26869;
  assign n26960 = n26874 ^ n26873;
  assign n26964 = n26963 ^ n26960;
  assign n26965 = n25336 ^ n18239;
  assign n26966 = n26965 ^ n1550;
  assign n26967 = n26966 ^ n2642;
  assign n26968 = n26871 & n26967;
  assign n26972 = n26971 ^ n26968;
  assign n26973 = n26872 ^ n26871;
  assign n26974 = n26973 ^ n26968;
  assign n26975 = n26972 & n26974;
  assign n26976 = n26975 ^ n26971;
  assign n26977 = n26976 ^ n26960;
  assign n26978 = n26964 & ~n26977;
  assign n26979 = n26978 ^ n26963;
  assign n26980 = n26979 ^ n26959;
  assign n26981 = n26875 ^ n26870;
  assign n26982 = n26981 ^ n26979;
  assign n26983 = n26980 & ~n26982;
  assign n26984 = n26983 ^ n26959;
  assign n26986 = n26985 ^ n26984;
  assign n26990 = n26989 ^ n26985;
  assign n26991 = n26986 & ~n26990;
  assign n26992 = n26991 ^ n26989;
  assign n26994 = n26993 ^ n26992;
  assign n26995 = n26993 ^ n1672;
  assign n26996 = ~n26994 & n26995;
  assign n26997 = n26996 ^ n1672;
  assign n26999 = n26998 ^ n26997;
  assign n27000 = n26998 ^ n1684;
  assign n27001 = n26999 & ~n27000;
  assign n27002 = n27001 ^ n1684;
  assign n1762 = n1754 ^ n1704;
  assign n1766 = n1765 ^ n1762;
  assign n1770 = n1769 ^ n1766;
  assign n27003 = n27002 ^ n1770;
  assign n27004 = n26883 ^ n26882;
  assign n27005 = n27004 ^ n27002;
  assign n27006 = n27003 & n27005;
  assign n27007 = n27006 ^ n1770;
  assign n27009 = n27008 ^ n27007;
  assign n27013 = n27012 ^ n27007;
  assign n27014 = ~n27009 & n27013;
  assign n27015 = n27014 ^ n27012;
  assign n27017 = n27016 ^ n27015;
  assign n27018 = n27016 ^ n1910;
  assign n27019 = ~n27017 & n27018;
  assign n27020 = n27019 ^ n1910;
  assign n27021 = n27020 ^ n26952;
  assign n27022 = n26956 & ~n27021;
  assign n27023 = n27022 ^ n26955;
  assign n27024 = n27023 ^ n26947;
  assign n27025 = ~n26951 & n27024;
  assign n27026 = n27025 ^ n26950;
  assign n27027 = n27026 ^ n26942;
  assign n27028 = n26946 & ~n27027;
  assign n27029 = n27028 ^ n26945;
  assign n27030 = n27029 ^ n26937;
  assign n27031 = n26941 & ~n27030;
  assign n27032 = n27031 ^ n26940;
  assign n27033 = n27032 ^ n26932;
  assign n27034 = ~n26936 & n27033;
  assign n27035 = n27034 ^ n26935;
  assign n27037 = n27036 ^ n27035;
  assign n27041 = n27040 ^ n27035;
  assign n27042 = n27037 & n27041;
  assign n27043 = n27042 ^ n27040;
  assign n27044 = n27043 ^ n26927;
  assign n27045 = ~n26931 & n27044;
  assign n27046 = n27045 ^ n26930;
  assign n27047 = n27046 ^ n26922;
  assign n27048 = ~n26926 & n27047;
  assign n27049 = n27048 ^ n26925;
  assign n27050 = n27049 ^ n26920;
  assign n27051 = ~n26921 & n27050;
  assign n27052 = n27051 ^ n675;
  assign n27056 = n27055 ^ n27052;
  assign n27057 = n26904 ^ n26903;
  assign n27058 = n27057 ^ n27052;
  assign n27059 = n27056 & n27058;
  assign n27060 = n27059 ^ n27055;
  assign n27061 = n27060 ^ n26918;
  assign n27062 = ~n26919 & n27061;
  assign n27063 = n27062 ^ n725;
  assign n27065 = n27064 ^ n27063;
  assign n27069 = n27068 ^ n27064;
  assign n27070 = ~n27065 & n27069;
  assign n27071 = n27070 ^ n27068;
  assign n27073 = n27072 ^ n27071;
  assign n27077 = n27076 ^ n27071;
  assign n27078 = ~n27073 & n27077;
  assign n27079 = n27078 ^ n27076;
  assign n27081 = n27080 ^ n27079;
  assign n27082 = n27079 ^ n1167;
  assign n27083 = ~n27081 & n27082;
  assign n27084 = n27083 ^ n1167;
  assign n27085 = n27084 ^ n26916;
  assign n27086 = n26917 & ~n27085;
  assign n27087 = n27086 ^ n1179;
  assign n27089 = n27088 ^ n27087;
  assign n1192 = n1152 ^ n1106;
  assign n1193 = n1192 ^ n1186;
  assign n1197 = n1196 ^ n1193;
  assign n27090 = n27088 ^ n1197;
  assign n27091 = n27089 & ~n27090;
  assign n27092 = n27091 ^ n1197;
  assign n27093 = n27092 ^ n26914;
  assign n27094 = ~n26915 & n27093;
  assign n27095 = n27094 ^ n1352;
  assign n27112 = n27111 ^ n27095;
  assign n2327 = n2306 ^ n2300;
  assign n2328 = n2327 ^ n1359;
  assign n2332 = n2331 ^ n2328;
  assign n27121 = n27095 ^ n2332;
  assign n27122 = ~n27112 & n27121;
  assign n27123 = n27122 ^ n2332;
  assign n27165 = n27139 ^ n27123;
  assign n27166 = n27140 & ~n27165;
  assign n27167 = n27166 ^ n2344;
  assign n27185 = n27184 ^ n27167;
  assign n2421 = n2420 ^ n2357;
  assign n2422 = n2421 ^ n2417;
  assign n2423 = n2422 ^ n2409;
  assign n27186 = n27185 ^ n2423;
  assign n25223 = n25222 ^ n25220;
  assign n25799 = n25798 ^ n25220;
  assign n25800 = ~n25223 & ~n25799;
  assign n25801 = n25800 ^ n25222;
  assign n27113 = n27112 ^ n2332;
  assign n27146 = ~n25801 & n27113;
  assign n27142 = n25822 ^ n25283;
  assign n27143 = n26315 ^ n25822;
  assign n27144 = n27142 & n27143;
  assign n27145 = n27144 ^ n25283;
  assign n27147 = n27146 ^ n27145;
  assign n27141 = n27140 ^ n27123;
  assign n27162 = n27145 ^ n27141;
  assign n27163 = n27147 & ~n27162;
  assign n27164 = n27163 ^ n27146;
  assign n27187 = n27186 ^ n27164;
  assign n27158 = n25957 ^ n25278;
  assign n27159 = n26311 ^ n25957;
  assign n27160 = ~n27158 & ~n27159;
  assign n27161 = n27160 ^ n25278;
  assign n27188 = n27187 ^ n27161;
  assign n27114 = n27113 ^ n25801;
  assign n27149 = ~n24350 & ~n27114;
  assign n27150 = n27149 ^ n24346;
  assign n27148 = n27147 ^ n27141;
  assign n27155 = n27149 ^ n27148;
  assign n27156 = n27150 & ~n27155;
  assign n27157 = n27156 ^ n24346;
  assign n27189 = n27188 ^ n27157;
  assign n27190 = n27189 ^ n24342;
  assign n27230 = n25211 ^ n1544;
  assign n27231 = n27230 ^ n2411;
  assign n27232 = n27231 ^ n2566;
  assign n27223 = n27175 ^ n27172;
  assign n27224 = n27176 & n27223;
  assign n27225 = n27224 ^ n27173;
  assign n27220 = n25918 ^ n24355;
  assign n27221 = n27220 ^ n25224;
  assign n27218 = n26529 ^ n1224;
  assign n27219 = n27218 ^ n26527;
  assign n27222 = n27221 ^ n27219;
  assign n27226 = n27225 ^ n27222;
  assign n27213 = n27182 ^ n23947;
  assign n27214 = n27182 ^ n27177;
  assign n27215 = ~n27213 & ~n27214;
  assign n27216 = n27215 ^ n23947;
  assign n27217 = n27216 ^ n23517;
  assign n27227 = n27226 ^ n27217;
  assign n27212 = ~n27168 & ~n27183;
  assign n27228 = n27227 ^ n27212;
  assign n27209 = n27167 ^ n2423;
  assign n27210 = n27185 & n27209;
  assign n27211 = n27210 ^ n2423;
  assign n27229 = n27228 ^ n27211;
  assign n27233 = n27232 ^ n27229;
  assign n27204 = n25818 ^ n25277;
  assign n27205 = n26307 ^ n25818;
  assign n27206 = n27204 & ~n27205;
  assign n27207 = n27206 ^ n25277;
  assign n27201 = n27186 ^ n27161;
  assign n27202 = n27187 & n27201;
  assign n27203 = n27202 ^ n27161;
  assign n27208 = n27207 ^ n27203;
  assign n27234 = n27233 ^ n27208;
  assign n27235 = n27234 ^ n24675;
  assign n27198 = n27188 ^ n24342;
  assign n27199 = ~n27189 & ~n27198;
  assign n27200 = n27199 ^ n24342;
  assign n27236 = n27235 ^ n27200;
  assign n27280 = n27190 & ~n27236;
  assign n27268 = n27212 & n27227;
  assign n27269 = n27268 ^ n25914;
  assign n2562 = n2561 ^ n2492;
  assign n2569 = n2568 ^ n2562;
  assign n2570 = n2569 ^ n1517;
  assign n27270 = n27269 ^ n2570;
  assign n27271 = n27270 ^ n26580;
  assign n27272 = n27271 ^ n25355;
  assign n27267 = n26532 ^ n26488;
  assign n27273 = n27272 ^ n27267;
  assign n27263 = n27226 ^ n23517;
  assign n27264 = n27226 ^ n27216;
  assign n27265 = ~n27263 & ~n27264;
  assign n27266 = n27265 ^ n23517;
  assign n27274 = n27273 ^ n27266;
  assign n27260 = n27232 ^ n27228;
  assign n27261 = n27229 & ~n27260;
  assign n27262 = n27261 ^ n27232;
  assign n27275 = n27274 ^ n27262;
  assign n27257 = n27225 ^ n27219;
  assign n27258 = n27222 & ~n27257;
  assign n27259 = n27258 ^ n27221;
  assign n27276 = n27275 ^ n27259;
  assign n27253 = n25814 ^ n25273;
  assign n27254 = n26302 ^ n25814;
  assign n27255 = ~n27253 & ~n27254;
  assign n27256 = n27255 ^ n25273;
  assign n27277 = n27276 ^ n27256;
  assign n27249 = n27233 ^ n27207;
  assign n27250 = n27233 ^ n27203;
  assign n27251 = n27249 & ~n27250;
  assign n27252 = n27251 ^ n27207;
  assign n27278 = n27277 ^ n27252;
  assign n27245 = n27234 ^ n27200;
  assign n27246 = ~n27235 & ~n27245;
  assign n27247 = n27246 ^ n24675;
  assign n27248 = n27247 ^ n24340;
  assign n27279 = n27278 ^ n27248;
  assign n27281 = n27280 ^ n27279;
  assign n27285 = n27284 ^ n27281;
  assign n27237 = n27236 ^ n27190;
  assign n27238 = n27237 ^ n27197;
  assign n1557 = n1556 ^ n1433;
  assign n1558 = n1557 ^ n1526;
  assign n1559 = n1558 ^ n1472;
  assign n27191 = n27190 ^ n1559;
  assign n27117 = n18359 ^ n2654;
  assign n27118 = n27117 ^ n22392;
  assign n27119 = n27118 ^ n1502;
  assign n27115 = n27114 ^ n24350;
  assign n27116 = n2636 & n27115;
  assign n27120 = n27119 ^ n27116;
  assign n27151 = n27150 ^ n27148;
  assign n27152 = n27151 ^ n27116;
  assign n27153 = n27120 & ~n27152;
  assign n27154 = n27153 ^ n27119;
  assign n27239 = n27154 ^ n1559;
  assign n27240 = n27191 & ~n27239;
  assign n27241 = n27240 ^ n27190;
  assign n27242 = n27241 ^ n27237;
  assign n27243 = n27238 & ~n27242;
  assign n27244 = n27243 ^ n27197;
  assign n27627 = n27281 ^ n27244;
  assign n27628 = n27285 & ~n27627;
  assign n27629 = n27628 ^ n27284;
  assign n27452 = n27278 ^ n24340;
  assign n27453 = n27278 ^ n27247;
  assign n27454 = n27452 & n27453;
  assign n27455 = n27454 ^ n24340;
  assign n27353 = n25810 ^ n25269;
  assign n27354 = n26300 ^ n25810;
  assign n27355 = n27353 & n27354;
  assign n27356 = n27355 ^ n25269;
  assign n27351 = n26967 ^ n26871;
  assign n27348 = n27256 ^ n27252;
  assign n27349 = n27277 & ~n27348;
  assign n27350 = n27349 ^ n27276;
  assign n27352 = n27351 ^ n27350;
  assign n27450 = n27356 ^ n27352;
  assign n27451 = n27450 ^ n24336;
  assign n27543 = n27455 ^ n27451;
  assign n27542 = ~n27279 & n27280;
  assign n27622 = n27543 ^ n27542;
  assign n27626 = n27625 ^ n27622;
  assign n27821 = n27629 ^ n27626;
  assign n27817 = n26674 ^ n26234;
  assign n27399 = n27020 ^ n26956;
  assign n27818 = n27399 ^ n26674;
  assign n27819 = n27817 & n27818;
  assign n27820 = n27819 ^ n26234;
  assign n27822 = n27821 ^ n27820;
  assign n27823 = n26286 ^ n26077;
  assign n27304 = n27017 ^ n1910;
  assign n27824 = n27304 ^ n26286;
  assign n27825 = n27823 & ~n27824;
  assign n27826 = n27825 ^ n26077;
  assign n27286 = n27285 ^ n27244;
  assign n27827 = n27826 ^ n27286;
  assign n28102 = n27241 ^ n27238;
  assign n27828 = n26661 ^ n26051;
  assign n27316 = n27004 ^ n1770;
  assign n27317 = n27316 ^ n27002;
  assign n27829 = n27317 ^ n26661;
  assign n27830 = ~n27828 & n27829;
  assign n27831 = n27830 ^ n26051;
  assign n27192 = n27191 ^ n27154;
  assign n27832 = n27831 ^ n27192;
  assign n27834 = n26653 ^ n25975;
  assign n27193 = n26999 ^ n1684;
  assign n27835 = n27193 ^ n26653;
  assign n27836 = ~n27834 & n27835;
  assign n27837 = n27836 ^ n25975;
  assign n27833 = n27151 ^ n27120;
  assign n27838 = n27837 ^ n27833;
  assign n28087 = n27115 ^ n2636;
  assign n28045 = n26642 ^ n25814;
  assign n27374 = n26989 ^ n26984;
  assign n27375 = n27374 ^ n26985;
  assign n28046 = n27375 ^ n26642;
  assign n28047 = ~n28045 & ~n28046;
  assign n28048 = n28047 ^ n25814;
  assign n28040 = n2646 ^ n2576;
  assign n28041 = n28040 ^ n2539;
  assign n28042 = n28041 ^ n2632;
  assign n27928 = n25914 ^ n25337;
  assign n27929 = n26607 ^ n25914;
  assign n27930 = n27928 & n27929;
  assign n27931 = n27930 ^ n25337;
  assign n27734 = n27084 ^ n1179;
  assign n27735 = n27734 ^ n26916;
  assign n27932 = n27931 ^ n27735;
  assign n27883 = n25918 ^ n25345;
  assign n27884 = n26603 ^ n25918;
  assign n27885 = ~n27883 & ~n27884;
  assign n27886 = n27885 ^ n25345;
  assign n27742 = n27081 ^ n1167;
  assign n27924 = n27886 ^ n27742;
  assign n27839 = n25934 ^ n25213;
  assign n27840 = n26598 ^ n25934;
  assign n27841 = n27839 & ~n27840;
  assign n27842 = n27841 ^ n25213;
  assign n27752 = n27076 ^ n27073;
  assign n27843 = n27842 ^ n27752;
  assign n27844 = n25927 ^ n25166;
  assign n27845 = n27267 ^ n25927;
  assign n27846 = ~n27844 & ~n27845;
  assign n27847 = n27846 ^ n25166;
  assign n27758 = n27068 ^ n27065;
  assign n27848 = n27847 ^ n27758;
  assign n27868 = n27060 ^ n26919;
  assign n27849 = n26582 ^ n25907;
  assign n27850 = n27173 ^ n26582;
  assign n27851 = n27849 & ~n27850;
  assign n27852 = n27851 ^ n25907;
  assign n27765 = n27057 ^ n27056;
  assign n27853 = n27852 ^ n27765;
  assign n27854 = n26559 ^ n25802;
  assign n27855 = n27135 ^ n26559;
  assign n27856 = n27854 & ~n27855;
  assign n27857 = n27856 ^ n25802;
  assign n27772 = n27049 ^ n26921;
  assign n27858 = n27857 ^ n27772;
  assign n27700 = n26473 ^ n25856;
  assign n27701 = n27106 ^ n26473;
  assign n27702 = n27700 & ~n27701;
  assign n27703 = n27702 ^ n25856;
  assign n27698 = n27046 ^ n26925;
  assign n27699 = n27698 ^ n26922;
  assign n27704 = n27703 ^ n27699;
  assign n27530 = n27043 ^ n26930;
  assign n27531 = n27530 ^ n26927;
  assign n27525 = n25840 ^ n25804;
  assign n27526 = n26857 ^ n25804;
  assign n27527 = ~n27525 & n27526;
  assign n27528 = n27527 ^ n25840;
  assign n27694 = n27531 ^ n27528;
  assign n27431 = n26380 ^ n25782;
  assign n27432 = n26718 ^ n26380;
  assign n27433 = ~n27431 & n27432;
  assign n27434 = n27433 ^ n25782;
  assign n27430 = n27040 ^ n27037;
  assign n27435 = n27434 ^ n27430;
  assign n27291 = n26267 ^ n25555;
  assign n27292 = n26708 ^ n26267;
  assign n27293 = n27291 & ~n27292;
  assign n27294 = n27293 ^ n25555;
  assign n27290 = n27032 ^ n26936;
  assign n27295 = n27294 ^ n27290;
  assign n27297 = n26327 ^ n25543;
  assign n27298 = n26327 ^ n26264;
  assign n27299 = n27297 & n27298;
  assign n27300 = n27299 ^ n25543;
  assign n27296 = n27029 ^ n26941;
  assign n27301 = n27300 ^ n27296;
  assign n27305 = n26284 ^ n25233;
  assign n27306 = n26284 ^ n26272;
  assign n27307 = n27305 & ~n27306;
  assign n27308 = n27307 ^ n25233;
  assign n27309 = n27308 ^ n27304;
  assign n27314 = n27012 ^ n27009;
  assign n27310 = n26289 ^ n25237;
  assign n27311 = n26289 ^ n26277;
  assign n27312 = ~n27310 & ~n27311;
  assign n27313 = n27312 ^ n25237;
  assign n27315 = n27314 ^ n27313;
  assign n27318 = n26339 ^ n25241;
  assign n27319 = n26674 ^ n26339;
  assign n27320 = ~n27318 & n27319;
  assign n27321 = n27320 ^ n25241;
  assign n27322 = n27321 ^ n27317;
  assign n27323 = n26258 ^ n25244;
  assign n27324 = n26286 ^ n26258;
  assign n27325 = ~n27323 & ~n27324;
  assign n27326 = n27325 ^ n25244;
  assign n27327 = n27326 ^ n27193;
  assign n27332 = n26994 ^ n1672;
  assign n27328 = n26234 ^ n25248;
  assign n27329 = n26288 ^ n26234;
  assign n27330 = n27328 & n27329;
  assign n27331 = n27330 ^ n25248;
  assign n27333 = n27332 ^ n27331;
  assign n27337 = n26051 ^ n25262;
  assign n27338 = n26295 ^ n26051;
  assign n27339 = ~n27337 & n27338;
  assign n27340 = n27339 ^ n25262;
  assign n27335 = n26976 ^ n26963;
  assign n27336 = n27335 ^ n26960;
  assign n27341 = n27340 ^ n27336;
  assign n27346 = n26973 ^ n26972;
  assign n27342 = n25975 ^ n25265;
  assign n27343 = n26642 ^ n25975;
  assign n27344 = n27342 & ~n27343;
  assign n27345 = n27344 ^ n25265;
  assign n27347 = n27346 ^ n27345;
  assign n27357 = n27356 ^ n27351;
  assign n27358 = n27352 & n27357;
  assign n27359 = n27358 ^ n27356;
  assign n27360 = n27359 ^ n27345;
  assign n27361 = n27347 & n27360;
  assign n27362 = n27361 ^ n27346;
  assign n27363 = n27362 ^ n27340;
  assign n27364 = n27341 & n27363;
  assign n27365 = n27364 ^ n27336;
  assign n27334 = n26981 ^ n26980;
  assign n27366 = n27365 ^ n27334;
  assign n27367 = n26064 ^ n25256;
  assign n27368 = n26653 ^ n26064;
  assign n27369 = ~n27367 & n27368;
  assign n27370 = n27369 ^ n25256;
  assign n27371 = n27370 ^ n27365;
  assign n27372 = n27366 & ~n27371;
  assign n27373 = n27372 ^ n27334;
  assign n27376 = n27375 ^ n27373;
  assign n27377 = n26077 ^ n25252;
  assign n27378 = n26661 ^ n26077;
  assign n27379 = ~n27377 & ~n27378;
  assign n27380 = n27379 ^ n25252;
  assign n27381 = n27380 ^ n27375;
  assign n27382 = n27376 & n27381;
  assign n27383 = n27382 ^ n27380;
  assign n27384 = n27383 ^ n27331;
  assign n27385 = ~n27333 & ~n27384;
  assign n27386 = n27385 ^ n27332;
  assign n27387 = n27386 ^ n27193;
  assign n27388 = n27327 & n27387;
  assign n27389 = n27388 ^ n27326;
  assign n27390 = n27389 ^ n27317;
  assign n27391 = n27322 & ~n27390;
  assign n27392 = n27391 ^ n27321;
  assign n27393 = n27392 ^ n27314;
  assign n27394 = n27315 & n27393;
  assign n27395 = n27394 ^ n27313;
  assign n27396 = n27395 ^ n27304;
  assign n27397 = ~n27309 & ~n27396;
  assign n27398 = n27397 ^ n27308;
  assign n27400 = n27399 ^ n27398;
  assign n27401 = n26334 ^ n25227;
  assign n27402 = n26334 ^ n26271;
  assign n27403 = n27401 & ~n27402;
  assign n27404 = n27403 ^ n25227;
  assign n27405 = n27404 ^ n27399;
  assign n27406 = n27400 & ~n27405;
  assign n27407 = n27406 ^ n27404;
  assign n27303 = n27023 ^ n26951;
  assign n27408 = n27407 ^ n27303;
  assign n27409 = n26278 ^ n25413;
  assign n27410 = n26278 ^ n26266;
  assign n27411 = ~n27409 & n27410;
  assign n27412 = n27411 ^ n25413;
  assign n27413 = n27412 ^ n27303;
  assign n27414 = ~n27408 & ~n27413;
  assign n27415 = n27414 ^ n27412;
  assign n27302 = n27026 ^ n26946;
  assign n27416 = n27415 ^ n27302;
  assign n27417 = n26274 ^ n25529;
  assign n27418 = n26697 ^ n26274;
  assign n27419 = n27417 & n27418;
  assign n27420 = n27419 ^ n25529;
  assign n27421 = n27420 ^ n27302;
  assign n27422 = ~n27416 & ~n27421;
  assign n27423 = n27422 ^ n27420;
  assign n27424 = n27423 ^ n27296;
  assign n27425 = n27301 & n27424;
  assign n27426 = n27425 ^ n27300;
  assign n27427 = n27426 ^ n27290;
  assign n27428 = n27295 & n27427;
  assign n27429 = n27428 ^ n27294;
  assign n27522 = n27430 ^ n27429;
  assign n27523 = ~n27435 & ~n27522;
  assign n27524 = n27523 ^ n27434;
  assign n27695 = n27531 ^ n27524;
  assign n27696 = ~n27694 & n27695;
  assign n27697 = n27696 ^ n27528;
  assign n27859 = n27703 ^ n27697;
  assign n27860 = n27704 & n27859;
  assign n27861 = n27860 ^ n27699;
  assign n27862 = n27861 ^ n27772;
  assign n27863 = ~n27858 & ~n27862;
  assign n27864 = n27863 ^ n27857;
  assign n27865 = n27864 ^ n27765;
  assign n27866 = ~n27853 & n27865;
  assign n27867 = n27866 ^ n27852;
  assign n27869 = n27868 ^ n27867;
  assign n27870 = n25792 ^ n25139;
  assign n27871 = n27219 ^ n25792;
  assign n27872 = ~n27870 & n27871;
  assign n27873 = n27872 ^ n25139;
  assign n27874 = n27873 ^ n27868;
  assign n27875 = n27869 & ~n27874;
  assign n27876 = n27875 ^ n27873;
  assign n27877 = n27876 ^ n27758;
  assign n27878 = ~n27848 & ~n27877;
  assign n27879 = n27878 ^ n27847;
  assign n27880 = n27879 ^ n27752;
  assign n27881 = ~n27843 & n27880;
  assign n27882 = n27881 ^ n27842;
  assign n27925 = n27882 ^ n27742;
  assign n27926 = n27924 & n27925;
  assign n27927 = n27926 ^ n27886;
  assign n27933 = n27932 ^ n27927;
  assign n27887 = n27886 ^ n27882;
  assign n27888 = n27887 ^ n27742;
  assign n27889 = n27888 ^ n24628;
  assign n27890 = n27879 ^ n27842;
  assign n27891 = n27890 ^ n27752;
  assign n27892 = n27891 ^ n24631;
  assign n27893 = n27876 ^ n27848;
  assign n27894 = n27893 ^ n24643;
  assign n27895 = n27873 ^ n27869;
  assign n27896 = n27895 ^ n24637;
  assign n27899 = n27861 ^ n27857;
  assign n27900 = n27899 ^ n27772;
  assign n27901 = n27900 ^ n25302;
  assign n27705 = n27704 ^ n27697;
  assign n27706 = n27705 ^ n25197;
  assign n27529 = n27528 ^ n27524;
  assign n27532 = n27531 ^ n27529;
  assign n27533 = n27532 ^ n25156;
  assign n27436 = n27435 ^ n27429;
  assign n27437 = n27436 ^ n25132;
  assign n27514 = n27426 ^ n27295;
  assign n27508 = n27423 ^ n27300;
  assign n27509 = n27508 ^ n27296;
  assign n27503 = n27420 ^ n27416;
  assign n27438 = n27412 ^ n27408;
  assign n27439 = n27438 ^ n24292;
  assign n27495 = n27404 ^ n27400;
  assign n27440 = n27395 ^ n27309;
  assign n27441 = n27440 ^ n24307;
  assign n27442 = n27392 ^ n27315;
  assign n27443 = n27442 ^ n24309;
  assign n27444 = n27386 ^ n27327;
  assign n27445 = n27444 ^ n24316;
  assign n27446 = n27380 ^ n27376;
  assign n27447 = n27446 ^ n24700;
  assign n27462 = n27362 ^ n27341;
  assign n27448 = n27359 ^ n27347;
  assign n27449 = n27448 ^ n24330;
  assign n27456 = n27455 ^ n27450;
  assign n27457 = n27451 & ~n27456;
  assign n27458 = n27457 ^ n24336;
  assign n27459 = n27458 ^ n27448;
  assign n27460 = ~n27449 & n27459;
  assign n27461 = n27460 ^ n24330;
  assign n27463 = n27462 ^ n27461;
  assign n27464 = n27462 ^ n24329;
  assign n27465 = ~n27463 & ~n27464;
  assign n27466 = n27465 ^ n24329;
  assign n27467 = n27466 ^ n24322;
  assign n27468 = n27370 ^ n27334;
  assign n27469 = n27468 ^ n27365;
  assign n27470 = n27469 ^ n27466;
  assign n27471 = ~n27467 & ~n27470;
  assign n27472 = n27471 ^ n24322;
  assign n27473 = n27472 ^ n27446;
  assign n27474 = ~n27447 & n27473;
  assign n27475 = n27474 ^ n24700;
  assign n27476 = n27475 ^ n24707;
  assign n27477 = n27383 ^ n27333;
  assign n27478 = n27477 ^ n27475;
  assign n27479 = n27476 & n27478;
  assign n27480 = n27479 ^ n24707;
  assign n27481 = n27480 ^ n27444;
  assign n27482 = n27445 & n27481;
  assign n27483 = n27482 ^ n24316;
  assign n27484 = n27483 ^ n24310;
  assign n27485 = n27389 ^ n27322;
  assign n27486 = n27485 ^ n27483;
  assign n27487 = n27484 & n27486;
  assign n27488 = n27487 ^ n24310;
  assign n27489 = n27488 ^ n27442;
  assign n27490 = ~n27443 & n27489;
  assign n27491 = n27490 ^ n24309;
  assign n27492 = n27491 ^ n27440;
  assign n27493 = ~n27441 & n27492;
  assign n27494 = n27493 ^ n24307;
  assign n27496 = n27495 ^ n27494;
  assign n27497 = n27495 ^ n24302;
  assign n27498 = ~n27496 & ~n27497;
  assign n27499 = n27498 ^ n24302;
  assign n27500 = n27499 ^ n27438;
  assign n27501 = ~n27439 & n27500;
  assign n27502 = n27501 ^ n24292;
  assign n27504 = n27503 ^ n27502;
  assign n27505 = n27503 ^ n24739;
  assign n27506 = ~n27504 & ~n27505;
  assign n27507 = n27506 ^ n24739;
  assign n27510 = n27509 ^ n27507;
  assign n27511 = n27509 ^ n24875;
  assign n27512 = n27510 & n27511;
  assign n27513 = n27512 ^ n24875;
  assign n27515 = n27514 ^ n27513;
  assign n27516 = n27514 ^ n24944;
  assign n27517 = n27515 & n27516;
  assign n27518 = n27517 ^ n24944;
  assign n27519 = n27518 ^ n27436;
  assign n27520 = n27437 & ~n27519;
  assign n27521 = n27520 ^ n25132;
  assign n27691 = n27532 ^ n27521;
  assign n27692 = ~n27533 & n27691;
  assign n27693 = n27692 ^ n25156;
  assign n27902 = n27705 ^ n27693;
  assign n27903 = ~n27706 & ~n27902;
  assign n27904 = n27903 ^ n25197;
  assign n27905 = n27904 ^ n27900;
  assign n27906 = ~n27901 & n27905;
  assign n27907 = n27906 ^ n25302;
  assign n27897 = n27864 ^ n27852;
  assign n27898 = n27897 ^ n27765;
  assign n27908 = n27907 ^ n27898;
  assign n27909 = n27898 ^ n25325;
  assign n27910 = ~n27908 & n27909;
  assign n27911 = n27910 ^ n25325;
  assign n27912 = n27911 ^ n27895;
  assign n27913 = n27896 & ~n27912;
  assign n27914 = n27913 ^ n24637;
  assign n27915 = n27914 ^ n27893;
  assign n27916 = ~n27894 & ~n27915;
  assign n27917 = n27916 ^ n24643;
  assign n27918 = n27917 ^ n27891;
  assign n27919 = n27892 & ~n27918;
  assign n27920 = n27919 ^ n24631;
  assign n27921 = n27920 ^ n27888;
  assign n27922 = n27889 & n27921;
  assign n27923 = n27922 ^ n24628;
  assign n27934 = n27933 ^ n27923;
  assign n27935 = n27934 ^ n24623;
  assign n27936 = n27920 ^ n24628;
  assign n27937 = n27936 ^ n27888;
  assign n27938 = n27904 ^ n25302;
  assign n27939 = n27938 ^ n27900;
  assign n27534 = n27533 ^ n27521;
  assign n27535 = n27515 ^ n24944;
  assign n27536 = n27488 ^ n27443;
  assign n27537 = n27477 ^ n24707;
  assign n27538 = n27537 ^ n27475;
  assign n27539 = n27469 ^ n27467;
  assign n27540 = n27463 ^ n24329;
  assign n27541 = n27458 ^ n27449;
  assign n27544 = ~n27542 & ~n27543;
  assign n27545 = ~n27541 & ~n27544;
  assign n27546 = ~n27540 & n27545;
  assign n27547 = ~n27539 & ~n27546;
  assign n27548 = n27472 ^ n27447;
  assign n27549 = n27547 & n27548;
  assign n27550 = ~n27538 & ~n27549;
  assign n27551 = n27480 ^ n27445;
  assign n27552 = n27550 & n27551;
  assign n27553 = n27485 ^ n24310;
  assign n27554 = n27553 ^ n27483;
  assign n27555 = n27552 & n27554;
  assign n27556 = n27536 & n27555;
  assign n27557 = n27491 ^ n27441;
  assign n27558 = ~n27556 & ~n27557;
  assign n27559 = n27496 ^ n24302;
  assign n27560 = ~n27558 & n27559;
  assign n27561 = n27499 ^ n24292;
  assign n27562 = n27561 ^ n27438;
  assign n27563 = n27560 & ~n27562;
  assign n27564 = n27504 ^ n24739;
  assign n27565 = n27563 & ~n27564;
  assign n27566 = n27510 ^ n24875;
  assign n27567 = ~n27565 & n27566;
  assign n27568 = n27535 & ~n27567;
  assign n27569 = n27518 ^ n25132;
  assign n27570 = n27569 ^ n27436;
  assign n27571 = n27568 & ~n27570;
  assign n27690 = ~n27534 & ~n27571;
  assign n27707 = n27706 ^ n27693;
  assign n27940 = n27690 & ~n27707;
  assign n27941 = n27939 & n27940;
  assign n27942 = n27908 ^ n25325;
  assign n27943 = ~n27941 & n27942;
  assign n27944 = n27911 ^ n27896;
  assign n27945 = n27943 & n27944;
  assign n27946 = n27914 ^ n27894;
  assign n27947 = n27945 & ~n27946;
  assign n27948 = n27917 ^ n27892;
  assign n27949 = n27947 & ~n27948;
  assign n27950 = n27937 & ~n27949;
  assign n27951 = n27935 & n27950;
  assign n27960 = n27927 ^ n27735;
  assign n27961 = ~n27932 & ~n27960;
  assign n27962 = n27961 ^ n27931;
  assign n27955 = n25833 ^ n25224;
  assign n27956 = n26617 ^ n25833;
  assign n27957 = ~n27955 & ~n27956;
  assign n27958 = n27957 ^ n25224;
  assign n27726 = n27087 ^ n1197;
  assign n27727 = n27726 ^ n27088;
  assign n27959 = n27958 ^ n27727;
  assign n27963 = n27962 ^ n27959;
  assign n27964 = n27963 ^ n24355;
  assign n27952 = n27933 ^ n24623;
  assign n27953 = ~n27934 & ~n27952;
  assign n27954 = n27953 ^ n24623;
  assign n27965 = n27964 ^ n27954;
  assign n28038 = n27951 & ~n27965;
  assign n28030 = n25829 ^ n25355;
  assign n28031 = n26592 ^ n25829;
  assign n28032 = ~n28030 & ~n28031;
  assign n28033 = n28032 ^ n25355;
  assign n28027 = n27962 ^ n27727;
  assign n28028 = ~n27959 & ~n28027;
  assign n28029 = n28028 ^ n27958;
  assign n28034 = n28033 ^ n28029;
  assign n27719 = n27092 ^ n1352;
  assign n27720 = n27719 ^ n26914;
  assign n28035 = n28034 ^ n27720;
  assign n28036 = n28035 ^ n24351;
  assign n28024 = n27963 ^ n27954;
  assign n28025 = ~n27964 & ~n28024;
  assign n28026 = n28025 ^ n24355;
  assign n28037 = n28036 ^ n28026;
  assign n28039 = n28038 ^ n28037;
  assign n28043 = n28042 ^ n28039;
  assign n27966 = n27965 ^ n27951;
  assign n27967 = n27966 ^ n2531;
  assign n27968 = n27950 ^ n27935;
  assign n2505 = n2457 ^ n2401;
  assign n2512 = n2511 ^ n2505;
  assign n2516 = n2515 ^ n2512;
  assign n27969 = n27968 ^ n2516;
  assign n27971 = n25775 ^ n2388;
  assign n27972 = n27971 ^ n22528;
  assign n27973 = n27972 ^ n2508;
  assign n27970 = n27949 ^ n27937;
  assign n27974 = n27973 ^ n27970;
  assign n28007 = n27948 ^ n27947;
  assign n27976 = n1381 ^ n1298;
  assign n27977 = n27976 ^ n1214;
  assign n27978 = n27977 ^ n17431;
  assign n27975 = n27946 ^ n27945;
  assign n27979 = n27978 ^ n27975;
  assign n27981 = n1372 ^ n1280;
  assign n27982 = n27981 ^ n22354;
  assign n27983 = n27982 ^ n1209;
  assign n27980 = n27944 ^ n27943;
  assign n27984 = n27983 ^ n27980;
  assign n27985 = n27942 ^ n27941;
  assign n27986 = n27985 ^ n1043;
  assign n27987 = n27940 ^ n27939;
  assign n27991 = n27990 ^ n27987;
  assign n27708 = n27707 ^ n27690;
  assign n27709 = n27708 ^ n887;
  assign n27572 = n27571 ^ n27534;
  assign n803 = n772 ^ n738;
  assign n804 = n803 ^ n800;
  assign n808 = n807 ^ n804;
  assign n27573 = n27572 ^ n808;
  assign n27574 = n27570 ^ n27568;
  assign n776 = n763 ^ n749;
  assign n789 = n788 ^ n776;
  assign n793 = n792 ^ n789;
  assign n27575 = n27574 ^ n793;
  assign n27576 = n27567 ^ n27535;
  assign n27580 = n27579 ^ n27576;
  assign n27582 = n25738 ^ n689;
  assign n27583 = n27582 ^ n22363;
  assign n27584 = n27583 ^ n17538;
  assign n27581 = n27566 ^ n27565;
  assign n27585 = n27584 ^ n27581;
  assign n27586 = n27564 ^ n27563;
  assign n27590 = n27589 ^ n27586;
  assign n27592 = n25727 ^ n18689;
  assign n27593 = n27592 ^ n22463;
  assign n27594 = n27593 ^ n524;
  assign n27591 = n27562 ^ n27560;
  assign n27595 = n27594 ^ n27591;
  assign n27597 = n25719 ^ n18694;
  assign n27598 = n27597 ^ n605;
  assign n27599 = n27598 ^ n17451;
  assign n27596 = n27559 ^ n27558;
  assign n27600 = n27599 ^ n27596;
  assign n27661 = n27557 ^ n27556;
  assign n27601 = n27555 ^ n27536;
  assign n27605 = n27604 ^ n27601;
  assign n27606 = n27554 ^ n27552;
  assign n27610 = n27609 ^ n27606;
  assign n27650 = n27551 ^ n27550;
  assign n27611 = n27549 ^ n27538;
  assign n27612 = n27611 ^ n2020;
  assign n27613 = n27546 ^ n27539;
  assign n27614 = n27613 ^ n1880;
  assign n27615 = n27545 ^ n27540;
  assign n1851 = n1790 ^ n1743;
  assign n1861 = n1860 ^ n1851;
  assign n1865 = n1864 ^ n1861;
  assign n27616 = n27615 ^ n1865;
  assign n27620 = n27544 ^ n27541;
  assign n27621 = n27620 ^ n27619;
  assign n27630 = n27629 ^ n27622;
  assign n27631 = n27626 & ~n27630;
  assign n27632 = n27631 ^ n27625;
  assign n27633 = n27632 ^ n27620;
  assign n27634 = ~n27621 & n27633;
  assign n27635 = n27634 ^ n27619;
  assign n27636 = n27635 ^ n27615;
  assign n27637 = n27616 & ~n27636;
  assign n27638 = n27637 ^ n1865;
  assign n27639 = n27638 ^ n27613;
  assign n27640 = n27614 & ~n27639;
  assign n27641 = n27640 ^ n1880;
  assign n27642 = n27641 ^ n2005;
  assign n27643 = n27548 ^ n27547;
  assign n27644 = n27643 ^ n27641;
  assign n27645 = n27642 & ~n27644;
  assign n27646 = n27645 ^ n2005;
  assign n27647 = n27646 ^ n27611;
  assign n27648 = ~n27612 & n27647;
  assign n27649 = n27648 ^ n2020;
  assign n27651 = n27650 ^ n27649;
  assign n27652 = n27649 ^ n2190;
  assign n27653 = n27651 & n27652;
  assign n27654 = n27653 ^ n2190;
  assign n27655 = n27654 ^ n27606;
  assign n27656 = ~n27610 & n27655;
  assign n27657 = n27656 ^ n27609;
  assign n27658 = n27657 ^ n27601;
  assign n27659 = ~n27605 & n27658;
  assign n27660 = n27659 ^ n27604;
  assign n27662 = n27661 ^ n27660;
  assign n27666 = n27665 ^ n27661;
  assign n27667 = ~n27662 & n27666;
  assign n27668 = n27667 ^ n27665;
  assign n27669 = n27668 ^ n27596;
  assign n27670 = n27600 & ~n27669;
  assign n27671 = n27670 ^ n27599;
  assign n27672 = n27671 ^ n27591;
  assign n27673 = n27595 & ~n27672;
  assign n27674 = n27673 ^ n27594;
  assign n27675 = n27674 ^ n27586;
  assign n27676 = n27590 & ~n27675;
  assign n27677 = n27676 ^ n27589;
  assign n27678 = n27677 ^ n27581;
  assign n27679 = ~n27585 & n27678;
  assign n27680 = n27679 ^ n27584;
  assign n27681 = n27680 ^ n27576;
  assign n27682 = n27580 & ~n27681;
  assign n27683 = n27682 ^ n27579;
  assign n27684 = n27683 ^ n27574;
  assign n27685 = n27575 & ~n27684;
  assign n27686 = n27685 ^ n793;
  assign n27687 = n27686 ^ n27572;
  assign n27688 = n27573 & ~n27687;
  assign n27689 = n27688 ^ n808;
  assign n27992 = n27689 ^ n887;
  assign n27993 = ~n27709 & ~n27992;
  assign n27994 = n27993 ^ n27708;
  assign n27995 = n27994 ^ n27987;
  assign n27996 = n27991 & n27995;
  assign n27997 = n27996 ^ n27990;
  assign n27998 = n27997 ^ n27985;
  assign n27999 = n27986 & ~n27998;
  assign n28000 = n27999 ^ n1043;
  assign n28001 = n28000 ^ n27980;
  assign n28002 = ~n27984 & n28001;
  assign n28003 = n28002 ^ n27983;
  assign n28004 = n28003 ^ n27975;
  assign n28005 = n27979 & ~n28004;
  assign n28006 = n28005 ^ n27978;
  assign n28008 = n28007 ^ n28006;
  assign n28009 = n2379 ^ n1396;
  assign n28010 = n28009 ^ n22347;
  assign n28011 = n28010 ^ n2276;
  assign n28012 = n28011 ^ n28007;
  assign n28013 = ~n28008 & n28012;
  assign n28014 = n28013 ^ n28011;
  assign n28015 = n28014 ^ n27973;
  assign n28016 = ~n27974 & ~n28015;
  assign n28017 = n28016 ^ n27970;
  assign n28018 = n28017 ^ n27968;
  assign n28019 = n27969 & n28018;
  assign n28020 = n28019 ^ n2516;
  assign n28021 = n28020 ^ n27966;
  assign n28022 = ~n27967 & n28021;
  assign n28023 = n28022 ^ n2531;
  assign n28044 = n28043 ^ n28023;
  assign n28049 = n28048 ^ n28044;
  assign n28051 = n26300 ^ n25818;
  assign n28052 = n27334 ^ n26300;
  assign n28053 = n28051 & n28052;
  assign n28054 = n28053 ^ n25818;
  assign n28050 = n28020 ^ n27967;
  assign n28055 = n28054 ^ n28050;
  assign n28058 = n26302 ^ n25957;
  assign n28059 = n27336 ^ n26302;
  assign n28060 = n28058 & ~n28059;
  assign n28061 = n28060 ^ n25957;
  assign n28056 = n28017 ^ n2516;
  assign n28057 = n28056 ^ n27968;
  assign n28062 = n28061 ^ n28057;
  assign n28069 = n26307 ^ n25822;
  assign n28070 = n27346 ^ n26307;
  assign n28071 = ~n28069 & ~n28070;
  assign n28072 = n28071 ^ n25822;
  assign n28063 = n28011 ^ n28008;
  assign n28064 = n26311 ^ n25220;
  assign n28065 = n27351 ^ n26311;
  assign n28066 = n28064 & ~n28065;
  assign n28067 = n28066 ^ n25220;
  assign n28068 = n28063 & n28067;
  assign n28073 = n28072 ^ n28068;
  assign n28074 = n28014 ^ n27974;
  assign n28075 = n28074 ^ n28068;
  assign n28076 = n28073 & n28075;
  assign n28077 = n28076 ^ n28072;
  assign n28078 = n28077 ^ n28057;
  assign n28079 = ~n28062 & n28078;
  assign n28080 = n28079 ^ n28061;
  assign n28081 = n28080 ^ n28050;
  assign n28082 = n28055 & n28081;
  assign n28083 = n28082 ^ n28054;
  assign n28084 = n28083 ^ n28044;
  assign n28085 = ~n28049 & ~n28084;
  assign n28086 = n28085 ^ n28048;
  assign n28088 = n28087 ^ n28086;
  assign n28089 = n26295 ^ n25810;
  assign n28090 = n27332 ^ n26295;
  assign n28091 = n28089 & ~n28090;
  assign n28092 = n28091 ^ n25810;
  assign n28093 = n28092 ^ n28086;
  assign n28094 = n28088 & ~n28093;
  assign n28095 = n28094 ^ n28087;
  assign n28096 = n28095 ^ n27833;
  assign n28097 = ~n27838 & ~n28096;
  assign n28098 = n28097 ^ n27837;
  assign n28099 = n28098 ^ n27192;
  assign n28100 = ~n27832 & n28099;
  assign n28101 = n28100 ^ n27831;
  assign n28103 = n28102 ^ n28101;
  assign n28104 = n26288 ^ n26064;
  assign n28105 = n27314 ^ n26288;
  assign n28106 = ~n28104 & ~n28105;
  assign n28107 = n28106 ^ n26064;
  assign n28108 = n28107 ^ n28101;
  assign n28109 = ~n28103 & ~n28108;
  assign n28110 = n28109 ^ n28102;
  assign n28111 = n28110 ^ n27286;
  assign n28112 = n27827 & ~n28111;
  assign n28113 = n28112 ^ n27826;
  assign n28114 = n28113 ^ n27820;
  assign n28115 = ~n27822 & n28114;
  assign n28116 = n28115 ^ n27821;
  assign n27814 = n27632 ^ n27619;
  assign n27815 = n27814 ^ n27620;
  assign n27810 = n26277 ^ n26258;
  assign n27811 = n27303 ^ n26277;
  assign n27812 = ~n27810 & ~n27811;
  assign n27813 = n27812 ^ n26258;
  assign n27816 = n27815 ^ n27813;
  assign n28217 = n28116 ^ n27816;
  assign n28218 = n28217 ^ n25244;
  assign n28219 = n28113 ^ n27822;
  assign n28220 = n28219 ^ n25248;
  assign n28221 = n28110 ^ n27827;
  assign n28222 = n28221 ^ n25252;
  assign n28223 = n28107 ^ n28102;
  assign n28224 = n28223 ^ n28101;
  assign n28225 = n28224 ^ n25256;
  assign n28226 = n28098 ^ n27831;
  assign n28227 = n28226 ^ n27192;
  assign n28228 = n28227 ^ n25262;
  assign n28251 = n28092 ^ n28087;
  assign n28252 = n28251 ^ n28086;
  assign n28229 = n28083 ^ n28049;
  assign n28230 = n28229 ^ n25273;
  assign n28231 = n28080 ^ n28055;
  assign n28232 = n28231 ^ n25277;
  assign n28233 = n28067 ^ n28063;
  assign n28234 = ~n25222 & n28233;
  assign n28235 = n28234 ^ n25283;
  assign n28236 = n28074 ^ n28073;
  assign n28237 = n28236 ^ n28234;
  assign n28238 = n28235 & n28237;
  assign n28239 = n28238 ^ n25283;
  assign n28240 = n28239 ^ n25278;
  assign n28241 = n28077 ^ n28062;
  assign n28242 = n28241 ^ n28239;
  assign n28243 = ~n28240 & n28242;
  assign n28244 = n28243 ^ n25278;
  assign n28245 = n28244 ^ n28231;
  assign n28246 = ~n28232 & n28245;
  assign n28247 = n28246 ^ n25277;
  assign n28248 = n28247 ^ n28229;
  assign n28249 = ~n28230 & n28248;
  assign n28250 = n28249 ^ n25273;
  assign n28253 = n28252 ^ n28250;
  assign n28254 = n28252 ^ n25269;
  assign n28255 = n28253 & n28254;
  assign n28256 = n28255 ^ n25269;
  assign n28257 = n28256 ^ n25265;
  assign n28258 = n28095 ^ n27837;
  assign n28259 = n28258 ^ n27833;
  assign n28260 = n28259 ^ n28256;
  assign n28261 = ~n28257 & n28260;
  assign n28262 = n28261 ^ n25265;
  assign n28263 = n28262 ^ n28227;
  assign n28264 = n28228 & n28263;
  assign n28265 = n28264 ^ n25262;
  assign n28266 = n28265 ^ n28224;
  assign n28267 = n28225 & ~n28266;
  assign n28268 = n28267 ^ n25256;
  assign n28269 = n28268 ^ n28221;
  assign n28270 = ~n28222 & ~n28269;
  assign n28271 = n28270 ^ n25252;
  assign n28272 = n28271 ^ n28219;
  assign n28273 = n28220 & ~n28272;
  assign n28274 = n28273 ^ n25248;
  assign n28275 = n28274 ^ n28217;
  assign n28276 = n28218 & ~n28275;
  assign n28277 = n28276 ^ n25244;
  assign n28117 = n28116 ^ n27813;
  assign n28118 = ~n27816 & ~n28117;
  assign n28119 = n28118 ^ n27815;
  assign n27808 = n27635 ^ n27616;
  assign n27804 = n26339 ^ n26272;
  assign n27805 = n27302 ^ n26272;
  assign n27806 = ~n27804 & n27805;
  assign n27807 = n27806 ^ n26339;
  assign n27809 = n27808 ^ n27807;
  assign n28215 = n28119 ^ n27809;
  assign n28216 = n28215 ^ n25241;
  assign n28350 = n28277 ^ n28216;
  assign n28351 = n28271 ^ n28220;
  assign n28352 = n28262 ^ n28228;
  assign n28353 = n28253 ^ n25269;
  assign n28354 = n28247 ^ n28230;
  assign n28355 = n28241 ^ n28240;
  assign n28356 = n28244 ^ n28232;
  assign n28357 = ~n28355 & ~n28356;
  assign n28358 = ~n28354 & n28357;
  assign n28359 = ~n28353 & ~n28358;
  assign n28360 = n28259 ^ n25265;
  assign n28361 = n28360 ^ n28256;
  assign n28362 = ~n28359 & ~n28361;
  assign n28363 = n28352 & n28362;
  assign n28364 = n28265 ^ n28225;
  assign n28365 = ~n28363 & n28364;
  assign n28366 = n28268 ^ n28222;
  assign n28367 = n28365 & ~n28366;
  assign n28368 = n28351 & ~n28367;
  assign n28369 = n28274 ^ n28218;
  assign n28370 = n28368 & n28369;
  assign n28371 = n28350 & n28370;
  assign n28120 = n28119 ^ n27807;
  assign n28121 = n27809 & n28120;
  assign n28122 = n28121 ^ n27808;
  assign n27802 = n27638 ^ n27614;
  assign n27798 = n26289 ^ n26271;
  assign n27799 = n27296 ^ n26271;
  assign n27800 = n27798 & n27799;
  assign n27801 = n27800 ^ n26289;
  assign n27803 = n27802 ^ n27801;
  assign n28281 = n28122 ^ n27803;
  assign n28348 = n28281 ^ n25237;
  assign n28278 = n28277 ^ n28215;
  assign n28279 = n28216 & ~n28278;
  assign n28280 = n28279 ^ n25241;
  assign n28349 = n28348 ^ n28280;
  assign n28489 = n28371 ^ n28349;
  assign n28493 = n28492 ^ n28489;
  assign n28494 = n28370 ^ n28350;
  assign n28498 = n28497 ^ n28494;
  assign n28571 = n28369 ^ n28368;
  assign n28566 = n28367 ^ n28351;
  assign n28499 = n28366 ^ n28365;
  assign n28500 = n28499 ^ n2124;
  assign n28502 = n26137 ^ n1948;
  assign n28503 = n28502 ^ n1760;
  assign n28504 = n28503 ^ n2118;
  assign n28501 = n28364 ^ n28363;
  assign n28505 = n28504 ^ n28501;
  assign n28552 = n28362 ^ n28352;
  assign n28506 = n28361 ^ n28359;
  assign n1644 = n1643 ^ n1629;
  assign n1654 = n1653 ^ n1644;
  assign n1658 = n1657 ^ n1654;
  assign n28507 = n28506 ^ n1658;
  assign n28511 = n28358 ^ n28353;
  assign n28512 = n28511 ^ n28510;
  assign n28516 = n28356 ^ n28355;
  assign n28513 = n26164 ^ n1478;
  assign n28514 = n28513 ^ n23119;
  assign n28515 = n28514 ^ n1574;
  assign n28517 = n28516 ^ n28515;
  assign n28521 = n28233 ^ n25222;
  assign n28522 = n28520 & ~n28521;
  assign n28526 = n28525 ^ n28522;
  assign n28527 = n28236 ^ n28235;
  assign n28528 = n28527 ^ n28525;
  assign n28529 = n28526 & n28528;
  assign n28530 = n28529 ^ n28522;
  assign n28531 = n28530 ^ n28355;
  assign n28535 = n28534 ^ n28530;
  assign n28536 = n28531 & n28535;
  assign n28537 = n28536 ^ n28534;
  assign n28538 = n28537 ^ n28516;
  assign n28539 = ~n28517 & n28538;
  assign n28540 = n28539 ^ n28515;
  assign n28541 = n28540 ^ n1584;
  assign n28542 = n28357 ^ n28354;
  assign n28543 = n28542 ^ n1584;
  assign n28544 = n28541 & ~n28543;
  assign n28545 = n28544 ^ n28540;
  assign n28546 = n28545 ^ n28511;
  assign n28547 = n28512 & ~n28546;
  assign n28548 = n28547 ^ n28510;
  assign n28549 = n28548 ^ n28506;
  assign n28550 = ~n28507 & n28549;
  assign n28551 = n28550 ^ n1658;
  assign n28553 = n28552 ^ n28551;
  assign n28557 = n28556 ^ n28552;
  assign n28558 = n28553 & ~n28557;
  assign n28559 = n28558 ^ n28556;
  assign n28560 = n28559 ^ n28504;
  assign n28561 = ~n28505 & ~n28560;
  assign n28562 = n28561 ^ n28501;
  assign n28563 = n28562 ^ n28499;
  assign n28564 = ~n28500 & ~n28563;
  assign n28565 = n28564 ^ n2124;
  assign n28567 = n28566 ^ n28565;
  assign n28568 = n28566 ^ n2139;
  assign n28569 = ~n28567 & n28568;
  assign n28570 = n28569 ^ n2139;
  assign n28572 = n28571 ^ n28570;
  assign n28573 = n28571 ^ n2157;
  assign n28574 = n28572 & ~n28573;
  assign n28575 = n28574 ^ n2157;
  assign n28576 = n28575 ^ n28494;
  assign n28577 = ~n28498 & n28576;
  assign n28578 = n28577 ^ n28497;
  assign n28579 = n28578 ^ n28489;
  assign n28580 = n28493 & ~n28579;
  assign n28581 = n28580 ^ n28492;
  assign n28869 = n28581 ^ n28487;
  assign n28372 = ~n28349 & n28371;
  assign n28282 = n28281 ^ n28280;
  assign n28283 = n28280 ^ n25237;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = n28284 ^ n25237;
  assign n28346 = n28285 ^ n25233;
  assign n28123 = n28122 ^ n27801;
  assign n28124 = ~n27803 & n28123;
  assign n28125 = n28124 ^ n27802;
  assign n27796 = n27643 ^ n27642;
  assign n27792 = n26284 ^ n26266;
  assign n27793 = n27290 ^ n26266;
  assign n27794 = ~n27792 & n27793;
  assign n27795 = n27794 ^ n26284;
  assign n27797 = n27796 ^ n27795;
  assign n28213 = n28125 ^ n27797;
  assign n28347 = n28346 ^ n28213;
  assign n28484 = n28372 ^ n28347;
  assign n28870 = n28869 ^ n28484;
  assign n27769 = n27665 ^ n27662;
  assign n30271 = n28870 ^ n27769;
  assign n29005 = n27302 ^ n26674;
  assign n27789 = n27646 ^ n2020;
  assign n27790 = n27789 ^ n27611;
  assign n29006 = n27790 ^ n27302;
  assign n29007 = ~n29005 & n29006;
  assign n29008 = n29007 ^ n26674;
  assign n28922 = n28545 ^ n28512;
  assign n29119 = n29008 ^ n28922;
  assign n28853 = n28542 ^ n28541;
  assign n28849 = n27303 ^ n26286;
  assign n28850 = n27796 ^ n27303;
  assign n28851 = ~n28849 & n28850;
  assign n28852 = n28851 ^ n26286;
  assign n28854 = n28853 ^ n28852;
  assign n28770 = n28537 ^ n28515;
  assign n28771 = n28770 ^ n28516;
  assign n28765 = n27399 ^ n26288;
  assign n28766 = n27802 ^ n27399;
  assign n28767 = n28765 & ~n28766;
  assign n28768 = n28767 ^ n26288;
  assign n28845 = n28771 ^ n28768;
  assign n28738 = n27314 ^ n26653;
  assign n28739 = n27815 ^ n27314;
  assign n28740 = n28738 & n28739;
  assign n28741 = n28740 ^ n26653;
  assign n28737 = n28527 ^ n28526;
  assign n28742 = n28741 ^ n28737;
  assign n28703 = n28521 ^ n28520;
  assign n28699 = n27317 ^ n26295;
  assign n28700 = n27821 ^ n27317;
  assign n28701 = ~n28699 & n28700;
  assign n28702 = n28701 ^ n26295;
  assign n28704 = n28703 ^ n28702;
  assign n27718 = n26603 ^ n25927;
  assign n27721 = n27720 ^ n26603;
  assign n27722 = ~n27718 & ~n27721;
  assign n27723 = n27722 ^ n25927;
  assign n27716 = n27686 ^ n808;
  assign n27717 = n27716 ^ n27572;
  assign n27724 = n27723 ^ n27717;
  assign n27731 = n27683 ^ n27575;
  assign n27725 = n26598 ^ n25792;
  assign n27728 = n27727 ^ n26598;
  assign n27729 = n27725 & ~n27728;
  assign n27730 = n27729 ^ n25792;
  assign n27732 = n27731 ^ n27730;
  assign n27739 = n27680 ^ n27580;
  assign n27733 = n27267 ^ n26582;
  assign n27736 = n27735 ^ n27267;
  assign n27737 = n27733 & ~n27736;
  assign n27738 = n27737 ^ n26582;
  assign n27740 = n27739 ^ n27738;
  assign n27746 = n27677 ^ n27584;
  assign n27747 = n27746 ^ n27581;
  assign n27741 = n27219 ^ n26559;
  assign n27743 = n27742 ^ n27219;
  assign n27744 = n27741 & ~n27743;
  assign n27745 = n27744 ^ n26559;
  assign n27748 = n27747 ^ n27745;
  assign n27751 = n27173 ^ n26473;
  assign n27753 = n27752 ^ n27173;
  assign n27754 = ~n27751 & ~n27753;
  assign n27755 = n27754 ^ n26473;
  assign n27749 = n27674 ^ n27589;
  assign n27750 = n27749 ^ n27586;
  assign n27756 = n27755 ^ n27750;
  assign n27762 = n27671 ^ n27595;
  assign n27757 = n27135 ^ n25804;
  assign n27759 = n27758 ^ n27135;
  assign n27760 = ~n27757 & ~n27759;
  assign n27761 = n27760 ^ n25804;
  assign n27763 = n27762 ^ n27761;
  assign n28150 = n27668 ^ n27600;
  assign n27764 = n26857 ^ n26267;
  assign n27766 = n27765 ^ n26857;
  assign n27767 = ~n27764 & n27766;
  assign n27768 = n27767 ^ n26267;
  assign n27770 = n27769 ^ n27768;
  assign n27776 = n27657 ^ n27605;
  assign n27771 = n26718 ^ n26327;
  assign n27773 = n27772 ^ n26718;
  assign n27774 = n27771 & n27773;
  assign n27775 = n27774 ^ n26327;
  assign n27777 = n27776 ^ n27775;
  assign n27782 = n27654 ^ n27609;
  assign n27783 = n27782 ^ n27606;
  assign n27778 = n26708 ^ n26274;
  assign n27779 = n27699 ^ n26708;
  assign n27780 = n27778 & ~n27779;
  assign n27781 = n27780 ^ n26274;
  assign n27784 = n27783 ^ n27781;
  assign n28132 = n27651 ^ n2190;
  assign n27785 = n26697 ^ n26334;
  assign n27786 = n27430 ^ n26697;
  assign n27787 = ~n27785 & n27786;
  assign n27788 = n27787 ^ n26334;
  assign n27791 = n27790 ^ n27788;
  assign n28126 = n28125 ^ n27796;
  assign n28127 = ~n27797 & ~n28126;
  assign n28128 = n28127 ^ n27795;
  assign n28129 = n28128 ^ n27790;
  assign n28130 = n27791 & ~n28129;
  assign n28131 = n28130 ^ n27788;
  assign n28133 = n28132 ^ n28131;
  assign n28134 = n26278 ^ n26264;
  assign n28135 = n27531 ^ n26264;
  assign n28136 = n28134 & ~n28135;
  assign n28137 = n28136 ^ n26278;
  assign n28138 = n28137 ^ n28132;
  assign n28139 = ~n28133 & n28138;
  assign n28140 = n28139 ^ n28137;
  assign n28141 = n28140 ^ n27783;
  assign n28142 = n27784 & ~n28141;
  assign n28143 = n28142 ^ n27781;
  assign n28144 = n28143 ^ n27775;
  assign n28145 = ~n27777 & n28144;
  assign n28146 = n28145 ^ n27776;
  assign n28147 = n28146 ^ n27769;
  assign n28148 = ~n27770 & n28147;
  assign n28149 = n28148 ^ n27768;
  assign n28151 = n28150 ^ n28149;
  assign n28152 = n27106 ^ n26380;
  assign n28153 = n27868 ^ n27106;
  assign n28154 = n28152 & ~n28153;
  assign n28155 = n28154 ^ n26380;
  assign n28156 = n28155 ^ n28150;
  assign n28157 = n28151 & ~n28156;
  assign n28158 = n28157 ^ n28155;
  assign n28159 = n28158 ^ n27762;
  assign n28160 = ~n27763 & n28159;
  assign n28161 = n28160 ^ n27761;
  assign n28162 = n28161 ^ n27750;
  assign n28163 = ~n27756 & n28162;
  assign n28164 = n28163 ^ n27755;
  assign n28165 = n28164 ^ n27747;
  assign n28166 = ~n27748 & ~n28165;
  assign n28167 = n28166 ^ n27745;
  assign n28168 = n28167 ^ n27739;
  assign n28169 = ~n27740 & n28168;
  assign n28170 = n28169 ^ n28167;
  assign n28171 = n28170 ^ n27731;
  assign n28172 = ~n27732 & ~n28171;
  assign n28173 = n28172 ^ n27730;
  assign n28174 = n28173 ^ n27717;
  assign n28175 = n27724 & n28174;
  assign n28176 = n28175 ^ n27723;
  assign n27711 = n26607 ^ n25934;
  assign n27712 = n27113 ^ n26607;
  assign n27713 = ~n27711 & ~n27712;
  assign n27714 = n27713 ^ n25934;
  assign n27710 = n27709 ^ n27689;
  assign n27715 = n27714 ^ n27710;
  assign n28188 = n28176 ^ n27715;
  assign n28189 = n28188 ^ n25213;
  assign n28190 = n28173 ^ n27723;
  assign n28191 = n28190 ^ n27717;
  assign n28192 = n28191 ^ n25166;
  assign n28319 = n28167 ^ n27740;
  assign n28193 = n28164 ^ n27745;
  assign n28194 = n28193 ^ n27747;
  assign n28195 = n28194 ^ n25802;
  assign n28196 = n28161 ^ n27755;
  assign n28197 = n28196 ^ n27750;
  assign n28198 = n28197 ^ n25856;
  assign n28199 = n28158 ^ n27761;
  assign n28200 = n28199 ^ n27762;
  assign n28201 = n28200 ^ n25840;
  assign n28202 = n28155 ^ n28151;
  assign n28203 = n28202 ^ n25782;
  assign n28204 = n28146 ^ n27768;
  assign n28205 = n28204 ^ n27769;
  assign n28206 = n28205 ^ n25555;
  assign n28207 = n28143 ^ n27777;
  assign n28208 = n28207 ^ n25543;
  assign n28209 = n28140 ^ n27784;
  assign n28210 = n28209 ^ n25529;
  assign n28211 = n28137 ^ n28133;
  assign n28212 = n28211 ^ n25413;
  assign n28289 = n28128 ^ n27788;
  assign n28290 = n28289 ^ n27790;
  assign n28214 = n28213 ^ n25233;
  assign n28286 = n28285 ^ n28213;
  assign n28287 = n28214 & n28286;
  assign n28288 = n28287 ^ n25233;
  assign n28291 = n28290 ^ n28288;
  assign n28292 = n28290 ^ n25227;
  assign n28293 = ~n28291 & n28292;
  assign n28294 = n28293 ^ n25227;
  assign n28295 = n28294 ^ n28211;
  assign n28296 = ~n28212 & ~n28295;
  assign n28297 = n28296 ^ n25413;
  assign n28298 = n28297 ^ n28209;
  assign n28299 = n28210 & n28298;
  assign n28300 = n28299 ^ n25529;
  assign n28301 = n28300 ^ n28207;
  assign n28302 = n28208 & n28301;
  assign n28303 = n28302 ^ n25543;
  assign n28304 = n28303 ^ n28205;
  assign n28305 = ~n28206 & ~n28304;
  assign n28306 = n28305 ^ n25555;
  assign n28307 = n28306 ^ n28202;
  assign n28308 = n28203 & n28307;
  assign n28309 = n28308 ^ n25782;
  assign n28310 = n28309 ^ n28200;
  assign n28311 = n28201 & ~n28310;
  assign n28312 = n28311 ^ n25840;
  assign n28313 = n28312 ^ n28197;
  assign n28314 = ~n28198 & ~n28313;
  assign n28315 = n28314 ^ n25856;
  assign n28316 = n28315 ^ n28194;
  assign n28317 = n28195 & n28316;
  assign n28318 = n28317 ^ n25802;
  assign n28320 = n28319 ^ n28318;
  assign n28321 = n28319 ^ n25907;
  assign n28322 = ~n28320 & n28321;
  assign n28323 = n28322 ^ n25907;
  assign n28324 = n28323 ^ n25139;
  assign n28325 = n28170 ^ n27732;
  assign n28326 = n28325 ^ n28323;
  assign n28327 = n28324 & n28326;
  assign n28328 = n28327 ^ n25139;
  assign n28329 = n28328 ^ n28191;
  assign n28330 = n28192 & n28329;
  assign n28331 = n28330 ^ n25166;
  assign n28332 = n28331 ^ n28188;
  assign n28333 = ~n28189 & n28332;
  assign n28334 = n28333 ^ n25213;
  assign n28181 = n26617 ^ n25918;
  assign n28182 = n27141 ^ n26617;
  assign n28183 = n28181 & n28182;
  assign n28184 = n28183 ^ n25918;
  assign n28180 = n27994 ^ n27991;
  assign n28185 = n28184 ^ n28180;
  assign n28177 = n28176 ^ n27710;
  assign n28178 = n27715 & n28177;
  assign n28179 = n28178 ^ n27714;
  assign n28186 = n28185 ^ n28179;
  assign n28187 = n28186 ^ n25345;
  assign n28335 = n28334 ^ n28187;
  assign n28336 = n28331 ^ n28189;
  assign n28337 = n28328 ^ n25166;
  assign n28338 = n28337 ^ n28191;
  assign n28339 = n28325 ^ n25139;
  assign n28340 = n28339 ^ n28323;
  assign n28341 = n28320 ^ n25907;
  assign n28342 = n28309 ^ n25840;
  assign n28343 = n28342 ^ n28200;
  assign n28344 = n28303 ^ n25555;
  assign n28345 = n28344 ^ n28205;
  assign n28373 = n28347 & ~n28372;
  assign n28374 = n28291 ^ n25227;
  assign n28375 = ~n28373 & n28374;
  assign n28376 = n28294 ^ n25413;
  assign n28377 = n28376 ^ n28211;
  assign n28378 = n28375 & ~n28377;
  assign n28379 = n28297 ^ n28210;
  assign n28380 = n28378 & ~n28379;
  assign n28381 = n28300 ^ n25543;
  assign n28382 = n28381 ^ n28207;
  assign n28383 = ~n28380 & ~n28382;
  assign n28384 = n28345 & ~n28383;
  assign n28385 = n28306 ^ n25782;
  assign n28386 = n28385 ^ n28202;
  assign n28387 = n28384 & n28386;
  assign n28388 = n28343 & ~n28387;
  assign n28389 = n28312 ^ n28198;
  assign n28390 = n28388 & ~n28389;
  assign n28391 = n28315 ^ n28195;
  assign n28392 = n28390 & ~n28391;
  assign n28393 = ~n28341 & ~n28392;
  assign n28394 = n28340 & n28393;
  assign n28395 = ~n28338 & n28394;
  assign n28396 = ~n28336 & n28395;
  assign n28397 = n28335 & ~n28396;
  assign n28408 = n28180 ^ n28179;
  assign n28409 = n28185 & ~n28408;
  assign n28410 = n28409 ^ n28184;
  assign n28403 = n26592 ^ n25914;
  assign n28404 = n27186 ^ n26592;
  assign n28405 = n28403 & ~n28404;
  assign n28406 = n28405 ^ n25914;
  assign n28402 = n27997 ^ n27986;
  assign n28407 = n28406 ^ n28402;
  assign n28411 = n28410 ^ n28407;
  assign n28398 = n28334 ^ n28186;
  assign n28399 = ~n28187 & ~n28398;
  assign n28400 = n28399 ^ n25345;
  assign n28401 = n28400 ^ n25337;
  assign n28412 = n28411 ^ n28401;
  assign n28413 = n28397 & ~n28412;
  assign n28425 = n28411 ^ n25337;
  assign n28426 = n28411 ^ n28400;
  assign n28427 = ~n28425 & ~n28426;
  assign n28428 = n28427 ^ n25337;
  assign n28418 = n25833 ^ n25798;
  assign n28419 = n27233 ^ n25798;
  assign n28420 = ~n28418 & n28419;
  assign n28421 = n28420 ^ n25833;
  assign n28415 = n28410 ^ n28402;
  assign n28416 = ~n28407 & n28415;
  assign n28417 = n28416 ^ n28406;
  assign n28422 = n28421 ^ n28417;
  assign n28414 = n28000 ^ n27984;
  assign n28423 = n28422 ^ n28414;
  assign n28424 = n28423 ^ n25224;
  assign n28429 = n28428 ^ n28424;
  assign n28659 = n28413 & n28429;
  assign n28654 = n28003 ^ n27979;
  assign n28650 = n28421 ^ n28414;
  assign n28651 = n28417 ^ n28414;
  assign n28652 = n28650 & ~n28651;
  assign n28653 = n28652 ^ n28421;
  assign n28655 = n28654 ^ n28653;
  assign n28646 = n26315 ^ n25829;
  assign n28647 = n27276 ^ n26315;
  assign n28648 = n28646 & ~n28647;
  assign n28649 = n28648 ^ n25829;
  assign n28656 = n28655 ^ n28649;
  assign n28642 = n28428 ^ n25224;
  assign n28643 = n28428 ^ n28423;
  assign n28644 = ~n28642 & ~n28643;
  assign n28645 = n28644 ^ n25224;
  assign n28657 = n28656 ^ n28645;
  assign n28658 = n28657 ^ n25355;
  assign n28660 = n28659 ^ n28658;
  assign n28638 = n26569 ^ n2608;
  assign n28639 = n28638 ^ n23223;
  assign n28640 = n28639 ^ n2561;
  assign n28431 = n26480 ^ n2584;
  assign n28432 = n28431 ^ n2429;
  assign n28433 = n28432 ^ n1544;
  assign n28430 = n28429 ^ n28413;
  assign n28434 = n28433 ^ n28430;
  assign n28436 = n26543 ^ n2595;
  assign n28437 = n28436 ^ n23044;
  assign n28438 = n28437 ^ n2420;
  assign n28435 = n28412 ^ n28397;
  assign n28439 = n28438 ^ n28435;
  assign n28440 = n28396 ^ n28335;
  assign n2319 = n2318 ^ n2282;
  assign n2320 = n2319 ^ n2315;
  assign n2324 = n2323 ^ n2320;
  assign n28441 = n28440 ^ n2324;
  assign n28621 = n28395 ^ n28336;
  assign n28442 = n28394 ^ n28338;
  assign n1318 = n1311 ^ n1224;
  assign n1325 = n1324 ^ n1318;
  assign n1329 = n1328 ^ n1325;
  assign n28443 = n28442 ^ n1329;
  assign n28444 = n28393 ^ n28340;
  assign n1148 = n1129 ^ n1056;
  assign n1149 = n1148 ^ n1145;
  assign n1153 = n1152 ^ n1149;
  assign n28445 = n28444 ^ n1153;
  assign n28446 = n28392 ^ n28341;
  assign n1133 = n1120 ^ n1061;
  assign n1134 = n1133 ^ n1020;
  assign n1138 = n1137 ^ n1134;
  assign n28447 = n28446 ^ n1138;
  assign n28448 = n28391 ^ n28390;
  assign n28449 = n28448 ^ n1010;
  assign n28450 = n28389 ^ n28388;
  assign n981 = n930 ^ n867;
  assign n991 = n990 ^ n981;
  assign n995 = n994 ^ n991;
  assign n28451 = n28450 ^ n995;
  assign n28452 = n28387 ^ n28343;
  assign n28456 = n28455 ^ n28452;
  assign n28457 = n28386 ^ n28384;
  assign n28461 = n28460 ^ n28457;
  assign n28465 = n28383 ^ n28345;
  assign n28466 = n28465 ^ n28464;
  assign n28468 = n26243 ^ n19314;
  assign n28469 = n28468 ^ n23067;
  assign n28470 = n28469 ^ n549;
  assign n28467 = n28382 ^ n28380;
  assign n28471 = n28470 ^ n28467;
  assign n28472 = n28379 ^ n28378;
  assign n28473 = n28472 ^ n644;
  assign n28475 = n26217 ^ n19321;
  assign n28476 = n28475 ^ n23074;
  assign n28477 = n28476 ^ n634;
  assign n28474 = n28377 ^ n28375;
  assign n28478 = n28477 ^ n28474;
  assign n28479 = n28374 ^ n28373;
  assign n28483 = n28482 ^ n28479;
  assign n28488 = n28487 ^ n28484;
  assign n28582 = n28581 ^ n28484;
  assign n28583 = ~n28488 & n28582;
  assign n28584 = n28583 ^ n28487;
  assign n28585 = n28584 ^ n28479;
  assign n28586 = n28483 & ~n28585;
  assign n28587 = n28586 ^ n28482;
  assign n28588 = n28587 ^ n28474;
  assign n28589 = n28478 & ~n28588;
  assign n28590 = n28589 ^ n28477;
  assign n28591 = n28590 ^ n28472;
  assign n28592 = n28473 & ~n28591;
  assign n28593 = n28592 ^ n644;
  assign n28594 = n28593 ^ n28467;
  assign n28595 = n28471 & ~n28594;
  assign n28596 = n28595 ^ n28470;
  assign n28597 = n28596 ^ n28465;
  assign n28598 = n28466 & ~n28597;
  assign n28599 = n28598 ^ n28464;
  assign n28600 = n28599 ^ n28457;
  assign n28601 = ~n28461 & n28600;
  assign n28602 = n28601 ^ n28460;
  assign n28603 = n28602 ^ n28452;
  assign n28604 = ~n28456 & n28603;
  assign n28605 = n28604 ^ n28455;
  assign n28606 = n28605 ^ n28450;
  assign n28607 = ~n28451 & n28606;
  assign n28608 = n28607 ^ n995;
  assign n28609 = n28608 ^ n28448;
  assign n28610 = ~n28449 & n28609;
  assign n28611 = n28610 ^ n1010;
  assign n28612 = n28611 ^ n28446;
  assign n28613 = ~n28447 & n28612;
  assign n28614 = n28613 ^ n1138;
  assign n28615 = n28614 ^ n28444;
  assign n28616 = ~n28445 & n28615;
  assign n28617 = n28616 ^ n1153;
  assign n28618 = n28617 ^ n28442;
  assign n28619 = n28443 & ~n28618;
  assign n28620 = n28619 ^ n1329;
  assign n28622 = n28621 ^ n28620;
  assign n28623 = n26487 ^ n19442;
  assign n28624 = n28623 ^ n1336;
  assign n28625 = n28624 ^ n2306;
  assign n28626 = n28625 ^ n28621;
  assign n28627 = ~n28622 & n28626;
  assign n28628 = n28627 ^ n28625;
  assign n28629 = n28628 ^ n28440;
  assign n28630 = ~n28441 & n28629;
  assign n28631 = n28630 ^ n2324;
  assign n28632 = n28631 ^ n28435;
  assign n28633 = ~n28439 & n28632;
  assign n28634 = n28633 ^ n28438;
  assign n28635 = n28634 ^ n28430;
  assign n28636 = n28434 & ~n28635;
  assign n28637 = n28636 ^ n28433;
  assign n28641 = n28640 ^ n28637;
  assign n28661 = n28660 ^ n28641;
  assign n27194 = n27193 ^ n26642;
  assign n27287 = n27286 ^ n27193;
  assign n27288 = n27194 & n27287;
  assign n27289 = n27288 ^ n26642;
  assign n28662 = n28661 ^ n27289;
  assign n28664 = n27332 ^ n26300;
  assign n28665 = n28102 ^ n27332;
  assign n28666 = ~n28664 & ~n28665;
  assign n28667 = n28666 ^ n26300;
  assign n28663 = n28634 ^ n28434;
  assign n28668 = n28667 ^ n28663;
  assign n28670 = n27375 ^ n26302;
  assign n28671 = n27375 ^ n27192;
  assign n28672 = ~n28670 & n28671;
  assign n28673 = n28672 ^ n26302;
  assign n28669 = n28631 ^ n28439;
  assign n28674 = n28673 ^ n28669;
  assign n28679 = n27336 ^ n26311;
  assign n28680 = n28087 ^ n27336;
  assign n28681 = n28679 & ~n28680;
  assign n28682 = n28681 ^ n26311;
  assign n28683 = n28625 ^ n28622;
  assign n28684 = n28682 & n28683;
  assign n28675 = n27334 ^ n26307;
  assign n28676 = n27833 ^ n27334;
  assign n28677 = ~n28675 & ~n28676;
  assign n28678 = n28677 ^ n26307;
  assign n28685 = n28684 ^ n28678;
  assign n28686 = n28628 ^ n28441;
  assign n28687 = n28686 ^ n28678;
  assign n28688 = ~n28685 & ~n28687;
  assign n28689 = n28688 ^ n28684;
  assign n28690 = n28689 ^ n28669;
  assign n28691 = ~n28674 & n28690;
  assign n28692 = n28691 ^ n28673;
  assign n28693 = n28692 ^ n28663;
  assign n28694 = ~n28668 & ~n28693;
  assign n28695 = n28694 ^ n28667;
  assign n28696 = n28695 ^ n28661;
  assign n28697 = n28662 & ~n28696;
  assign n28698 = n28697 ^ n27289;
  assign n28734 = n28703 ^ n28698;
  assign n28735 = ~n28704 & ~n28734;
  assign n28736 = n28735 ^ n28702;
  assign n28753 = n28737 ^ n28736;
  assign n28754 = ~n28742 & n28753;
  assign n28755 = n28754 ^ n28741;
  assign n28752 = n28534 ^ n28531;
  assign n28756 = n28755 ^ n28752;
  assign n28748 = n27304 ^ n26661;
  assign n28749 = n27808 ^ n27304;
  assign n28750 = n28748 & ~n28749;
  assign n28751 = n28750 ^ n26661;
  assign n28762 = n28752 ^ n28751;
  assign n28763 = n28756 & ~n28762;
  assign n28764 = n28763 ^ n28751;
  assign n28846 = n28771 ^ n28764;
  assign n28847 = ~n28845 & n28846;
  assign n28848 = n28847 ^ n28768;
  assign n29001 = n28852 ^ n28848;
  assign n29002 = n28854 & ~n29001;
  assign n29003 = n29002 ^ n28853;
  assign n29120 = n29119 ^ n29003;
  assign n29121 = n29120 ^ n26234;
  assign n28769 = n28768 ^ n28764;
  assign n28772 = n28771 ^ n28769;
  assign n28773 = n28772 ^ n26064;
  assign n28757 = n28756 ^ n28751;
  assign n28743 = n28742 ^ n28736;
  assign n28705 = n28704 ^ n28698;
  assign n28706 = n28705 ^ n25810;
  assign n28707 = n28695 ^ n27289;
  assign n28708 = n28707 ^ n28661;
  assign n28709 = n28708 ^ n25814;
  assign n28710 = n28692 ^ n28667;
  assign n28711 = n28710 ^ n28663;
  assign n28712 = n28711 ^ n25818;
  assign n28720 = n28689 ^ n28674;
  assign n28713 = n28683 ^ n28682;
  assign n28714 = n25220 & n28713;
  assign n28715 = n28714 ^ n25822;
  assign n28716 = n28686 ^ n28685;
  assign n28717 = n28716 ^ n28714;
  assign n28718 = n28715 & ~n28717;
  assign n28719 = n28718 ^ n25822;
  assign n28721 = n28720 ^ n28719;
  assign n28722 = n28720 ^ n25957;
  assign n28723 = n28721 & ~n28722;
  assign n28724 = n28723 ^ n25957;
  assign n28725 = n28724 ^ n28711;
  assign n28726 = n28712 & n28725;
  assign n28727 = n28726 ^ n25818;
  assign n28728 = n28727 ^ n28708;
  assign n28729 = ~n28709 & ~n28728;
  assign n28730 = n28729 ^ n25814;
  assign n28731 = n28730 ^ n28705;
  assign n28732 = n28706 & ~n28731;
  assign n28733 = n28732 ^ n25810;
  assign n28744 = n28743 ^ n28733;
  assign n28745 = n28743 ^ n25975;
  assign n28746 = n28744 & n28745;
  assign n28747 = n28746 ^ n25975;
  assign n28758 = n28757 ^ n28747;
  assign n28759 = n28757 ^ n26051;
  assign n28760 = ~n28758 & n28759;
  assign n28761 = n28760 ^ n26051;
  assign n28857 = n28772 ^ n28761;
  assign n28858 = n28773 & ~n28857;
  assign n28859 = n28858 ^ n26064;
  assign n29122 = n28859 ^ n26077;
  assign n28855 = n28854 ^ n28848;
  assign n29123 = n28859 ^ n28855;
  assign n29124 = ~n29122 & n29123;
  assign n29125 = n29124 ^ n26077;
  assign n29126 = n29125 ^ n29120;
  assign n29127 = n29121 & n29126;
  assign n29128 = n29127 ^ n26234;
  assign n29004 = n29003 ^ n28922;
  assign n29009 = n29008 ^ n29003;
  assign n29010 = n29004 & n29009;
  assign n29011 = n29010 ^ n28922;
  assign n28999 = n28548 ^ n28507;
  assign n28995 = n27296 ^ n26277;
  assign n28996 = n28132 ^ n27296;
  assign n28997 = ~n28995 & n28996;
  assign n28998 = n28997 ^ n26277;
  assign n29000 = n28999 ^ n28998;
  assign n29117 = n29011 ^ n29000;
  assign n29118 = n29117 ^ n26258;
  assign n29213 = n29128 ^ n29118;
  assign n28856 = n28855 ^ n26077;
  assign n28860 = n28859 ^ n28856;
  assign n28774 = n28773 ^ n28761;
  assign n28775 = n28721 ^ n25957;
  assign n28776 = n28724 ^ n28712;
  assign n28777 = n28775 & ~n28776;
  assign n28778 = n28727 ^ n28709;
  assign n28779 = n28777 & ~n28778;
  assign n28780 = n28730 ^ n28706;
  assign n28781 = ~n28779 & n28780;
  assign n28782 = n28744 ^ n25975;
  assign n28783 = ~n28781 & ~n28782;
  assign n28784 = n28758 ^ n26051;
  assign n28785 = n28783 & n28784;
  assign n28861 = ~n28774 & ~n28785;
  assign n29210 = ~n28860 & n28861;
  assign n29211 = n29125 ^ n29121;
  assign n29212 = ~n29210 & ~n29211;
  assign n29321 = n29213 ^ n29212;
  assign n29325 = n29324 ^ n29321;
  assign n29329 = n29211 ^ n29210;
  assign n28862 = n28861 ^ n28860;
  assign n28786 = n28785 ^ n28774;
  assign n1828 = n1820 ^ n1770;
  assign n1835 = n1834 ^ n1828;
  assign n1839 = n1838 ^ n1835;
  assign n28787 = n28786 ^ n1839;
  assign n28788 = n28784 ^ n28783;
  assign n28789 = n28788 ^ n1744;
  assign n28790 = n28782 ^ n28781;
  assign n28791 = n28790 ^ n1729;
  assign n28795 = n28780 ^ n28779;
  assign n28796 = n28795 ^ n28794;
  assign n28800 = n28776 ^ n28775;
  assign n28804 = n28803 ^ n28800;
  assign n28808 = n28807 ^ n28775;
  assign n28814 = n26967 ^ n19680;
  assign n28815 = n28814 ^ n1553;
  assign n28816 = n28815 ^ n18359;
  assign n28809 = n20097 ^ n2570;
  assign n28810 = n28809 ^ n2648;
  assign n28811 = n28810 ^ n1520;
  assign n28812 = n28713 ^ n25220;
  assign n28813 = n28811 & n28812;
  assign n28817 = n28816 ^ n28813;
  assign n28818 = n28716 ^ n28715;
  assign n28819 = n28818 ^ n28816;
  assign n28820 = n28817 & ~n28819;
  assign n28821 = n28820 ^ n28813;
  assign n28822 = n28821 ^ n28775;
  assign n28823 = n28808 & ~n28822;
  assign n28824 = n28823 ^ n28807;
  assign n28825 = n28824 ^ n28800;
  assign n28826 = n28804 & ~n28825;
  assign n28827 = n28826 ^ n28803;
  assign n28828 = n28827 ^ n28799;
  assign n28829 = n28778 ^ n28777;
  assign n28830 = n28829 ^ n28827;
  assign n28831 = n28828 & ~n28830;
  assign n28832 = n28831 ^ n28799;
  assign n28833 = n28832 ^ n28795;
  assign n28834 = ~n28796 & n28833;
  assign n28835 = n28834 ^ n28794;
  assign n28836 = n28835 ^ n28790;
  assign n28837 = ~n28791 & n28836;
  assign n28838 = n28837 ^ n1729;
  assign n28839 = n28838 ^ n28788;
  assign n28840 = ~n28789 & n28839;
  assign n28841 = n28840 ^ n1744;
  assign n28842 = n28841 ^ n1839;
  assign n28843 = n28787 & ~n28842;
  assign n28844 = n28843 ^ n28786;
  assign n28863 = n28862 ^ n28844;
  assign n29326 = n28866 ^ n28844;
  assign n29327 = n28863 & n29326;
  assign n29328 = n29327 ^ n28866;
  assign n29330 = n29329 ^ n29328;
  assign n29331 = n29329 ^ n1997;
  assign n29332 = n29330 & ~n29331;
  assign n29333 = n29332 ^ n1997;
  assign n29334 = n29333 ^ n29321;
  assign n29335 = ~n29325 & n29334;
  assign n29336 = n29335 ^ n29324;
  assign n29129 = n29128 ^ n29117;
  assign n29130 = n29118 & n29129;
  assign n29131 = n29130 ^ n26258;
  assign n29012 = n29011 ^ n28999;
  assign n29013 = n29000 & n29012;
  assign n29014 = n29013 ^ n28998;
  assign n28990 = n27290 ^ n26272;
  assign n28991 = n27783 ^ n27290;
  assign n28992 = n28990 & ~n28991;
  assign n28993 = n28992 ^ n26272;
  assign n29114 = n29014 ^ n28993;
  assign n28988 = n28556 ^ n28551;
  assign n28989 = n28988 ^ n28552;
  assign n29115 = n29114 ^ n28989;
  assign n29116 = n29115 ^ n26339;
  assign n29215 = n29131 ^ n29116;
  assign n29214 = n29212 & n29213;
  assign n29316 = n29215 ^ n29214;
  assign n29320 = n29319 ^ n29316;
  assign n29781 = n29336 ^ n29320;
  assign n30272 = n29781 ^ n28870;
  assign n30273 = ~n30271 & ~n30272;
  assign n30274 = n30273 ^ n27769;
  assign n28876 = n28578 ^ n28493;
  assign n29835 = n28876 ^ n27776;
  assign n29742 = n29333 ^ n29325;
  assign n29836 = n29742 ^ n28876;
  assign n29837 = ~n29835 & n29836;
  assign n29838 = n29837 ^ n27776;
  assign n29472 = n27815 ^ n27193;
  assign n29473 = n28853 ^ n27815;
  assign n29474 = n29472 & n29473;
  assign n29475 = n29474 ^ n27193;
  assign n29464 = n28617 ^ n1329;
  assign n29465 = n29464 ^ n28442;
  assign n29407 = n28614 ^ n1153;
  assign n29408 = n29407 ^ n28444;
  assign n29402 = n27351 ^ n25798;
  assign n29403 = n28050 ^ n27351;
  assign n29404 = n29402 & n29403;
  assign n29405 = n29404 ^ n25798;
  assign n29460 = n29408 ^ n29405;
  assign n29198 = n28608 ^ n28449;
  assign n29086 = n28605 ^ n28451;
  assign n29081 = n27186 ^ n26607;
  assign n29082 = n28063 ^ n27186;
  assign n29083 = ~n29081 & n29082;
  assign n29084 = n29083 ^ n26607;
  assign n29194 = n29086 ^ n29084;
  assign n28932 = n27141 ^ n26603;
  assign n28933 = n28654 ^ n27141;
  assign n28934 = ~n28932 & ~n28933;
  assign n28935 = n28934 ^ n26603;
  assign n28931 = n28602 ^ n28456;
  assign n28936 = n28935 ^ n28931;
  assign n28941 = n28599 ^ n28461;
  assign n28937 = n27113 ^ n26598;
  assign n28938 = n28414 ^ n27113;
  assign n28939 = ~n28937 & n28938;
  assign n28940 = n28939 ^ n26598;
  assign n28942 = n28941 ^ n28940;
  assign n28947 = n28596 ^ n28466;
  assign n28943 = n27720 ^ n27267;
  assign n28944 = n28402 ^ n27720;
  assign n28945 = ~n28943 & n28944;
  assign n28946 = n28945 ^ n27267;
  assign n28948 = n28947 ^ n28946;
  assign n29063 = n28593 ^ n28471;
  assign n28950 = n27735 ^ n27173;
  assign n28951 = n27735 ^ n27710;
  assign n28952 = n28950 & n28951;
  assign n28953 = n28952 ^ n27173;
  assign n28949 = n28590 ^ n28473;
  assign n28954 = n28953 ^ n28949;
  assign n28957 = n27742 ^ n27135;
  assign n28958 = n27742 ^ n27717;
  assign n28959 = n28957 & ~n28958;
  assign n28960 = n28959 ^ n27135;
  assign n28955 = n28587 ^ n28477;
  assign n28956 = n28955 ^ n28474;
  assign n28961 = n28960 ^ n28956;
  assign n28963 = n27868 ^ n26718;
  assign n28964 = n27868 ^ n27747;
  assign n28965 = ~n28963 & ~n28964;
  assign n28966 = n28965 ^ n26718;
  assign n28967 = n28966 ^ n28876;
  assign n29030 = n27765 ^ n26708;
  assign n29031 = n27765 ^ n27750;
  assign n29032 = n29030 & n29031;
  assign n29033 = n29032 ^ n26708;
  assign n28968 = n27772 ^ n26264;
  assign n28969 = n27772 ^ n27762;
  assign n28970 = n28968 & n28969;
  assign n28971 = n28970 ^ n26264;
  assign n28891 = n28572 ^ n2157;
  assign n28972 = n28971 ^ n28891;
  assign n28973 = n27699 ^ n26697;
  assign n28974 = n28150 ^ n27699;
  assign n28975 = ~n28973 & n28974;
  assign n28976 = n28975 ^ n26697;
  assign n28899 = n28567 ^ n2139;
  assign n28977 = n28976 ^ n28899;
  assign n28978 = n27531 ^ n26266;
  assign n28979 = n27769 ^ n27531;
  assign n28980 = ~n28978 & n28979;
  assign n28981 = n28980 ^ n26266;
  assign n28906 = n28562 ^ n28500;
  assign n28982 = n28981 ^ n28906;
  assign n28983 = n27430 ^ n26271;
  assign n28984 = n27776 ^ n27430;
  assign n28985 = n28983 & ~n28984;
  assign n28986 = n28985 ^ n26271;
  assign n28914 = n28559 ^ n28505;
  assign n28987 = n28986 ^ n28914;
  assign n28994 = n28993 ^ n28989;
  assign n29015 = n29014 ^ n28989;
  assign n29016 = n28994 & ~n29015;
  assign n29017 = n29016 ^ n28993;
  assign n29018 = n29017 ^ n28914;
  assign n29019 = n28987 & ~n29018;
  assign n29020 = n29019 ^ n28986;
  assign n29021 = n29020 ^ n28906;
  assign n29022 = n28982 & n29021;
  assign n29023 = n29022 ^ n28981;
  assign n29024 = n29023 ^ n28899;
  assign n29025 = n28977 & ~n29024;
  assign n29026 = n29025 ^ n28976;
  assign n29027 = n29026 ^ n28971;
  assign n29028 = n28972 & n29027;
  assign n29029 = n29028 ^ n28891;
  assign n29034 = n29033 ^ n29029;
  assign n28884 = n28575 ^ n28497;
  assign n28885 = n28884 ^ n28494;
  assign n29035 = n29029 ^ n28885;
  assign n29036 = ~n29034 & n29035;
  assign n29037 = n29036 ^ n28885;
  assign n29038 = n29037 ^ n28876;
  assign n29039 = n28967 & n29038;
  assign n29040 = n29039 ^ n28966;
  assign n29041 = n29040 ^ n28870;
  assign n29042 = n27758 ^ n26857;
  assign n29043 = n27758 ^ n27739;
  assign n29044 = n29042 & ~n29043;
  assign n29045 = n29044 ^ n26857;
  assign n29046 = n29045 ^ n29040;
  assign n29047 = ~n29041 & ~n29046;
  assign n29048 = n29047 ^ n28870;
  assign n28962 = n28584 ^ n28483;
  assign n29049 = n29048 ^ n28962;
  assign n29050 = n27752 ^ n27106;
  assign n29051 = n27752 ^ n27731;
  assign n29052 = ~n29050 & ~n29051;
  assign n29053 = n29052 ^ n27106;
  assign n29054 = n29053 ^ n28962;
  assign n29055 = n29049 & ~n29054;
  assign n29056 = n29055 ^ n29053;
  assign n29057 = n29056 ^ n28960;
  assign n29058 = n28961 & n29057;
  assign n29059 = n29058 ^ n28956;
  assign n29060 = n29059 ^ n28949;
  assign n29061 = n28954 & ~n29060;
  assign n29062 = n29061 ^ n28953;
  assign n29064 = n29063 ^ n29062;
  assign n29065 = n27727 ^ n27219;
  assign n29066 = n28180 ^ n27727;
  assign n29067 = ~n29065 & ~n29066;
  assign n29068 = n29067 ^ n27219;
  assign n29069 = n29068 ^ n29063;
  assign n29070 = ~n29064 & n29069;
  assign n29071 = n29070 ^ n29068;
  assign n29072 = n29071 ^ n28946;
  assign n29073 = n28948 & ~n29072;
  assign n29074 = n29073 ^ n28947;
  assign n29075 = n29074 ^ n28941;
  assign n29076 = n28942 & n29075;
  assign n29077 = n29076 ^ n28940;
  assign n29078 = n29077 ^ n28931;
  assign n29079 = n28936 & ~n29078;
  assign n29080 = n29079 ^ n28935;
  assign n29195 = n29086 ^ n29080;
  assign n29196 = ~n29194 & ~n29195;
  assign n29197 = n29196 ^ n29084;
  assign n29199 = n29198 ^ n29197;
  assign n29190 = n27233 ^ n26617;
  assign n29191 = n28074 ^ n27233;
  assign n29192 = n29190 & ~n29191;
  assign n29193 = n29192 ^ n26617;
  assign n29250 = n29198 ^ n29193;
  assign n29251 = n29199 & n29250;
  assign n29252 = n29251 ^ n29193;
  assign n29249 = n28611 ^ n28447;
  assign n29253 = n29252 ^ n29249;
  assign n29245 = n27276 ^ n26592;
  assign n29246 = n28057 ^ n27276;
  assign n29247 = n29245 & ~n29246;
  assign n29248 = n29247 ^ n26592;
  assign n29399 = n29249 ^ n29248;
  assign n29400 = ~n29253 & n29399;
  assign n29401 = n29400 ^ n29248;
  assign n29461 = n29408 ^ n29401;
  assign n29462 = ~n29460 & ~n29461;
  assign n29463 = n29462 ^ n29405;
  assign n29466 = n29465 ^ n29463;
  assign n29456 = n27346 ^ n26315;
  assign n29457 = n28044 ^ n27346;
  assign n29458 = n29456 & ~n29457;
  assign n29459 = n29458 ^ n26315;
  assign n29467 = n29466 ^ n29459;
  assign n29406 = n29405 ^ n29401;
  assign n29409 = n29408 ^ n29406;
  assign n29410 = n29409 ^ n25833;
  assign n29254 = n29253 ^ n29248;
  assign n29200 = n29199 ^ n29193;
  assign n29201 = n29200 ^ n25918;
  assign n29085 = n29084 ^ n29080;
  assign n29087 = n29086 ^ n29085;
  assign n29088 = n29087 ^ n25934;
  assign n29177 = n29074 ^ n28940;
  assign n29178 = n29177 ^ n28941;
  assign n29091 = n29071 ^ n28948;
  assign n29092 = n29091 ^ n26582;
  assign n29093 = n29068 ^ n29064;
  assign n29094 = n29093 ^ n26559;
  assign n29165 = n29059 ^ n28953;
  assign n29166 = n29165 ^ n28949;
  assign n29095 = n29056 ^ n28961;
  assign n29096 = n29095 ^ n25804;
  assign n29097 = n29053 ^ n29049;
  assign n29098 = n29097 ^ n26380;
  assign n29099 = n29045 ^ n28870;
  assign n29100 = n29099 ^ n29040;
  assign n29101 = n29100 ^ n26267;
  assign n29102 = n29037 ^ n28967;
  assign n29103 = n29102 ^ n26327;
  assign n29104 = n29033 ^ n28885;
  assign n29105 = n29104 ^ n29029;
  assign n29106 = n29105 ^ n26274;
  assign n29107 = n29026 ^ n28972;
  assign n29108 = n29107 ^ n26278;
  assign n29109 = n29023 ^ n28977;
  assign n29110 = n29109 ^ n26334;
  assign n29138 = n29020 ^ n28981;
  assign n29139 = n29138 ^ n28906;
  assign n29111 = n29017 ^ n28986;
  assign n29112 = n29111 ^ n28914;
  assign n29113 = n29112 ^ n26289;
  assign n29132 = n29131 ^ n29115;
  assign n29133 = ~n29116 & n29132;
  assign n29134 = n29133 ^ n26339;
  assign n29135 = n29134 ^ n29112;
  assign n29136 = n29113 & n29135;
  assign n29137 = n29136 ^ n26289;
  assign n29140 = n29139 ^ n29137;
  assign n29141 = n29139 ^ n26284;
  assign n29142 = ~n29140 & n29141;
  assign n29143 = n29142 ^ n26284;
  assign n29144 = n29143 ^ n29109;
  assign n29145 = ~n29110 & n29144;
  assign n29146 = n29145 ^ n26334;
  assign n29147 = n29146 ^ n29107;
  assign n29148 = ~n29108 & n29147;
  assign n29149 = n29148 ^ n26278;
  assign n29150 = n29149 ^ n29105;
  assign n29151 = n29106 & ~n29150;
  assign n29152 = n29151 ^ n26274;
  assign n29153 = n29152 ^ n29102;
  assign n29154 = ~n29103 & ~n29153;
  assign n29155 = n29154 ^ n26327;
  assign n29156 = n29155 ^ n29100;
  assign n29157 = n29101 & n29156;
  assign n29158 = n29157 ^ n26267;
  assign n29159 = n29158 ^ n29097;
  assign n29160 = ~n29098 & n29159;
  assign n29161 = n29160 ^ n26380;
  assign n29162 = n29161 ^ n29095;
  assign n29163 = n29096 & ~n29162;
  assign n29164 = n29163 ^ n25804;
  assign n29167 = n29166 ^ n29164;
  assign n29168 = n29166 ^ n26473;
  assign n29169 = n29167 & ~n29168;
  assign n29170 = n29169 ^ n26473;
  assign n29171 = n29170 ^ n29093;
  assign n29172 = n29094 & n29171;
  assign n29173 = n29172 ^ n26559;
  assign n29174 = n29173 ^ n29091;
  assign n29175 = n29092 & ~n29174;
  assign n29176 = n29175 ^ n26582;
  assign n29179 = n29178 ^ n29176;
  assign n29180 = n29178 ^ n25792;
  assign n29181 = ~n29179 & ~n29180;
  assign n29182 = n29181 ^ n25792;
  assign n29089 = n29077 ^ n28935;
  assign n29090 = n29089 ^ n28931;
  assign n29183 = n29182 ^ n29090;
  assign n29184 = n29090 ^ n25927;
  assign n29185 = ~n29183 & ~n29184;
  assign n29186 = n29185 ^ n25927;
  assign n29187 = n29186 ^ n29087;
  assign n29188 = ~n29088 & ~n29187;
  assign n29189 = n29188 ^ n25934;
  assign n29242 = n29200 ^ n29189;
  assign n29243 = ~n29201 & n29242;
  assign n29244 = n29243 ^ n25918;
  assign n29255 = n29254 ^ n29244;
  assign n29396 = n29254 ^ n25914;
  assign n29397 = ~n29255 & n29396;
  assign n29398 = n29397 ^ n25914;
  assign n29452 = n29409 ^ n29398;
  assign n29453 = ~n29410 & n29452;
  assign n29454 = n29453 ^ n25833;
  assign n29455 = n29454 ^ n25829;
  assign n29468 = n29467 ^ n29455;
  assign n29411 = n29410 ^ n29398;
  assign n29202 = n29201 ^ n29189;
  assign n29203 = n29186 ^ n25934;
  assign n29204 = n29203 ^ n29087;
  assign n29205 = n29183 ^ n25927;
  assign n29206 = n29179 ^ n25792;
  assign n29207 = n29158 ^ n29098;
  assign n29208 = n29149 ^ n29106;
  assign n29209 = n29140 ^ n26284;
  assign n29216 = n29214 & n29215;
  assign n29217 = n29134 ^ n29113;
  assign n29218 = n29216 & ~n29217;
  assign n29219 = ~n29209 & ~n29218;
  assign n29220 = n29143 ^ n29110;
  assign n29221 = ~n29219 & ~n29220;
  assign n29222 = n29146 ^ n29108;
  assign n29223 = n29221 & ~n29222;
  assign n29224 = n29208 & n29223;
  assign n29225 = n29152 ^ n29103;
  assign n29226 = ~n29224 & n29225;
  assign n29227 = n29155 ^ n29101;
  assign n29228 = ~n29226 & ~n29227;
  assign n29229 = ~n29207 & n29228;
  assign n29230 = n29161 ^ n29096;
  assign n29231 = ~n29229 & ~n29230;
  assign n29232 = n29167 ^ n26473;
  assign n29233 = n29231 & n29232;
  assign n29234 = n29170 ^ n29094;
  assign n29235 = n29233 & ~n29234;
  assign n29236 = n29173 ^ n29092;
  assign n29237 = ~n29235 & ~n29236;
  assign n29238 = n29206 & n29237;
  assign n29239 = ~n29205 & n29238;
  assign n29240 = n29204 & n29239;
  assign n29241 = n29202 & ~n29240;
  assign n29256 = n29255 ^ n25914;
  assign n29412 = n29241 & ~n29256;
  assign n29451 = n29411 & n29412;
  assign n29469 = n29468 ^ n29451;
  assign n29447 = n27232 ^ n1547;
  assign n29448 = n29447 ^ n2480;
  assign n29449 = n29448 ^ n2646;
  assign n29413 = n29412 ^ n29411;
  assign n29257 = n29256 ^ n29241;
  assign n29258 = n29257 ^ n2404;
  assign n29259 = n29240 ^ n29202;
  assign n2372 = n2348 ^ n2332;
  assign n2385 = n2384 ^ n2372;
  assign n2389 = n2388 ^ n2385;
  assign n29260 = n29259 ^ n2389;
  assign n29262 = n2289 ^ n1352;
  assign n29263 = n29262 ^ n23810;
  assign n29264 = n29263 ^ n2379;
  assign n29261 = n29239 ^ n29204;
  assign n29265 = n29264 ^ n29261;
  assign n29266 = n29238 ^ n29205;
  assign n1294 = n1251 ^ n1197;
  assign n1295 = n1294 ^ n1288;
  assign n1299 = n1298 ^ n1295;
  assign n29267 = n29266 ^ n1299;
  assign n29268 = n29237 ^ n29206;
  assign n1276 = n1236 ^ n1179;
  assign n1277 = n1276 ^ n1273;
  assign n1281 = n1280 ^ n1277;
  assign n29269 = n29268 ^ n1281;
  assign n29270 = n29236 ^ n29235;
  assign n29271 = n29270 ^ n1266;
  assign n29272 = n29234 ^ n29233;
  assign n29276 = n29275 ^ n29272;
  assign n29367 = n29232 ^ n29231;
  assign n29277 = n29230 ^ n29229;
  assign n29278 = n29277 ^ n773;
  assign n29280 = n27055 ^ n19974;
  assign n29281 = n29280 ^ n706;
  assign n29282 = n29281 ^ n763;
  assign n29279 = n29228 ^ n29207;
  assign n29283 = n29282 ^ n29279;
  assign n29284 = n29227 ^ n29226;
  assign n682 = n675 ^ n564;
  assign n695 = n694 ^ n682;
  assign n699 = n698 ^ n695;
  assign n29285 = n29284 ^ n699;
  assign n29287 = n26925 ^ n661;
  assign n29288 = n29287 ^ n23832;
  assign n29289 = n29288 ^ n689;
  assign n29286 = n29225 ^ n29224;
  assign n29290 = n29289 ^ n29286;
  assign n29292 = n26930 ^ n652;
  assign n29293 = n29292 ^ n23837;
  assign n29294 = n29293 ^ n18684;
  assign n29291 = n29223 ^ n29208;
  assign n29295 = n29294 ^ n29291;
  assign n29296 = n29222 ^ n29221;
  assign n29300 = n29299 ^ n29296;
  assign n29301 = n29220 ^ n29219;
  assign n29305 = n29304 ^ n29301;
  assign n29306 = n29218 ^ n29209;
  assign n29310 = n29309 ^ n29306;
  assign n29311 = n29217 ^ n29216;
  assign n29315 = n29314 ^ n29311;
  assign n29337 = n29336 ^ n29316;
  assign n29338 = ~n29320 & n29337;
  assign n29339 = n29338 ^ n29319;
  assign n29340 = n29339 ^ n29311;
  assign n29341 = n29315 & ~n29340;
  assign n29342 = n29341 ^ n29314;
  assign n29343 = n29342 ^ n29306;
  assign n29344 = n29310 & ~n29343;
  assign n29345 = n29344 ^ n29309;
  assign n29346 = n29345 ^ n29301;
  assign n29347 = ~n29305 & n29346;
  assign n29348 = n29347 ^ n29304;
  assign n29349 = n29348 ^ n29296;
  assign n29350 = n29300 & ~n29349;
  assign n29351 = n29350 ^ n29299;
  assign n29352 = n29351 ^ n29291;
  assign n29353 = ~n29295 & n29352;
  assign n29354 = n29353 ^ n29294;
  assign n29355 = n29354 ^ n29286;
  assign n29356 = ~n29290 & n29355;
  assign n29357 = n29356 ^ n29289;
  assign n29358 = n29357 ^ n699;
  assign n29359 = ~n29285 & ~n29358;
  assign n29360 = n29359 ^ n29284;
  assign n29361 = n29360 ^ n29282;
  assign n29362 = n29283 & n29361;
  assign n29363 = n29362 ^ n29279;
  assign n29364 = n29363 ^ n29277;
  assign n29365 = n29278 & ~n29364;
  assign n29366 = n29365 ^ n773;
  assign n29368 = n29367 ^ n29366;
  assign n29372 = n29371 ^ n29367;
  assign n29373 = ~n29368 & n29372;
  assign n29374 = n29373 ^ n29371;
  assign n29375 = n29374 ^ n29272;
  assign n29376 = ~n29276 & n29375;
  assign n29377 = n29376 ^ n29275;
  assign n29378 = n29377 ^ n29270;
  assign n29379 = ~n29271 & n29378;
  assign n29380 = n29379 ^ n1266;
  assign n29381 = n29380 ^ n29268;
  assign n29382 = ~n29269 & n29381;
  assign n29383 = n29382 ^ n1281;
  assign n29384 = n29383 ^ n29266;
  assign n29385 = n29267 & ~n29384;
  assign n29386 = n29385 ^ n1299;
  assign n29387 = n29386 ^ n29261;
  assign n29388 = ~n29265 & n29387;
  assign n29389 = n29388 ^ n29264;
  assign n29390 = n29389 ^ n29259;
  assign n29391 = ~n29260 & n29390;
  assign n29392 = n29391 ^ n2389;
  assign n29393 = n29392 ^ n29257;
  assign n29394 = ~n29258 & n29393;
  assign n29395 = n29394 ^ n2404;
  assign n29414 = n29413 ^ n29395;
  assign n2494 = n2486 ^ n2423;
  assign n2498 = n2497 ^ n2494;
  assign n2499 = n2498 ^ n2478;
  assign n29444 = n29413 ^ n2499;
  assign n29445 = ~n29414 & n29444;
  assign n29446 = n29445 ^ n2499;
  assign n29450 = n29449 ^ n29446;
  assign n29470 = n29469 ^ n29450;
  assign n29415 = n29414 ^ n2499;
  assign n28927 = n27821 ^ n27332;
  assign n28928 = n28771 ^ n27821;
  assign n28929 = n28927 & n28928;
  assign n28930 = n28929 ^ n27332;
  assign n29416 = n29415 ^ n28930;
  assign n29421 = n29392 ^ n29258;
  assign n29417 = n27375 ^ n27286;
  assign n29418 = n28752 ^ n27286;
  assign n29419 = ~n29417 & n29418;
  assign n29420 = n29419 ^ n27375;
  assign n29422 = n29421 ^ n29420;
  assign n29424 = n28102 ^ n27334;
  assign n29425 = n28737 ^ n28102;
  assign n29426 = n29424 & n29425;
  assign n29427 = n29426 ^ n27334;
  assign n29423 = n29389 ^ n29260;
  assign n29428 = n29427 ^ n29423;
  assign n29429 = n27336 ^ n27192;
  assign n29430 = n28703 ^ n27192;
  assign n29431 = n29429 & n29430;
  assign n29432 = n29431 ^ n27336;
  assign n29433 = n29386 ^ n29265;
  assign n29434 = n29432 & ~n29433;
  assign n29435 = n29434 ^ n29423;
  assign n29436 = n29428 & ~n29435;
  assign n29437 = n29436 ^ n29434;
  assign n29438 = n29437 ^ n29420;
  assign n29439 = n29422 & n29438;
  assign n29440 = n29439 ^ n29421;
  assign n29441 = n29440 ^ n29415;
  assign n29442 = n29416 & n29441;
  assign n29443 = n29442 ^ n28930;
  assign n29471 = n29470 ^ n29443;
  assign n29530 = n29475 ^ n29471;
  assign n29531 = n29530 ^ n26642;
  assign n29532 = n29440 ^ n29416;
  assign n29533 = n29532 ^ n26300;
  assign n29534 = n29437 ^ n29422;
  assign n29535 = n29534 ^ n26302;
  assign n29536 = n29433 ^ n29432;
  assign n29537 = n26311 & ~n29536;
  assign n29538 = n29537 ^ n26307;
  assign n29539 = n29434 ^ n29427;
  assign n29540 = n29539 ^ n29423;
  assign n29541 = n29540 ^ n29537;
  assign n29542 = ~n29538 & n29541;
  assign n29543 = n29542 ^ n26307;
  assign n29544 = n29543 ^ n29534;
  assign n29545 = n29535 & n29544;
  assign n29546 = n29545 ^ n26302;
  assign n29547 = n29546 ^ n29532;
  assign n29548 = n29533 & n29547;
  assign n29549 = n29548 ^ n26300;
  assign n29550 = n29549 ^ n29530;
  assign n29551 = n29531 & ~n29550;
  assign n29552 = n29551 ^ n26642;
  assign n29553 = n29552 ^ n26295;
  assign n29476 = n29475 ^ n29470;
  assign n29477 = ~n29471 & ~n29476;
  assign n29478 = n29477 ^ n29475;
  assign n28921 = n27808 ^ n27317;
  assign n28923 = n28922 ^ n27808;
  assign n28924 = ~n28921 & ~n28923;
  assign n28925 = n28924 ^ n27317;
  assign n28920 = n28812 ^ n28811;
  assign n28926 = n28925 ^ n28920;
  assign n29554 = n29478 ^ n28926;
  assign n29555 = n29554 ^ n29552;
  assign n29556 = ~n29553 & n29555;
  assign n29557 = n29556 ^ n26295;
  assign n29484 = n27802 ^ n27314;
  assign n29485 = n28999 ^ n27802;
  assign n29486 = n29484 & n29485;
  assign n29487 = n29486 ^ n27314;
  assign n29482 = n28818 ^ n28817;
  assign n29479 = n29478 ^ n28925;
  assign n29480 = ~n28926 & ~n29479;
  assign n29481 = n29480 ^ n28920;
  assign n29483 = n29482 ^ n29481;
  assign n29528 = n29487 ^ n29483;
  assign n29529 = n29528 ^ n26653;
  assign n29617 = n29557 ^ n29529;
  assign n29608 = n29549 ^ n29531;
  assign n29609 = n29543 ^ n26302;
  assign n29610 = n29609 ^ n29534;
  assign n29611 = n29546 ^ n26300;
  assign n29612 = n29611 ^ n29532;
  assign n29613 = n29610 & ~n29612;
  assign n29614 = n29608 & n29613;
  assign n29615 = n29554 ^ n29553;
  assign n29616 = ~n29614 & ~n29615;
  assign n29700 = n29617 ^ n29616;
  assign n29659 = n29615 ^ n29614;
  assign n29663 = n29662 ^ n29659;
  assign n29667 = n29612 ^ n29610;
  assign n1560 = n1559 ^ n1436;
  assign n1561 = n1560 ^ n1529;
  assign n1562 = n1561 ^ n1478;
  assign n29668 = n29667 ^ n1562;
  assign n29672 = n28042 ^ n2652;
  assign n29673 = n29672 ^ n2617;
  assign n29674 = n29673 ^ n19479;
  assign n29675 = n29536 ^ n26311;
  assign n29676 = n29674 & ~n29675;
  assign n29680 = n29679 ^ n29676;
  assign n29681 = n29540 ^ n29538;
  assign n29682 = n29681 ^ n29679;
  assign n29683 = n29680 & ~n29682;
  assign n29684 = n29683 ^ n29676;
  assign n29669 = n27119 ^ n20253;
  assign n29670 = n29669 ^ n24199;
  assign n29671 = n29670 ^ n1505;
  assign n29685 = n29684 ^ n29671;
  assign n29686 = n29684 ^ n29610;
  assign n29687 = n29685 & ~n29686;
  assign n29688 = n29687 ^ n29671;
  assign n29689 = n29688 ^ n29667;
  assign n29690 = n29668 & ~n29689;
  assign n29691 = n29690 ^ n1562;
  assign n29692 = n29691 ^ n29666;
  assign n29693 = n29613 ^ n29608;
  assign n29694 = n29693 ^ n29691;
  assign n29695 = n29692 & n29694;
  assign n29696 = n29695 ^ n29666;
  assign n29697 = n29696 ^ n29662;
  assign n29698 = n29663 & ~n29697;
  assign n29699 = n29698 ^ n29659;
  assign n29701 = n29700 ^ n29699;
  assign n29834 = n29704 ^ n29701;
  assign n29839 = n29838 ^ n29834;
  assign n29844 = n29696 ^ n29663;
  assign n29840 = n28885 ^ n27783;
  assign n29591 = n29330 ^ n1997;
  assign n29841 = n29591 ^ n28885;
  assign n29842 = n29840 & ~n29841;
  assign n29843 = n29842 ^ n27783;
  assign n29845 = n29844 ^ n29843;
  assign n29850 = n29693 ^ n29666;
  assign n29851 = n29850 ^ n29691;
  assign n29846 = n28891 ^ n28132;
  assign n28867 = n28866 ^ n28863;
  assign n29847 = n28891 ^ n28867;
  assign n29848 = n29846 & ~n29847;
  assign n29849 = n29848 ^ n28132;
  assign n29852 = n29851 ^ n29849;
  assign n29861 = n29685 ^ n29610;
  assign n29857 = n28906 ^ n27796;
  assign n28881 = n28838 ^ n1744;
  assign n28882 = n28881 ^ n28788;
  assign n29858 = n28906 ^ n28882;
  assign n29859 = n29857 & n29858;
  assign n29860 = n29859 ^ n27796;
  assign n29862 = n29861 ^ n29860;
  assign n30244 = n29681 ^ n29680;
  assign n30235 = n29675 ^ n29674;
  assign n30188 = n27833 ^ n27346;
  assign n30189 = n28661 ^ n27833;
  assign n30190 = ~n30188 & n30189;
  assign n30191 = n30190 ^ n27346;
  assign n30187 = n29383 ^ n29267;
  assign n30192 = n30191 ^ n30187;
  assign n29971 = n29377 ^ n1266;
  assign n29972 = n29971 ^ n29270;
  assign n29966 = n28044 ^ n27276;
  assign n29967 = n28669 ^ n28044;
  assign n29968 = n29966 & ~n29967;
  assign n29969 = n29968 ^ n27276;
  assign n30048 = n29972 ^ n29969;
  assign n29869 = n28050 ^ n27233;
  assign n29870 = n28686 ^ n28050;
  assign n29871 = n29869 & ~n29870;
  assign n29872 = n29871 ^ n27233;
  assign n29867 = n29374 ^ n29275;
  assign n29868 = n29867 ^ n29272;
  assign n29873 = n29872 ^ n29868;
  assign n29874 = n28057 ^ n27186;
  assign n29875 = n28683 ^ n28057;
  assign n29876 = n29874 & n29875;
  assign n29877 = n29876 ^ n27186;
  assign n29790 = n29371 ^ n29368;
  assign n29878 = n29877 ^ n29790;
  assign n29879 = n28074 ^ n27141;
  assign n29880 = n29465 ^ n28074;
  assign n29881 = ~n29879 & n29880;
  assign n29882 = n29881 ^ n27141;
  assign n29797 = n29363 ^ n29278;
  assign n29883 = n29882 ^ n29797;
  assign n29884 = n28063 ^ n27113;
  assign n29885 = n29408 ^ n28063;
  assign n29886 = n29884 & n29885;
  assign n29887 = n29886 ^ n27113;
  assign n29804 = n29360 ^ n29283;
  assign n29888 = n29887 ^ n29804;
  assign n29945 = n29357 ^ n29285;
  assign n29893 = n29354 ^ n29289;
  assign n29894 = n29893 ^ n29286;
  assign n29889 = n28414 ^ n27727;
  assign n29890 = n29198 ^ n28414;
  assign n29891 = n29889 & ~n29890;
  assign n29892 = n29891 ^ n27727;
  assign n29895 = n29894 ^ n29892;
  assign n29898 = n27758 ^ n27717;
  assign n29899 = n28947 ^ n27717;
  assign n29900 = n29898 & ~n29899;
  assign n29901 = n29900 ^ n27758;
  assign n29897 = n29342 ^ n29310;
  assign n29902 = n29901 ^ n29897;
  assign n29903 = n27868 ^ n27731;
  assign n29904 = n29063 ^ n27731;
  assign n29905 = ~n29903 & ~n29904;
  assign n29906 = n29905 ^ n27868;
  assign n29828 = n29339 ^ n29315;
  assign n29907 = n29906 ^ n29828;
  assign n29777 = n27765 ^ n27739;
  assign n29778 = n28949 ^ n27739;
  assign n29779 = ~n29777 & ~n29778;
  assign n29780 = n29779 ^ n27765;
  assign n29743 = n27772 ^ n27747;
  assign n29744 = n28956 ^ n27747;
  assign n29745 = n29743 & n29744;
  assign n29746 = n29745 ^ n27772;
  assign n29773 = n29746 ^ n29742;
  assign n29592 = n27750 ^ n27699;
  assign n29593 = n28962 ^ n27750;
  assign n29594 = ~n29592 & ~n29593;
  assign n29595 = n29594 ^ n27699;
  assign n29596 = n29595 ^ n29591;
  assign n28868 = n27762 ^ n27531;
  assign n28871 = n28870 ^ n27762;
  assign n28872 = ~n28868 & n28871;
  assign n28873 = n28872 ^ n27531;
  assign n29597 = n28873 ^ n28867;
  assign n28875 = n28150 ^ n27430;
  assign n28877 = n28876 ^ n28150;
  assign n28878 = ~n28875 & ~n28877;
  assign n28879 = n28878 ^ n27430;
  assign n28874 = n28841 ^ n28787;
  assign n28880 = n28879 ^ n28874;
  assign n28883 = n27769 ^ n27290;
  assign n28886 = n28885 ^ n27769;
  assign n28887 = ~n28883 & n28886;
  assign n28888 = n28887 ^ n27290;
  assign n28889 = n28888 ^ n28882;
  assign n28895 = n28835 ^ n28791;
  assign n28890 = n27776 ^ n27296;
  assign n28892 = n28891 ^ n27776;
  assign n28893 = ~n28890 & ~n28892;
  assign n28894 = n28893 ^ n27296;
  assign n28896 = n28895 ^ n28894;
  assign n28898 = n27783 ^ n27302;
  assign n28900 = n28899 ^ n27783;
  assign n28901 = ~n28898 & n28900;
  assign n28902 = n28901 ^ n27302;
  assign n28897 = n28832 ^ n28796;
  assign n28903 = n28902 ^ n28897;
  assign n28905 = n28132 ^ n27303;
  assign n28907 = n28906 ^ n28132;
  assign n28908 = n28905 & n28907;
  assign n28909 = n28908 ^ n27303;
  assign n28904 = n28829 ^ n28828;
  assign n28910 = n28909 ^ n28904;
  assign n28913 = n27790 ^ n27399;
  assign n28915 = n28914 ^ n27790;
  assign n28916 = ~n28913 & ~n28915;
  assign n28917 = n28916 ^ n27399;
  assign n28911 = n28824 ^ n28803;
  assign n28912 = n28911 ^ n28800;
  assign n28918 = n28917 ^ n28912;
  assign n29488 = n29487 ^ n29482;
  assign n29489 = ~n29483 & n29488;
  assign n29490 = n29489 ^ n29487;
  assign n28919 = n28821 ^ n28808;
  assign n29491 = n29490 ^ n28919;
  assign n29492 = n27796 ^ n27304;
  assign n29493 = n28989 ^ n27796;
  assign n29494 = n29492 & n29493;
  assign n29495 = n29494 ^ n27304;
  assign n29496 = n29495 ^ n28919;
  assign n29497 = ~n29491 & n29496;
  assign n29498 = n29497 ^ n29495;
  assign n29499 = n29498 ^ n28912;
  assign n29500 = n28918 & ~n29499;
  assign n29501 = n29500 ^ n28917;
  assign n29502 = n29501 ^ n28909;
  assign n29503 = ~n28910 & n29502;
  assign n29504 = n29503 ^ n28904;
  assign n29505 = n29504 ^ n28902;
  assign n29506 = ~n28903 & ~n29505;
  assign n29507 = n29506 ^ n28897;
  assign n29508 = n29507 ^ n28895;
  assign n29509 = ~n28896 & ~n29508;
  assign n29510 = n29509 ^ n28894;
  assign n29511 = n29510 ^ n28888;
  assign n29512 = n28889 & n29511;
  assign n29513 = n29512 ^ n28882;
  assign n29514 = n29513 ^ n28874;
  assign n29515 = ~n28880 & n29514;
  assign n29516 = n29515 ^ n28879;
  assign n29598 = n29516 ^ n28867;
  assign n29599 = n29597 & ~n29598;
  assign n29600 = n29599 ^ n28873;
  assign n29747 = n29600 ^ n29595;
  assign n29748 = n29596 & ~n29747;
  assign n29749 = n29748 ^ n29591;
  assign n29774 = n29749 ^ n29742;
  assign n29775 = n29773 & ~n29774;
  assign n29776 = n29775 ^ n29746;
  assign n29908 = n29780 ^ n29776;
  assign n29909 = n29781 ^ n29776;
  assign n29910 = n29908 & ~n29909;
  assign n29911 = n29910 ^ n29780;
  assign n29912 = n29911 ^ n29906;
  assign n29913 = ~n29907 & ~n29912;
  assign n29914 = n29913 ^ n29828;
  assign n29915 = n29914 ^ n29897;
  assign n29916 = n29902 & ~n29915;
  assign n29917 = n29916 ^ n29901;
  assign n29896 = n29345 ^ n29305;
  assign n29918 = n29917 ^ n29896;
  assign n29919 = n27752 ^ n27710;
  assign n29920 = n28941 ^ n27710;
  assign n29921 = ~n29919 & ~n29920;
  assign n29922 = n29921 ^ n27752;
  assign n29923 = n29922 ^ n29896;
  assign n29924 = n29918 & ~n29923;
  assign n29925 = n29924 ^ n29922;
  assign n29818 = n29348 ^ n29300;
  assign n29926 = n29925 ^ n29818;
  assign n29927 = n28180 ^ n27742;
  assign n29928 = n28931 ^ n28180;
  assign n29929 = ~n29927 & ~n29928;
  assign n29930 = n29929 ^ n27742;
  assign n29931 = n29930 ^ n29925;
  assign n29932 = n29926 & ~n29931;
  assign n29933 = n29932 ^ n29818;
  assign n29811 = n29351 ^ n29295;
  assign n29934 = n29933 ^ n29811;
  assign n29935 = n28402 ^ n27735;
  assign n29936 = n29086 ^ n28402;
  assign n29937 = n29935 & n29936;
  assign n29938 = n29937 ^ n27735;
  assign n29939 = n29938 ^ n29933;
  assign n29940 = ~n29934 & ~n29939;
  assign n29941 = n29940 ^ n29811;
  assign n29942 = n29941 ^ n29894;
  assign n29943 = n29895 & ~n29942;
  assign n29944 = n29943 ^ n29892;
  assign n29946 = n29945 ^ n29944;
  assign n29947 = n28654 ^ n27720;
  assign n29948 = n29249 ^ n28654;
  assign n29949 = ~n29947 & n29948;
  assign n29950 = n29949 ^ n27720;
  assign n29951 = n29950 ^ n29945;
  assign n29952 = ~n29946 & n29951;
  assign n29953 = n29952 ^ n29950;
  assign n29954 = n29953 ^ n29804;
  assign n29955 = ~n29888 & ~n29954;
  assign n29956 = n29955 ^ n29887;
  assign n29957 = n29956 ^ n29797;
  assign n29958 = n29883 & ~n29957;
  assign n29959 = n29958 ^ n29882;
  assign n29960 = n29959 ^ n29790;
  assign n29961 = ~n29878 & ~n29960;
  assign n29962 = n29961 ^ n29877;
  assign n29963 = n29962 ^ n29868;
  assign n29964 = n29873 & ~n29963;
  assign n29965 = n29964 ^ n29872;
  assign n30049 = n29972 ^ n29965;
  assign n30050 = n30048 & ~n30049;
  assign n30051 = n30050 ^ n29969;
  assign n30047 = n29380 ^ n29269;
  assign n30052 = n30051 ^ n30047;
  assign n30043 = n28087 ^ n27351;
  assign n30044 = n28663 ^ n28087;
  assign n30045 = n30043 & ~n30044;
  assign n30046 = n30045 ^ n27351;
  assign n30184 = n30047 ^ n30046;
  assign n30185 = ~n30052 & ~n30184;
  assign n30186 = n30185 ^ n30046;
  assign n30193 = n30192 ^ n30186;
  assign n30194 = n30193 ^ n26315;
  assign n30053 = n30052 ^ n30046;
  assign n30054 = n30053 ^ n25798;
  assign n29970 = n29969 ^ n29965;
  assign n29973 = n29972 ^ n29970;
  assign n29974 = n29973 ^ n26592;
  assign n29975 = n29962 ^ n29872;
  assign n29976 = n29975 ^ n29868;
  assign n29977 = n29976 ^ n26617;
  assign n29978 = n29959 ^ n29877;
  assign n29979 = n29978 ^ n29790;
  assign n29980 = n29979 ^ n26607;
  assign n29981 = n29956 ^ n29883;
  assign n29982 = n29981 ^ n26603;
  assign n29983 = n29953 ^ n29887;
  assign n29984 = n29983 ^ n29804;
  assign n29985 = n29984 ^ n26598;
  assign n29986 = n29950 ^ n29946;
  assign n29987 = n29986 ^ n27267;
  assign n30019 = n29941 ^ n29892;
  assign n30020 = n30019 ^ n29894;
  assign n29988 = n29938 ^ n29811;
  assign n29989 = n29988 ^ n29933;
  assign n29990 = n29989 ^ n27173;
  assign n29991 = n29930 ^ n29818;
  assign n29992 = n29991 ^ n29925;
  assign n29993 = n29992 ^ n27135;
  assign n29994 = n29922 ^ n29918;
  assign n29995 = n29994 ^ n27106;
  assign n29996 = n29914 ^ n29902;
  assign n29997 = n29996 ^ n26857;
  assign n29998 = n29911 ^ n29907;
  assign n29999 = n29998 ^ n26718;
  assign n29782 = n29781 ^ n29780;
  assign n29783 = n29782 ^ n29776;
  assign n29750 = n29749 ^ n29746;
  assign n29751 = n29750 ^ n29742;
  assign n29752 = n29751 ^ n26264;
  assign n29601 = n29600 ^ n29596;
  assign n29517 = n29516 ^ n28873;
  assign n29518 = n29517 ^ n28867;
  assign n29519 = n29518 ^ n26266;
  assign n29520 = n29513 ^ n28880;
  assign n29521 = n29520 ^ n26271;
  assign n29580 = n29510 ^ n28889;
  assign n29522 = n29507 ^ n28896;
  assign n29523 = n29522 ^ n26277;
  assign n29572 = n29504 ^ n28903;
  assign n29524 = n29498 ^ n28918;
  assign n29525 = n29524 ^ n26288;
  assign n29526 = n29495 ^ n29491;
  assign n29527 = n29526 ^ n26661;
  assign n29558 = n29557 ^ n29528;
  assign n29559 = n29529 & ~n29558;
  assign n29560 = n29559 ^ n26653;
  assign n29561 = n29560 ^ n29526;
  assign n29562 = n29527 & ~n29561;
  assign n29563 = n29562 ^ n26661;
  assign n29564 = n29563 ^ n29524;
  assign n29565 = n29525 & ~n29564;
  assign n29566 = n29565 ^ n26288;
  assign n29567 = n29566 ^ n26286;
  assign n29568 = n29501 ^ n28910;
  assign n29569 = n29568 ^ n29566;
  assign n29570 = n29567 & n29569;
  assign n29571 = n29570 ^ n26286;
  assign n29573 = n29572 ^ n29571;
  assign n29574 = n29572 ^ n26674;
  assign n29575 = n29573 & n29574;
  assign n29576 = n29575 ^ n26674;
  assign n29577 = n29576 ^ n29522;
  assign n29578 = ~n29523 & n29577;
  assign n29579 = n29578 ^ n26277;
  assign n29581 = n29580 ^ n29579;
  assign n29582 = n29580 ^ n26272;
  assign n29583 = n29581 & ~n29582;
  assign n29584 = n29583 ^ n26272;
  assign n29585 = n29584 ^ n29520;
  assign n29586 = ~n29521 & n29585;
  assign n29587 = n29586 ^ n26271;
  assign n29588 = n29587 ^ n29518;
  assign n29589 = ~n29519 & ~n29588;
  assign n29590 = n29589 ^ n26266;
  assign n29602 = n29601 ^ n29590;
  assign n29753 = n29601 ^ n26697;
  assign n29754 = n29602 & ~n29753;
  assign n29755 = n29754 ^ n26697;
  assign n29770 = n29755 ^ n29751;
  assign n29771 = n29752 & n29770;
  assign n29772 = n29771 ^ n26264;
  assign n30000 = n29783 ^ n29772;
  assign n30001 = n29772 ^ n26708;
  assign n30002 = ~n30000 & n30001;
  assign n30003 = n30002 ^ n26708;
  assign n30004 = n30003 ^ n29998;
  assign n30005 = n29999 & n30004;
  assign n30006 = n30005 ^ n26718;
  assign n30007 = n30006 ^ n29996;
  assign n30008 = n29997 & ~n30007;
  assign n30009 = n30008 ^ n26857;
  assign n30010 = n30009 ^ n29994;
  assign n30011 = n29995 & n30010;
  assign n30012 = n30011 ^ n27106;
  assign n30013 = n30012 ^ n29992;
  assign n30014 = n29993 & n30013;
  assign n30015 = n30014 ^ n27135;
  assign n30016 = n30015 ^ n29989;
  assign n30017 = ~n29990 & n30016;
  assign n30018 = n30017 ^ n27173;
  assign n30021 = n30020 ^ n30018;
  assign n30022 = n30020 ^ n27219;
  assign n30023 = n30021 & ~n30022;
  assign n30024 = n30023 ^ n27219;
  assign n30025 = n30024 ^ n29986;
  assign n30026 = ~n29987 & n30025;
  assign n30027 = n30026 ^ n27267;
  assign n30028 = n30027 ^ n29984;
  assign n30029 = ~n29985 & ~n30028;
  assign n30030 = n30029 ^ n26598;
  assign n30031 = n30030 ^ n29981;
  assign n30032 = ~n29982 & n30031;
  assign n30033 = n30032 ^ n26603;
  assign n30034 = n30033 ^ n29979;
  assign n30035 = ~n29980 & ~n30034;
  assign n30036 = n30035 ^ n26607;
  assign n30037 = n30036 ^ n29976;
  assign n30038 = n29977 & n30037;
  assign n30039 = n30038 ^ n26617;
  assign n30040 = n30039 ^ n29973;
  assign n30041 = n29974 & ~n30040;
  assign n30042 = n30041 ^ n26592;
  assign n30181 = n30053 ^ n30042;
  assign n30182 = n30054 & n30181;
  assign n30183 = n30182 ^ n25798;
  assign n30195 = n30194 ^ n30183;
  assign n30055 = n30054 ^ n30042;
  assign n30056 = n30039 ^ n26592;
  assign n30057 = n30056 ^ n29973;
  assign n30058 = n30036 ^ n29977;
  assign n30059 = n30015 ^ n27173;
  assign n30060 = n30059 ^ n29989;
  assign n30061 = n30009 ^ n29995;
  assign n29784 = n29783 ^ n26708;
  assign n29785 = n29784 ^ n29772;
  assign n29756 = n29755 ^ n29752;
  assign n29603 = n29602 ^ n26697;
  assign n29604 = n29568 ^ n26286;
  assign n29605 = n29604 ^ n29566;
  assign n29606 = n29563 ^ n26288;
  assign n29607 = n29606 ^ n29524;
  assign n29618 = ~n29616 & ~n29617;
  assign n29619 = n29560 ^ n29527;
  assign n29620 = n29618 & ~n29619;
  assign n29621 = n29607 & ~n29620;
  assign n29622 = ~n29605 & n29621;
  assign n29623 = n29573 ^ n26674;
  assign n29624 = ~n29622 & ~n29623;
  assign n29625 = n29576 ^ n29523;
  assign n29626 = n29624 & ~n29625;
  assign n29627 = n29581 ^ n26272;
  assign n29628 = n29626 & ~n29627;
  assign n29629 = n29584 ^ n29521;
  assign n29630 = n29628 & ~n29629;
  assign n29631 = n29587 ^ n29519;
  assign n29632 = ~n29630 & n29631;
  assign n29757 = n29603 & ~n29632;
  assign n29786 = ~n29756 & n29757;
  assign n30062 = n29785 & n29786;
  assign n30063 = n30003 ^ n29999;
  assign n30064 = ~n30062 & ~n30063;
  assign n30065 = n30006 ^ n26857;
  assign n30066 = n30065 ^ n29996;
  assign n30067 = ~n30064 & ~n30066;
  assign n30068 = ~n30061 & n30067;
  assign n30069 = n30012 ^ n29993;
  assign n30070 = ~n30068 & ~n30069;
  assign n30071 = ~n30060 & n30070;
  assign n30072 = n30021 ^ n27219;
  assign n30073 = n30071 & ~n30072;
  assign n30074 = n30024 ^ n27267;
  assign n30075 = n30074 ^ n29986;
  assign n30076 = ~n30073 & n30075;
  assign n30077 = n30027 ^ n29985;
  assign n30078 = n30076 & n30077;
  assign n30079 = n30030 ^ n29982;
  assign n30080 = n30078 & ~n30079;
  assign n30081 = n30033 ^ n26607;
  assign n30082 = n30081 ^ n29979;
  assign n30083 = n30080 & ~n30082;
  assign n30084 = n30058 & ~n30083;
  assign n30085 = ~n30057 & n30084;
  assign n30180 = ~n30055 & n30085;
  assign n30196 = n30195 ^ n30180;
  assign n30086 = n30085 ^ n30055;
  assign n2592 = n2516 ^ n2466;
  assign n2599 = n2598 ^ n2592;
  assign n2600 = n2599 ^ n2584;
  assign n30087 = n30086 ^ n2600;
  assign n30089 = n27973 ^ n2440;
  assign n30090 = n30089 ^ n24538;
  assign n30091 = n30090 ^ n2595;
  assign n30088 = n30084 ^ n30057;
  assign n30092 = n30091 ^ n30088;
  assign n30094 = n28011 ^ n2455;
  assign n30095 = n30094 ^ n24543;
  assign n30096 = n30095 ^ n2318;
  assign n30093 = n30083 ^ n30058;
  assign n30097 = n30096 ^ n30093;
  assign n30099 = n27978 ^ n1406;
  assign n30100 = n30099 ^ n1316;
  assign n30101 = n30100 ^ n19442;
  assign n30098 = n30082 ^ n30080;
  assign n30102 = n30101 ^ n30098;
  assign n30159 = n30079 ^ n30078;
  assign n30103 = n30077 ^ n30076;
  assign n30104 = n30103 ^ n1130;
  assign n30105 = n30075 ^ n30073;
  assign n30109 = n30108 ^ n30105;
  assign n30110 = n30072 ^ n30071;
  assign n30111 = n30110 ^ n969;
  assign n30112 = n30070 ^ n30060;
  assign n863 = n832 ^ n808;
  assign n864 = n863 ^ n860;
  assign n868 = n867 ^ n864;
  assign n30113 = n30112 ^ n868;
  assign n30114 = n30069 ^ n30068;
  assign n836 = n823 ^ n793;
  assign n849 = n848 ^ n836;
  assign n853 = n852 ^ n849;
  assign n30115 = n30114 ^ n853;
  assign n30116 = n30067 ^ n30061;
  assign n30120 = n30119 ^ n30116;
  assign n30133 = n30066 ^ n30064;
  assign n30121 = n30063 ^ n30062;
  assign n30125 = n30124 ^ n30121;
  assign n29787 = n29786 ^ n29785;
  assign n29758 = n29757 ^ n29756;
  assign n29633 = n29632 ^ n29603;
  assign n29637 = n29636 ^ n29633;
  assign n29731 = n29631 ^ n29630;
  assign n29638 = n29629 ^ n29628;
  assign n29642 = n29641 ^ n29638;
  assign n29643 = n29627 ^ n29626;
  assign n29647 = n29646 ^ n29643;
  assign n29648 = n29625 ^ n29624;
  assign n29649 = n29648 ^ n2110;
  assign n29650 = n29623 ^ n29622;
  assign n29651 = n29650 ^ n2095;
  assign n29714 = n29621 ^ n29605;
  assign n29652 = n29620 ^ n29607;
  assign n1935 = n1865 ^ n1809;
  assign n1945 = n1944 ^ n1935;
  assign n1949 = n1948 ^ n1945;
  assign n29653 = n29652 ^ n1949;
  assign n29657 = n29619 ^ n29618;
  assign n29654 = n27619 ^ n1794;
  assign n29655 = n29654 ^ n24182;
  assign n29656 = n29655 ^ n1942;
  assign n29658 = n29657 ^ n29656;
  assign n29705 = n29704 ^ n29700;
  assign n29706 = n29701 & ~n29705;
  assign n29707 = n29706 ^ n29704;
  assign n29708 = n29707 ^ n29657;
  assign n29709 = n29658 & ~n29708;
  assign n29710 = n29709 ^ n29656;
  assign n29711 = n29710 ^ n29652;
  assign n29712 = ~n29653 & n29711;
  assign n29713 = n29712 ^ n1949;
  assign n29715 = n29714 ^ n29713;
  assign n29716 = n29714 ^ n1964;
  assign n29717 = n29715 & ~n29716;
  assign n29718 = n29717 ^ n1964;
  assign n29719 = n29718 ^ n29650;
  assign n29720 = ~n29651 & n29719;
  assign n29721 = n29720 ^ n2095;
  assign n29722 = n29721 ^ n29648;
  assign n29723 = n29649 & ~n29722;
  assign n29724 = n29723 ^ n2110;
  assign n29725 = n29724 ^ n29643;
  assign n29726 = n29647 & ~n29725;
  assign n29727 = n29726 ^ n29646;
  assign n29728 = n29727 ^ n29638;
  assign n29729 = n29642 & ~n29728;
  assign n29730 = n29729 ^ n29641;
  assign n29732 = n29731 ^ n29730;
  assign n29736 = n29735 ^ n29730;
  assign n29737 = n29732 & n29736;
  assign n29738 = n29737 ^ n29735;
  assign n29739 = n29738 ^ n29633;
  assign n29740 = n29637 & ~n29739;
  assign n29741 = n29740 ^ n29636;
  assign n29759 = n29758 ^ n29741;
  assign n29760 = n27599 ^ n20610;
  assign n29761 = n29760 ^ n614;
  assign n29762 = n29761 ^ n19321;
  assign n29763 = n29762 ^ n29758;
  assign n29764 = ~n29759 & n29763;
  assign n29765 = n29764 ^ n29762;
  assign n30126 = n29787 ^ n29765;
  assign n29766 = n27594 ^ n20605;
  assign n29767 = n29766 ^ n24266;
  assign n29768 = n29767 ^ n530;
  assign n30127 = n29787 ^ n29768;
  assign n30128 = n30126 & ~n30127;
  assign n30129 = n30128 ^ n29768;
  assign n30130 = n30129 ^ n30121;
  assign n30131 = n30125 & ~n30130;
  assign n30132 = n30131 ^ n30124;
  assign n30134 = n30133 ^ n30132;
  assign n30135 = n27584 ^ n747;
  assign n30136 = n30135 ^ n24290;
  assign n30137 = n30136 ^ n19407;
  assign n30138 = n30137 ^ n30133;
  assign n30139 = n30134 & ~n30138;
  assign n30140 = n30139 ^ n30137;
  assign n30141 = n30140 ^ n30116;
  assign n30142 = n30120 & ~n30141;
  assign n30143 = n30142 ^ n30119;
  assign n30144 = n30143 ^ n853;
  assign n30145 = n30115 & ~n30144;
  assign n30146 = n30145 ^ n30114;
  assign n30147 = n30146 ^ n30112;
  assign n30148 = ~n30113 & n30147;
  assign n30149 = n30148 ^ n868;
  assign n30150 = n30149 ^ n30110;
  assign n30151 = ~n30111 & n30150;
  assign n30152 = n30151 ^ n969;
  assign n30153 = n30152 ^ n30105;
  assign n30154 = n30109 & ~n30153;
  assign n30155 = n30154 ^ n30108;
  assign n30156 = n30155 ^ n30103;
  assign n30157 = ~n30104 & n30156;
  assign n30158 = n30157 ^ n1130;
  assign n30160 = n30159 ^ n30158;
  assign n30161 = n27983 ^ n1388;
  assign n30162 = n30161 ^ n24550;
  assign n30163 = n30162 ^ n1311;
  assign n30164 = n30163 ^ n30159;
  assign n30165 = ~n30160 & n30164;
  assign n30166 = n30165 ^ n30163;
  assign n30167 = n30166 ^ n30098;
  assign n30168 = n30102 & ~n30167;
  assign n30169 = n30168 ^ n30101;
  assign n30170 = n30169 ^ n30093;
  assign n30171 = ~n30097 & n30170;
  assign n30172 = n30171 ^ n30096;
  assign n30173 = n30172 ^ n30088;
  assign n30174 = ~n30092 & n30173;
  assign n30175 = n30174 ^ n30091;
  assign n30176 = n30175 ^ n30086;
  assign n30177 = ~n30087 & n30176;
  assign n30178 = n30177 ^ n2600;
  assign n30179 = n30178 ^ n2609;
  assign n30197 = n30196 ^ n30179;
  assign n29863 = n28999 ^ n27815;
  assign n29864 = n28999 ^ n28904;
  assign n29865 = n29863 & n29864;
  assign n29866 = n29865 ^ n27815;
  assign n30198 = n30197 ^ n29866;
  assign n30215 = n28853 ^ n27286;
  assign n30216 = n28919 ^ n28853;
  assign n30217 = n30215 & ~n30216;
  assign n30218 = n30217 ^ n27286;
  assign n30206 = n28771 ^ n28102;
  assign n30207 = n29482 ^ n28771;
  assign n30208 = ~n30206 & n30207;
  assign n30209 = n30208 ^ n28102;
  assign n30200 = n30166 ^ n30102;
  assign n30201 = n28752 ^ n27192;
  assign n30202 = n28920 ^ n28752;
  assign n30203 = ~n30201 & n30202;
  assign n30204 = n30203 ^ n27192;
  assign n30205 = n30200 & n30204;
  assign n30210 = n30209 ^ n30205;
  assign n30211 = n30169 ^ n30097;
  assign n30212 = n30211 ^ n30205;
  assign n30213 = n30210 & n30212;
  assign n30214 = n30213 ^ n30209;
  assign n30219 = n30218 ^ n30214;
  assign n30220 = n30172 ^ n30092;
  assign n30221 = n30220 ^ n30214;
  assign n30222 = n30219 & n30221;
  assign n30223 = n30222 ^ n30218;
  assign n30199 = n30175 ^ n30087;
  assign n30224 = n30223 ^ n30199;
  assign n30225 = n28922 ^ n27821;
  assign n30226 = n28922 ^ n28912;
  assign n30227 = n30225 & ~n30226;
  assign n30228 = n30227 ^ n27821;
  assign n30229 = n30228 ^ n30223;
  assign n30230 = ~n30224 & ~n30229;
  assign n30231 = n30230 ^ n30199;
  assign n30232 = n30231 ^ n30197;
  assign n30233 = n30198 & ~n30232;
  assign n30234 = n30233 ^ n29866;
  assign n30236 = n30235 ^ n30234;
  assign n30237 = n28989 ^ n27808;
  assign n30238 = n28989 ^ n28897;
  assign n30239 = ~n30237 & ~n30238;
  assign n30240 = n30239 ^ n27808;
  assign n30241 = n30240 ^ n30235;
  assign n30242 = ~n30236 & ~n30241;
  assign n30243 = n30242 ^ n30240;
  assign n30245 = n30244 ^ n30243;
  assign n30246 = n28914 ^ n27802;
  assign n30247 = n28914 ^ n28895;
  assign n30248 = ~n30246 & ~n30247;
  assign n30249 = n30248 ^ n27802;
  assign n30250 = n30249 ^ n30244;
  assign n30251 = ~n30245 & n30250;
  assign n30252 = n30251 ^ n30249;
  assign n30253 = n30252 ^ n29860;
  assign n30254 = n29862 & ~n30253;
  assign n30255 = n30254 ^ n29861;
  assign n29853 = n28899 ^ n27790;
  assign n29854 = n28899 ^ n28874;
  assign n29855 = ~n29853 & ~n29854;
  assign n29856 = n29855 ^ n27790;
  assign n30256 = n30255 ^ n29856;
  assign n30257 = n29688 ^ n29668;
  assign n30258 = n30257 ^ n30255;
  assign n30259 = n30256 & n30258;
  assign n30260 = n30259 ^ n30257;
  assign n30261 = n30260 ^ n29849;
  assign n30262 = n29852 & n30261;
  assign n30263 = n30262 ^ n29851;
  assign n30264 = n30263 ^ n29844;
  assign n30265 = ~n29845 & n30264;
  assign n30266 = n30265 ^ n29843;
  assign n30267 = n30266 ^ n29838;
  assign n30268 = n29839 & ~n30267;
  assign n30269 = n30268 ^ n29834;
  assign n29833 = n29707 ^ n29658;
  assign n30270 = n30269 ^ n29833;
  assign n30422 = n30274 ^ n30270;
  assign n30417 = n30266 ^ n29839;
  assign n30411 = n30263 ^ n29843;
  assign n30412 = n30411 ^ n29844;
  assign n30361 = n30260 ^ n29852;
  assign n30362 = n30361 ^ n27303;
  assign n30363 = n30252 ^ n29862;
  assign n30364 = n30363 ^ n27304;
  assign n30365 = n30249 ^ n30245;
  assign n30366 = n30365 ^ n27314;
  assign n30367 = n30240 ^ n30236;
  assign n30368 = n30367 ^ n27317;
  assign n30369 = n30231 ^ n29866;
  assign n30370 = n30369 ^ n30197;
  assign n30371 = n30370 ^ n27193;
  assign n30372 = n30204 ^ n30200;
  assign n30373 = n27336 & n30372;
  assign n30374 = n30373 ^ n27334;
  assign n30375 = n30211 ^ n30210;
  assign n30376 = n30375 ^ n30373;
  assign n30377 = n30374 & n30376;
  assign n30378 = n30377 ^ n27334;
  assign n30379 = n30378 ^ n27375;
  assign n30380 = n30220 ^ n30219;
  assign n30381 = n30380 ^ n30378;
  assign n30382 = ~n30379 & n30381;
  assign n30383 = n30382 ^ n27375;
  assign n30384 = n30383 ^ n27332;
  assign n30385 = n30228 ^ n30199;
  assign n30386 = n30385 ^ n30223;
  assign n30387 = n30386 ^ n30383;
  assign n30388 = ~n30384 & ~n30387;
  assign n30389 = n30388 ^ n27332;
  assign n30390 = n30389 ^ n30370;
  assign n30391 = n30371 & n30390;
  assign n30392 = n30391 ^ n27193;
  assign n30393 = n30392 ^ n30367;
  assign n30394 = ~n30368 & n30393;
  assign n30395 = n30394 ^ n27317;
  assign n30396 = n30395 ^ n30365;
  assign n30397 = n30366 & n30396;
  assign n30398 = n30397 ^ n27314;
  assign n30399 = n30398 ^ n30363;
  assign n30400 = n30364 & ~n30399;
  assign n30401 = n30400 ^ n27304;
  assign n30402 = n30401 ^ n27399;
  assign n30403 = n30257 ^ n29856;
  assign n30404 = n30403 ^ n30255;
  assign n30405 = n30404 ^ n30401;
  assign n30406 = n30402 & n30405;
  assign n30407 = n30406 ^ n27399;
  assign n30408 = n30407 ^ n30361;
  assign n30409 = ~n30362 & ~n30408;
  assign n30410 = n30409 ^ n27303;
  assign n30413 = n30412 ^ n30410;
  assign n30414 = n30412 ^ n27302;
  assign n30415 = n30413 & n30414;
  assign n30416 = n30415 ^ n27302;
  assign n30418 = n30417 ^ n30416;
  assign n30419 = n30417 ^ n27296;
  assign n30420 = n30418 & ~n30419;
  assign n30421 = n30420 ^ n27296;
  assign n30423 = n30422 ^ n30421;
  assign n30424 = n30422 ^ n27290;
  assign n30425 = n30423 & n30424;
  assign n30426 = n30425 ^ n27290;
  assign n30275 = n30274 ^ n29833;
  assign n30276 = n30270 & n30275;
  assign n30277 = n30276 ^ n30274;
  assign n29827 = n28962 ^ n28150;
  assign n29829 = n29828 ^ n28962;
  assign n29830 = n29827 & ~n29829;
  assign n29831 = n29830 ^ n28150;
  assign n29825 = n29710 ^ n1949;
  assign n29826 = n29825 ^ n29652;
  assign n29832 = n29831 ^ n29826;
  assign n30359 = n30277 ^ n29832;
  assign n30360 = n30359 ^ n27430;
  assign n30478 = n30426 ^ n30360;
  assign n30479 = n30423 ^ n27290;
  assign n30480 = n30407 ^ n30362;
  assign n30481 = n30404 ^ n27399;
  assign n30482 = n30481 ^ n30401;
  assign n30483 = n30398 ^ n30364;
  assign n30484 = n30395 ^ n27314;
  assign n30485 = n30484 ^ n30365;
  assign n30486 = n30380 ^ n30379;
  assign n30487 = n30386 ^ n27332;
  assign n30488 = n30487 ^ n30383;
  assign n30489 = ~n30486 & ~n30488;
  assign n30490 = n30389 ^ n27193;
  assign n30491 = n30490 ^ n30370;
  assign n30492 = n30489 & ~n30491;
  assign n30493 = n30392 ^ n27317;
  assign n30494 = n30493 ^ n30367;
  assign n30495 = ~n30492 & n30494;
  assign n30496 = n30485 & ~n30495;
  assign n30497 = ~n30483 & n30496;
  assign n30498 = ~n30482 & ~n30497;
  assign n30499 = ~n30480 & n30498;
  assign n30500 = n30413 ^ n27302;
  assign n30501 = ~n30499 & n30500;
  assign n30502 = n30418 ^ n27296;
  assign n30503 = n30501 & n30502;
  assign n30504 = ~n30479 & n30503;
  assign n30505 = n30478 & n30504;
  assign n30427 = n30426 ^ n30359;
  assign n30428 = n30360 & ~n30427;
  assign n30429 = n30428 ^ n27430;
  assign n30283 = n28956 ^ n27762;
  assign n30284 = n29897 ^ n28956;
  assign n30285 = n30283 & ~n30284;
  assign n30286 = n30285 ^ n27762;
  assign n30281 = n29715 ^ n1964;
  assign n30356 = n30286 ^ n30281;
  assign n30278 = n30277 ^ n29826;
  assign n30279 = ~n29832 & n30278;
  assign n30280 = n30279 ^ n29831;
  assign n30357 = n30356 ^ n30280;
  assign n30358 = n30357 ^ n27531;
  assign n30477 = n30429 ^ n30358;
  assign n30570 = n30505 ^ n30477;
  assign n30574 = n30573 ^ n30570;
  assign n2257 = n2214 ^ n2157;
  assign n2258 = n2257 ^ n2250;
  assign n2262 = n2261 ^ n2258;
  assign n30575 = n30503 ^ n30479;
  assign n30576 = ~n2262 & ~n30575;
  assign n30580 = n30504 ^ n30478;
  assign n30581 = ~n30579 & n30580;
  assign n30582 = ~n30576 & ~n30581;
  assign n30583 = n30502 ^ n30501;
  assign n30584 = n2244 & ~n30583;
  assign n30585 = n30500 ^ n30499;
  assign n30586 = n30585 ^ n2229;
  assign n30592 = n28504 ^ n2038;
  assign n30593 = n30592 ^ n1826;
  assign n30594 = n30593 ^ n2223;
  assign n30595 = n30498 ^ n30480;
  assign n30598 = ~n30594 & n30595;
  assign n30590 = n30497 ^ n30482;
  assign n30591 = n30589 & n30590;
  assign n30596 = n30595 ^ n30594;
  assign n30597 = ~n30591 & ~n30596;
  assign n30599 = n30598 ^ n30597;
  assign n30600 = n30599 ^ n30585;
  assign n30601 = n30586 & n30600;
  assign n30602 = n30601 ^ n2229;
  assign n30603 = ~n30584 & ~n30602;
  assign n30659 = ~n2229 & ~n30585;
  assign n30660 = ~n30589 & ~n30590;
  assign n30661 = ~n30598 & ~n30660;
  assign n30662 = ~n30659 & n30661;
  assign n30604 = n30496 ^ n30483;
  assign n1695 = n1694 ^ n1658;
  assign n1705 = n1704 ^ n1695;
  assign n1709 = n1708 ^ n1705;
  assign n30605 = n30604 ^ n1709;
  assign n30609 = n30495 ^ n30485;
  assign n30610 = n30609 ^ n30608;
  assign n30611 = n28515 ^ n1484;
  assign n30612 = n30611 ^ n25000;
  assign n30613 = n30612 ^ n1609;
  assign n30614 = n30491 ^ n30489;
  assign n30615 = ~n30613 & ~n30614;
  assign n30616 = n30494 ^ n30492;
  assign n30617 = ~n1619 & n30616;
  assign n30618 = ~n30615 & ~n30617;
  assign n30639 = n30488 ^ n30486;
  assign n30619 = n28640 ^ n21370;
  assign n30620 = n30619 ^ n25336;
  assign n30621 = n30620 ^ n20097;
  assign n30622 = n30372 ^ n27336;
  assign n30623 = n30621 & n30622;
  assign n30627 = n30626 ^ n30623;
  assign n30628 = n30375 ^ n30374;
  assign n30629 = n30628 ^ n30626;
  assign n30630 = n30627 & n30629;
  assign n30631 = n30630 ^ n30623;
  assign n30635 = n30634 ^ n30631;
  assign n30636 = n30631 ^ n30486;
  assign n30637 = n30635 & n30636;
  assign n30638 = n30637 ^ n30634;
  assign n30640 = n30639 ^ n30638;
  assign n30644 = n30643 ^ n30639;
  assign n30645 = n30640 & ~n30644;
  assign n30646 = n30645 ^ n30643;
  assign n30647 = n30618 & n30646;
  assign n30648 = n30613 & n30614;
  assign n30649 = n30616 ^ n1619;
  assign n30650 = ~n30648 & ~n30649;
  assign n30651 = n30650 ^ n30617;
  assign n30652 = ~n30647 & n30651;
  assign n30653 = n30652 ^ n30609;
  assign n30654 = n30610 & n30653;
  assign n30655 = n30654 ^ n30608;
  assign n30656 = n30655 ^ n30604;
  assign n30657 = n30605 & ~n30656;
  assign n30658 = n30657 ^ n1709;
  assign n30663 = n30662 ^ n30658;
  assign n30664 = ~n2244 & n30583;
  assign n30665 = n30664 ^ n30662;
  assign n30666 = n30662 & ~n30665;
  assign n30667 = n30666 ^ n30662;
  assign n30668 = n30663 & n30667;
  assign n30669 = n30668 ^ n30666;
  assign n30670 = n30669 ^ n30662;
  assign n30671 = n30670 ^ n30664;
  assign n30672 = n30603 & ~n30671;
  assign n30673 = n30672 ^ n30664;
  assign n30674 = n30582 & ~n30673;
  assign n30675 = n2262 & n30575;
  assign n30676 = n30580 ^ n30579;
  assign n30677 = ~n30675 & ~n30676;
  assign n30678 = n30677 ^ n30581;
  assign n30679 = ~n30674 & n30678;
  assign n30680 = n30679 ^ n30570;
  assign n30681 = n30574 & n30680;
  assign n30682 = n30681 ^ n30573;
  assign n30430 = n30429 ^ n30357;
  assign n30431 = n30358 & ~n30430;
  assign n30432 = n30431 ^ n27531;
  assign n30292 = n28949 ^ n27750;
  assign n30293 = n29896 ^ n28949;
  assign n30294 = n30292 & n30293;
  assign n30295 = n30294 ^ n27750;
  assign n30290 = n29718 ^ n29651;
  assign n30282 = n30281 ^ n30280;
  assign n30287 = n30286 ^ n30280;
  assign n30288 = ~n30282 & ~n30287;
  assign n30289 = n30288 ^ n30281;
  assign n30291 = n30290 ^ n30289;
  assign n30354 = n30295 ^ n30291;
  assign n30355 = n30354 ^ n27699;
  assign n30507 = n30432 ^ n30355;
  assign n30506 = ~n30477 & ~n30505;
  assign n30565 = n30507 ^ n30506;
  assign n30569 = n30568 ^ n30565;
  assign n31398 = n30682 ^ n30569;
  assign n29802 = n29738 ^ n29637;
  assign n32873 = n31398 ^ n29802;
  assign n30898 = n29742 ^ n28891;
  assign n30899 = n30281 ^ n29742;
  assign n30900 = n30898 & ~n30899;
  assign n30901 = n30900 ^ n28891;
  assign n30887 = n30614 ^ n30613;
  assign n30897 = n30887 ^ n30646;
  assign n30902 = n30901 ^ n30897;
  assign n30907 = n30643 ^ n30640;
  assign n30903 = n29591 ^ n28899;
  assign n30904 = n29826 ^ n29591;
  assign n30905 = ~n30903 & ~n30904;
  assign n30906 = n30905 ^ n28899;
  assign n30908 = n30907 ^ n30906;
  assign n30913 = n30622 ^ n30621;
  assign n30909 = n28989 ^ n28882;
  assign n30910 = n29844 ^ n28882;
  assign n30911 = n30909 & n30910;
  assign n30912 = n30911 ^ n28989;
  assign n30914 = n30913 ^ n30912;
  assign n30974 = n28433 ^ n21357;
  assign n30975 = n30974 ^ n2492;
  assign n30976 = n30975 ^ n1547;
  assign n30796 = n30149 ^ n30111;
  assign n30792 = n28663 ^ n28050;
  assign n30793 = n29423 ^ n28663;
  assign n30794 = ~n30792 & n30793;
  assign n30795 = n30794 ^ n28050;
  assign n30797 = n30796 ^ n30795;
  assign n30764 = n30146 ^ n30113;
  assign n30543 = n28686 ^ n28074;
  assign n30544 = n30187 ^ n28686;
  assign n30545 = n30543 & n30544;
  assign n30546 = n30545 ^ n28074;
  assign n30542 = n30143 ^ n30115;
  assign n30547 = n30546 ^ n30542;
  assign n30530 = n28683 ^ n28063;
  assign n30531 = n30047 ^ n28683;
  assign n30532 = n30530 & n30531;
  assign n30533 = n30532 ^ n28063;
  assign n30529 = n30140 ^ n30120;
  assign n30534 = n30533 ^ n30529;
  assign n30468 = n30137 ^ n30134;
  assign n30463 = n29465 ^ n28654;
  assign n30464 = n29972 ^ n29465;
  assign n30465 = n30463 & n30464;
  assign n30466 = n30465 ^ n28654;
  assign n30525 = n30468 ^ n30466;
  assign n30332 = n29408 ^ n28414;
  assign n30333 = n29868 ^ n29408;
  assign n30334 = n30332 & ~n30333;
  assign n30335 = n30334 ^ n28414;
  assign n30331 = n30129 ^ n30125;
  assign n30336 = n30335 ^ n30331;
  assign n29789 = n29249 ^ n28402;
  assign n29791 = n29790 ^ n29249;
  assign n29792 = ~n29789 & n29791;
  assign n29793 = n29792 ^ n28402;
  assign n29769 = n29768 ^ n29765;
  assign n29788 = n29787 ^ n29769;
  assign n29794 = n29793 ^ n29788;
  assign n29796 = n29198 ^ n28180;
  assign n29798 = n29797 ^ n29198;
  assign n29799 = n29796 & n29798;
  assign n29800 = n29799 ^ n28180;
  assign n29795 = n29762 ^ n29759;
  assign n29801 = n29800 ^ n29795;
  assign n29803 = n29086 ^ n27710;
  assign n29805 = n29804 ^ n29086;
  assign n29806 = n29803 & ~n29805;
  assign n29807 = n29806 ^ n27710;
  assign n29808 = n29807 ^ n29802;
  assign n30305 = n29727 ^ n29642;
  assign n29815 = n29724 ^ n29647;
  assign n29810 = n28947 ^ n27739;
  assign n29812 = n29811 ^ n28947;
  assign n29813 = n29810 & n29812;
  assign n29814 = n29813 ^ n27739;
  assign n29816 = n29815 ^ n29814;
  assign n29822 = n29721 ^ n2110;
  assign n29823 = n29822 ^ n29648;
  assign n29817 = n29063 ^ n27747;
  assign n29819 = n29818 ^ n29063;
  assign n29820 = ~n29817 & ~n29819;
  assign n29821 = n29820 ^ n27747;
  assign n29824 = n29823 ^ n29821;
  assign n30296 = n30295 ^ n30290;
  assign n30297 = ~n30291 & ~n30296;
  assign n30298 = n30297 ^ n30295;
  assign n30299 = n30298 ^ n29823;
  assign n30300 = ~n29824 & ~n30299;
  assign n30301 = n30300 ^ n29821;
  assign n30302 = n30301 ^ n29815;
  assign n30303 = n29816 & n30302;
  assign n30304 = n30303 ^ n29814;
  assign n30306 = n30305 ^ n30304;
  assign n30307 = n28941 ^ n27731;
  assign n30308 = n29894 ^ n28941;
  assign n30309 = ~n30307 & ~n30308;
  assign n30310 = n30309 ^ n27731;
  assign n30311 = n30310 ^ n30305;
  assign n30312 = ~n30306 & n30311;
  assign n30313 = n30312 ^ n30310;
  assign n29809 = n29735 ^ n29732;
  assign n30314 = n30313 ^ n29809;
  assign n30315 = n28931 ^ n27717;
  assign n30316 = n29945 ^ n28931;
  assign n30317 = ~n30315 & ~n30316;
  assign n30318 = n30317 ^ n27717;
  assign n30319 = n30318 ^ n29809;
  assign n30320 = n30314 & ~n30319;
  assign n30321 = n30320 ^ n30318;
  assign n30322 = n30321 ^ n29802;
  assign n30323 = ~n29808 & ~n30322;
  assign n30324 = n30323 ^ n29807;
  assign n30325 = n30324 ^ n29800;
  assign n30326 = ~n29801 & ~n30325;
  assign n30327 = n30326 ^ n29795;
  assign n30328 = n30327 ^ n29788;
  assign n30329 = ~n29794 & n30328;
  assign n30330 = n30329 ^ n29793;
  assign n30460 = n30331 ^ n30330;
  assign n30461 = ~n30336 & ~n30460;
  assign n30462 = n30461 ^ n30335;
  assign n30526 = n30468 ^ n30462;
  assign n30527 = ~n30525 & ~n30526;
  assign n30528 = n30527 ^ n30466;
  assign n30548 = n30533 ^ n30528;
  assign n30549 = n30534 & ~n30548;
  assign n30550 = n30549 ^ n30529;
  assign n30761 = n30550 ^ n30546;
  assign n30762 = ~n30547 & n30761;
  assign n30763 = n30762 ^ n30542;
  assign n30765 = n30764 ^ n30763;
  assign n30766 = n28669 ^ n28057;
  assign n30767 = n29433 ^ n28669;
  assign n30768 = n30766 & ~n30767;
  assign n30769 = n30768 ^ n28057;
  assign n30789 = n30769 ^ n30764;
  assign n30790 = n30765 & n30789;
  assign n30791 = n30790 ^ n30769;
  assign n30843 = n30795 ^ n30791;
  assign n30844 = n30797 & ~n30843;
  assign n30845 = n30844 ^ n30796;
  assign n30841 = n30152 ^ n30109;
  assign n30837 = n28661 ^ n28044;
  assign n30838 = n29421 ^ n28661;
  assign n30839 = n30837 & ~n30838;
  assign n30840 = n30839 ^ n28044;
  assign n30842 = n30841 ^ n30840;
  assign n30846 = n30845 ^ n30842;
  assign n30847 = n30846 ^ n27276;
  assign n30798 = n30797 ^ n30791;
  assign n30799 = n30798 ^ n27233;
  assign n30770 = n30769 ^ n30765;
  assign n30771 = n30770 ^ n27186;
  assign n30551 = n30550 ^ n30547;
  assign n30552 = n30551 ^ n27141;
  assign n30535 = n30534 ^ n30528;
  assign n30536 = n30535 ^ n27113;
  assign n30467 = n30466 ^ n30462;
  assign n30469 = n30468 ^ n30467;
  assign n30337 = n30336 ^ n30330;
  assign n30338 = n30337 ^ n27727;
  assign n30339 = n30327 ^ n29793;
  assign n30340 = n30339 ^ n29788;
  assign n30341 = n30340 ^ n27735;
  assign n30342 = n30324 ^ n29801;
  assign n30343 = n30342 ^ n27742;
  assign n30344 = n30321 ^ n29808;
  assign n30345 = n30344 ^ n27752;
  assign n30346 = n30318 ^ n30314;
  assign n30347 = n30346 ^ n27758;
  assign n30348 = n30310 ^ n30306;
  assign n30349 = n30348 ^ n27868;
  assign n30350 = n30301 ^ n29816;
  assign n30351 = n30350 ^ n27765;
  assign n30352 = n30298 ^ n29824;
  assign n30353 = n30352 ^ n27772;
  assign n30433 = n30432 ^ n30354;
  assign n30434 = ~n30355 & n30433;
  assign n30435 = n30434 ^ n27699;
  assign n30436 = n30435 ^ n30352;
  assign n30437 = n30353 & ~n30436;
  assign n30438 = n30437 ^ n27772;
  assign n30439 = n30438 ^ n30350;
  assign n30440 = n30351 & ~n30439;
  assign n30441 = n30440 ^ n27765;
  assign n30442 = n30441 ^ n30348;
  assign n30443 = ~n30349 & n30442;
  assign n30444 = n30443 ^ n27868;
  assign n30445 = n30444 ^ n30346;
  assign n30446 = ~n30347 & ~n30445;
  assign n30447 = n30446 ^ n27758;
  assign n30448 = n30447 ^ n30344;
  assign n30449 = ~n30345 & n30448;
  assign n30450 = n30449 ^ n27752;
  assign n30451 = n30450 ^ n30342;
  assign n30452 = n30343 & ~n30451;
  assign n30453 = n30452 ^ n27742;
  assign n30454 = n30453 ^ n30340;
  assign n30455 = ~n30341 & n30454;
  assign n30456 = n30455 ^ n27735;
  assign n30457 = n30456 ^ n30337;
  assign n30458 = n30338 & n30457;
  assign n30459 = n30458 ^ n27727;
  assign n30470 = n30469 ^ n30459;
  assign n30522 = n30469 ^ n27720;
  assign n30523 = n30470 & ~n30522;
  assign n30524 = n30523 ^ n27720;
  assign n30539 = n30535 ^ n30524;
  assign n30540 = n30536 & n30539;
  assign n30541 = n30540 ^ n27113;
  assign n30772 = n30551 ^ n30541;
  assign n30773 = ~n30552 & n30772;
  assign n30774 = n30773 ^ n27141;
  assign n30786 = n30774 ^ n30770;
  assign n30787 = ~n30771 & ~n30786;
  assign n30788 = n30787 ^ n27186;
  assign n30834 = n30798 ^ n30788;
  assign n30835 = n30799 & ~n30834;
  assign n30836 = n30835 ^ n27233;
  assign n30931 = n30846 ^ n30836;
  assign n30932 = ~n30847 & n30931;
  assign n30933 = n30932 ^ n27276;
  assign n30924 = n28703 ^ n28087;
  assign n30925 = n29415 ^ n28703;
  assign n30926 = ~n30924 & n30925;
  assign n30927 = n30926 ^ n28087;
  assign n30921 = n30845 ^ n30841;
  assign n30922 = ~n30842 & n30921;
  assign n30923 = n30922 ^ n30840;
  assign n30928 = n30927 ^ n30923;
  assign n30919 = n30155 ^ n1130;
  assign n30920 = n30919 ^ n30103;
  assign n30929 = n30928 ^ n30920;
  assign n30930 = n30929 ^ n27351;
  assign n30934 = n30933 ^ n30930;
  assign n30848 = n30847 ^ n30836;
  assign n30800 = n30799 ^ n30788;
  assign n30471 = n30470 ^ n27720;
  assign n30472 = n30456 ^ n27727;
  assign n30473 = n30472 ^ n30337;
  assign n30474 = n30453 ^ n30341;
  assign n30475 = n30450 ^ n30343;
  assign n30476 = n30438 ^ n30351;
  assign n30508 = ~n30506 & ~n30507;
  assign n30509 = n30435 ^ n30353;
  assign n30510 = n30508 & n30509;
  assign n30511 = n30476 & n30510;
  assign n30512 = n30441 ^ n30349;
  assign n30513 = ~n30511 & n30512;
  assign n30514 = n30444 ^ n30347;
  assign n30515 = ~n30513 & ~n30514;
  assign n30516 = n30447 ^ n30345;
  assign n30517 = n30515 & n30516;
  assign n30518 = n30475 & ~n30517;
  assign n30519 = ~n30474 & n30518;
  assign n30520 = n30473 & n30519;
  assign n30521 = ~n30471 & ~n30520;
  assign n30537 = n30536 ^ n30524;
  assign n30538 = n30521 & n30537;
  assign n30553 = n30552 ^ n30541;
  assign n30760 = n30538 & n30553;
  assign n30775 = n30774 ^ n30771;
  assign n30801 = n30760 & n30775;
  assign n30849 = ~n30800 & ~n30801;
  assign n30935 = n30848 & n30849;
  assign n30972 = ~n30934 & n30935;
  assign n30965 = n28737 ^ n27833;
  assign n30966 = n29470 ^ n28737;
  assign n30967 = ~n30965 & n30966;
  assign n30968 = n30967 ^ n27833;
  assign n30961 = n30927 ^ n30920;
  assign n30962 = n30923 ^ n30920;
  assign n30963 = ~n30961 & ~n30962;
  assign n30964 = n30963 ^ n30927;
  assign n30969 = n30968 ^ n30964;
  assign n30960 = n30163 ^ n30160;
  assign n30970 = n30969 ^ n30960;
  assign n30955 = n30933 ^ n27351;
  assign n30956 = n30933 ^ n30929;
  assign n30957 = ~n30955 & n30956;
  assign n30958 = n30957 ^ n27351;
  assign n30959 = n30958 ^ n27346;
  assign n30971 = n30970 ^ n30959;
  assign n30973 = n30972 ^ n30971;
  assign n30977 = n30976 ^ n30973;
  assign n30937 = n28438 ^ n21328;
  assign n30938 = n30937 ^ n25211;
  assign n30939 = n30938 ^ n2486;
  assign n30936 = n30935 ^ n30934;
  assign n30940 = n30939 ^ n30936;
  assign n30683 = n30682 ^ n30565;
  assign n30684 = ~n30569 & n30683;
  assign n30685 = n30684 ^ n30568;
  assign n30689 = n30516 ^ n30515;
  assign n30690 = ~n30688 & n30689;
  assign n30694 = n30517 ^ n30475;
  assign n30695 = ~n30693 & n30694;
  assign n30696 = ~n30690 & ~n30695;
  assign n30700 = n30518 ^ n30474;
  assign n30701 = ~n30699 & n30700;
  assign n645 = n644 ^ n539;
  assign n658 = n657 ^ n645;
  assign n662 = n661 ^ n658;
  assign n30702 = n30512 ^ n30511;
  assign n30703 = ~n662 & n30702;
  assign n30707 = n30509 ^ n30508;
  assign n30708 = ~n30706 & n30707;
  assign n30709 = n30510 ^ n30476;
  assign n30710 = n28477 ^ n21143;
  assign n30711 = n30710 ^ n24965;
  assign n30712 = n30711 ^ n652;
  assign n30713 = n30709 & ~n30712;
  assign n30714 = ~n30708 & ~n30713;
  assign n30715 = n28470 ^ n21136;
  assign n30716 = n30715 ^ n25080;
  assign n30717 = n30716 ^ n564;
  assign n30718 = n30514 ^ n30513;
  assign n30719 = ~n30717 & n30718;
  assign n30720 = n30714 & ~n30719;
  assign n30721 = ~n30703 & n30720;
  assign n1078 = n995 ^ n939;
  assign n1088 = n1087 ^ n1078;
  assign n1089 = n1088 ^ n1071;
  assign n30722 = n30519 ^ n30473;
  assign n30723 = ~n1089 & ~n30722;
  assign n30724 = n30721 & ~n30723;
  assign n30725 = ~n30701 & n30724;
  assign n30726 = n30696 & n30725;
  assign n30727 = n30685 & n30726;
  assign n30728 = n30722 ^ n1089;
  assign n30729 = n30718 ^ n30717;
  assign n30730 = n30702 ^ n662;
  assign n30731 = n30712 ^ n30709;
  assign n30732 = n30706 & ~n30707;
  assign n30733 = ~n30731 & ~n30732;
  assign n30734 = n30733 ^ n30713;
  assign n30735 = n30734 ^ n30702;
  assign n30736 = ~n30730 & ~n30735;
  assign n30737 = n30736 ^ n662;
  assign n30738 = ~n30729 & ~n30737;
  assign n30739 = n30738 ^ n30719;
  assign n30740 = n30696 & ~n30739;
  assign n30741 = n30688 & ~n30689;
  assign n30742 = n30694 ^ n30693;
  assign n30743 = ~n30741 & ~n30742;
  assign n30744 = n30743 ^ n30695;
  assign n30745 = ~n30740 & n30744;
  assign n30746 = n30699 & ~n30700;
  assign n30747 = ~n30701 & ~n30746;
  assign n30748 = ~n30745 & n30747;
  assign n30749 = n30748 ^ n30746;
  assign n30750 = n30749 ^ n30722;
  assign n30751 = n30728 & ~n30750;
  assign n30752 = n30751 ^ n1089;
  assign n30753 = ~n30727 & ~n30752;
  assign n1232 = n1219 ^ n1138;
  assign n1233 = n1232 ^ n1106;
  assign n1237 = n1236 ^ n1233;
  assign n30560 = n30537 ^ n30521;
  assign n30563 = ~n1237 & n30560;
  assign n30558 = n30520 ^ n30471;
  assign n30754 = ~n1097 & n30558;
  assign n30755 = ~n30563 & ~n30754;
  assign n1247 = n1228 ^ n1153;
  assign n1248 = n1247 ^ n1244;
  assign n1252 = n1251 ^ n1248;
  assign n30554 = n30553 ^ n30538;
  assign n30555 = ~n1252 & n30554;
  assign n2297 = n2273 ^ n1329;
  assign n2301 = n2300 ^ n2297;
  assign n2302 = n2301 ^ n2289;
  assign n30776 = n30775 ^ n30760;
  assign n30807 = ~n2302 & n30776;
  assign n30808 = ~n30555 & ~n30807;
  assign n30809 = n30755 & n30808;
  assign n30810 = ~n30753 & n30809;
  assign n30777 = n30776 ^ n2302;
  assign n30556 = n1252 & ~n30554;
  assign n30557 = ~n30555 & ~n30556;
  assign n30559 = n1097 & ~n30558;
  assign n30561 = n30560 ^ n1237;
  assign n30562 = ~n30559 & ~n30561;
  assign n30564 = n30563 ^ n30562;
  assign n30811 = n30557 & n30564;
  assign n30812 = n30811 ^ n30555;
  assign n30813 = n30812 ^ n30776;
  assign n30814 = ~n30777 & ~n30813;
  assign n30815 = n30814 ^ n2302;
  assign n30816 = ~n30810 & ~n30815;
  assign n2364 = n2363 ^ n2324;
  assign n2365 = n2364 ^ n2357;
  assign n2369 = n2368 ^ n2365;
  assign n30850 = n30849 ^ n30848;
  assign n30851 = ~n2369 & ~n30850;
  assign n30802 = n30801 ^ n30800;
  assign n30803 = n28625 ^ n21278;
  assign n30804 = n30803 ^ n2295;
  assign n30805 = n30804 ^ n2348;
  assign n30941 = ~n30802 & ~n30805;
  assign n30942 = ~n30851 & ~n30941;
  assign n30943 = ~n30816 & n30942;
  assign n30944 = n30943 ^ n30936;
  assign n30945 = n30944 ^ n30936;
  assign n30852 = n2369 & n30850;
  assign n30853 = ~n30851 & ~n30852;
  assign n30946 = n30802 & n30805;
  assign n30947 = n30853 & n30946;
  assign n30948 = n30947 ^ n30852;
  assign n30949 = n30948 ^ n30936;
  assign n30950 = n30949 ^ n30936;
  assign n30951 = ~n30945 & ~n30950;
  assign n30952 = n30951 ^ n30936;
  assign n30953 = ~n30940 & ~n30952;
  assign n30954 = n30953 ^ n30939;
  assign n30978 = n30977 ^ n30954;
  assign n30915 = n28999 ^ n28895;
  assign n30916 = n29851 ^ n28895;
  assign n30917 = n30915 & ~n30916;
  assign n30918 = n30917 ^ n28999;
  assign n30979 = n30978 ^ n30918;
  assign n30985 = n28922 ^ n28897;
  assign n30986 = n30257 ^ n28897;
  assign n30987 = ~n30985 & n30986;
  assign n30988 = n30987 ^ n28922;
  assign n30980 = n30850 ^ n2369;
  assign n30806 = n30805 ^ n30802;
  assign n30831 = n30816 ^ n30802;
  assign n30832 = n30806 & n30831;
  assign n30833 = n30832 ^ n30805;
  assign n30981 = n30850 ^ n30833;
  assign n30982 = n30980 & ~n30981;
  assign n30983 = n30982 ^ n2369;
  assign n30984 = n30983 ^ n30940;
  assign n30989 = n30988 ^ n30984;
  assign n30855 = n28904 ^ n28853;
  assign n30856 = n29861 ^ n28904;
  assign n30857 = n30855 & ~n30856;
  assign n30858 = n30857 ^ n28853;
  assign n30854 = n30853 ^ n30833;
  assign n30859 = n30858 ^ n30854;
  assign n30756 = ~n30753 & n30755;
  assign n30757 = n30564 & ~n30756;
  assign n30758 = n30557 & ~n30757;
  assign n30759 = n30758 ^ n30556;
  assign n30778 = n30777 ^ n30759;
  assign n30779 = n28919 ^ n28752;
  assign n30780 = n30235 ^ n28919;
  assign n30781 = ~n30779 & n30780;
  assign n30782 = n30781 ^ n28752;
  assign n30822 = ~n30778 & ~n30782;
  assign n30818 = n28912 ^ n28771;
  assign n30819 = n30244 ^ n28912;
  assign n30820 = ~n30818 & ~n30819;
  assign n30821 = n30820 ^ n28771;
  assign n30823 = n30822 ^ n30821;
  assign n30817 = n30816 ^ n30806;
  assign n30828 = n30821 ^ n30817;
  assign n30829 = ~n30823 & ~n30828;
  assign n30830 = n30829 ^ n30822;
  assign n30990 = n30854 ^ n30830;
  assign n30991 = n30859 & ~n30990;
  assign n30992 = n30991 ^ n30858;
  assign n30993 = n30992 ^ n30984;
  assign n30994 = ~n30989 & n30993;
  assign n30995 = n30994 ^ n30988;
  assign n30996 = n30995 ^ n30978;
  assign n30997 = ~n30979 & ~n30996;
  assign n30998 = n30997 ^ n30918;
  assign n30999 = n30998 ^ n30913;
  assign n31000 = ~n30914 & n30999;
  assign n31001 = n31000 ^ n30912;
  assign n31002 = n30628 ^ n30627;
  assign n31003 = n28914 ^ n28874;
  assign n31004 = n29834 ^ n28874;
  assign n31005 = ~n31003 & n31004;
  assign n31006 = n31005 ^ n28914;
  assign n31007 = n31002 & n31006;
  assign n31008 = n30634 ^ n30486;
  assign n31009 = n31008 ^ n30631;
  assign n31010 = n28906 ^ n28867;
  assign n31011 = n29833 ^ n28867;
  assign n31012 = ~n31010 & n31011;
  assign n31013 = n31012 ^ n28906;
  assign n31014 = n31009 & ~n31013;
  assign n31015 = ~n31007 & ~n31014;
  assign n31016 = ~n31001 & n31015;
  assign n31017 = n31013 ^ n31009;
  assign n31018 = ~n31002 & ~n31006;
  assign n31019 = n31018 ^ n31013;
  assign n31020 = ~n31017 & ~n31019;
  assign n31021 = n31020 ^ n31009;
  assign n31022 = ~n31016 & n31021;
  assign n31023 = n31022 ^ n30907;
  assign n31024 = ~n30908 & ~n31023;
  assign n31025 = n31024 ^ n30906;
  assign n31026 = n31025 ^ n30897;
  assign n31027 = ~n30902 & ~n31026;
  assign n31028 = n31027 ^ n30901;
  assign n30892 = n29781 ^ n28885;
  assign n30893 = n30290 ^ n29781;
  assign n30894 = n30892 & ~n30893;
  assign n30895 = n30894 ^ n28885;
  assign n30888 = n30646 ^ n30614;
  assign n30889 = n30887 & ~n30888;
  assign n30890 = n30889 ^ n30613;
  assign n30891 = n30890 ^ n30649;
  assign n30896 = n30895 ^ n30891;
  assign n31045 = n31028 ^ n30896;
  assign n31046 = n31045 ^ n27783;
  assign n31047 = n31025 ^ n30902;
  assign n31048 = n31047 ^ n28132;
  assign n31049 = n31022 ^ n30908;
  assign n31050 = n31049 ^ n27790;
  assign n31051 = n31006 ^ n31002;
  assign n31052 = n31002 ^ n31001;
  assign n31053 = n31051 & ~n31052;
  assign n31054 = n31053 ^ n31006;
  assign n31055 = n31054 ^ n31017;
  assign n31056 = n31055 ^ n27796;
  assign n31057 = n31051 ^ n31001;
  assign n31058 = n31057 ^ n27802;
  assign n31059 = n30998 ^ n30914;
  assign n31060 = n31059 ^ n27808;
  assign n31061 = n30995 ^ n30979;
  assign n31062 = n31061 ^ n27815;
  assign n31063 = n30992 ^ n30989;
  assign n31064 = n31063 ^ n27821;
  assign n30860 = n30859 ^ n30830;
  assign n30861 = n30860 ^ n27286;
  assign n30783 = n30782 ^ n30778;
  assign n30784 = n27192 & n30783;
  assign n30785 = n30784 ^ n28102;
  assign n30824 = n30823 ^ n30817;
  assign n30825 = n30824 ^ n30784;
  assign n30826 = n30785 & ~n30825;
  assign n30827 = n30826 ^ n28102;
  assign n31065 = n30860 ^ n30827;
  assign n31066 = n30861 & ~n31065;
  assign n31067 = n31066 ^ n27286;
  assign n31068 = n31067 ^ n31063;
  assign n31069 = ~n31064 & n31068;
  assign n31070 = n31069 ^ n27821;
  assign n31071 = n31070 ^ n31061;
  assign n31072 = n31062 & n31071;
  assign n31073 = n31072 ^ n27815;
  assign n31074 = n31073 ^ n31059;
  assign n31075 = n31060 & n31074;
  assign n31076 = n31075 ^ n27808;
  assign n31077 = n31076 ^ n31057;
  assign n31078 = ~n31058 & n31077;
  assign n31079 = n31078 ^ n27802;
  assign n31080 = n31079 ^ n31055;
  assign n31081 = n31056 & ~n31080;
  assign n31082 = n31081 ^ n27796;
  assign n31083 = n31082 ^ n31049;
  assign n31084 = ~n31050 & ~n31083;
  assign n31085 = n31084 ^ n27790;
  assign n31086 = n31085 ^ n31047;
  assign n31087 = n31048 & ~n31086;
  assign n31088 = n31087 ^ n28132;
  assign n31089 = n31088 ^ n31045;
  assign n31090 = n31046 & ~n31089;
  assign n31091 = n31090 ^ n27783;
  assign n31029 = n31028 ^ n30891;
  assign n31030 = n30896 & ~n31029;
  assign n31031 = n31030 ^ n30895;
  assign n30882 = n29828 ^ n28876;
  assign n30883 = n29828 ^ n29823;
  assign n30884 = n30882 & ~n30883;
  assign n30885 = n30884 ^ n28876;
  assign n30881 = n30652 ^ n30610;
  assign n30886 = n30885 ^ n30881;
  assign n31043 = n31031 ^ n30886;
  assign n31044 = n31043 ^ n27776;
  assign n31096 = n31091 ^ n31044;
  assign n31097 = n31088 ^ n31046;
  assign n31098 = n31085 ^ n31048;
  assign n31099 = n31076 ^ n31058;
  assign n31100 = n31073 ^ n31060;
  assign n30862 = n30861 ^ n30827;
  assign n31101 = n31067 ^ n31064;
  assign n31102 = ~n30862 & n31101;
  assign n31103 = n31070 ^ n31062;
  assign n31104 = n31102 & ~n31103;
  assign n31105 = ~n31100 & ~n31104;
  assign n31106 = n31099 & ~n31105;
  assign n31107 = n31079 ^ n31056;
  assign n31108 = n31106 & ~n31107;
  assign n31109 = n31082 ^ n31050;
  assign n31110 = ~n31108 & ~n31109;
  assign n31111 = ~n31098 & n31110;
  assign n31112 = n31097 & ~n31111;
  assign n31113 = ~n31096 & n31112;
  assign n31092 = n31091 ^ n31043;
  assign n31093 = ~n31044 & n31092;
  assign n31094 = n31093 ^ n27776;
  assign n31036 = n29897 ^ n28870;
  assign n31037 = n29897 ^ n29815;
  assign n31038 = ~n31036 & ~n31037;
  assign n31039 = n31038 ^ n28870;
  assign n31035 = n30655 ^ n30605;
  assign n31040 = n31039 ^ n31035;
  assign n31032 = n31031 ^ n30881;
  assign n31033 = ~n30886 & ~n31032;
  assign n31034 = n31033 ^ n30885;
  assign n31041 = n31040 ^ n31034;
  assign n31042 = n31041 ^ n27769;
  assign n31095 = n31094 ^ n31042;
  assign n31209 = n31113 ^ n31095;
  assign n31213 = n31212 ^ n31209;
  assign n31214 = n31112 ^ n31096;
  assign n31215 = n31214 ^ n2087;
  assign n31216 = n31111 ^ n31097;
  assign n31220 = n31219 ^ n31216;
  assign n31221 = n31110 ^ n31098;
  assign n1912 = n1908 ^ n1839;
  assign n1919 = n1918 ^ n1912;
  assign n1923 = n1922 ^ n1919;
  assign n31222 = n31221 ^ n1923;
  assign n31223 = n31109 ^ n31108;
  assign n31224 = n31223 ^ n1810;
  assign n31225 = n31107 ^ n31106;
  assign n1778 = n1765 ^ n1729;
  assign n1791 = n1790 ^ n1778;
  assign n1795 = n1794 ^ n1791;
  assign n31226 = n31225 ^ n1795;
  assign n31230 = n31105 ^ n31099;
  assign n31231 = n31230 ^ n31229;
  assign n31235 = n31104 ^ n31100;
  assign n31236 = n31235 ^ n31234;
  assign n31237 = n31103 ^ n31102;
  assign n31241 = n31240 ^ n31237;
  assign n31242 = n31101 ^ n30862;
  assign n31246 = n31245 ^ n31242;
  assign n30872 = n28811 ^ n21568;
  assign n30873 = n30872 ^ n2654;
  assign n30874 = n30873 ^ n1523;
  assign n30867 = n29449 ^ n1550;
  assign n30868 = n30867 ^ n2555;
  assign n30869 = n30868 ^ n2652;
  assign n30870 = n30783 ^ n27192;
  assign n30871 = n30869 & n30870;
  assign n30875 = n30874 ^ n30871;
  assign n30876 = n30824 ^ n30785;
  assign n30877 = n30876 ^ n30874;
  assign n30878 = n30875 & ~n30877;
  assign n30879 = n30878 ^ n30871;
  assign n31247 = n30879 ^ n30862;
  assign n30863 = n28816 ^ n21572;
  assign n30864 = n30863 ^ n1556;
  assign n30865 = n30864 ^ n20253;
  assign n31248 = n30879 ^ n30865;
  assign n31249 = ~n31247 & ~n31248;
  assign n31250 = n31249 ^ n30862;
  assign n31251 = n31250 ^ n31242;
  assign n31252 = n31246 & n31251;
  assign n31253 = n31252 ^ n31245;
  assign n31254 = n31253 ^ n31237;
  assign n31255 = n31241 & ~n31254;
  assign n31256 = n31255 ^ n31240;
  assign n31257 = n31256 ^ n31235;
  assign n31258 = n31236 & ~n31257;
  assign n31259 = n31258 ^ n31234;
  assign n31260 = n31259 ^ n31230;
  assign n31261 = n31231 & ~n31260;
  assign n31262 = n31261 ^ n31229;
  assign n31263 = n31262 ^ n31225;
  assign n31264 = n31226 & ~n31263;
  assign n31265 = n31264 ^ n1795;
  assign n31266 = n31265 ^ n31223;
  assign n31267 = n31224 & ~n31266;
  assign n31268 = n31267 ^ n1810;
  assign n31269 = n31268 ^ n31221;
  assign n31270 = ~n31222 & n31269;
  assign n31271 = n31270 ^ n1923;
  assign n31272 = n31271 ^ n31216;
  assign n31273 = n31220 & ~n31272;
  assign n31274 = n31273 ^ n31219;
  assign n31275 = n31274 ^ n31214;
  assign n31276 = n31215 & ~n31275;
  assign n31277 = n31276 ^ n2087;
  assign n31278 = n31277 ^ n31209;
  assign n31279 = n31213 & ~n31278;
  assign n31280 = n31279 ^ n31212;
  assign n31125 = n31035 ^ n31034;
  assign n31126 = ~n31040 & ~n31125;
  assign n31127 = n31126 ^ n31039;
  assign n31122 = n30590 ^ n30589;
  assign n31123 = n31122 ^ n30658;
  assign n31118 = n29896 ^ n28962;
  assign n31119 = n30305 ^ n29896;
  assign n31120 = ~n31118 & n31119;
  assign n31121 = n31120 ^ n28962;
  assign n31124 = n31123 ^ n31121;
  assign n31128 = n31127 ^ n31124;
  assign n31129 = n31128 ^ n28150;
  assign n31115 = n31094 ^ n31041;
  assign n31116 = ~n31042 & ~n31115;
  assign n31117 = n31116 ^ n27769;
  assign n31130 = n31129 ^ n31117;
  assign n31114 = ~n31095 & n31113;
  assign n31204 = n31130 ^ n31114;
  assign n31208 = n31207 ^ n31204;
  assign n32019 = n31280 ^ n31208;
  assign n32874 = n32019 ^ n31398;
  assign n32875 = ~n32873 & ~n32874;
  assign n32876 = n32875 ^ n29802;
  assign n31333 = n30870 ^ n30869;
  assign n31329 = n29833 ^ n28882;
  assign n31330 = n30891 ^ n29833;
  assign n31331 = ~n31329 & n31330;
  assign n31332 = n31331 ^ n28882;
  assign n31334 = n31333 ^ n31332;
  assign n31704 = n29834 ^ n28895;
  assign n31705 = n30897 ^ n29834;
  assign n31706 = n31704 & n31705;
  assign n31707 = n31706 ^ n28895;
  assign n31537 = n30558 ^ n1097;
  assign n31538 = n31537 ^ n30753;
  assign n31533 = n29470 ^ n28661;
  assign n31534 = n30220 ^ n29470;
  assign n31535 = ~n31533 & n31534;
  assign n31536 = n31535 ^ n28661;
  assign n31539 = n31538 ^ n31536;
  assign n31339 = n30685 & n30721;
  assign n31340 = n30739 & ~n31339;
  assign n31341 = n30696 & ~n31340;
  assign n31342 = n30744 & ~n31341;
  assign n31463 = n30747 & ~n31342;
  assign n31464 = n31463 ^ n30746;
  assign n31465 = n31464 ^ n30728;
  assign n31459 = n29415 ^ n28663;
  assign n31460 = n30211 ^ n29415;
  assign n31461 = n31459 & n31460;
  assign n31462 = n31461 ^ n28663;
  assign n31466 = n31465 ^ n31462;
  assign n31343 = n31342 ^ n30699;
  assign n31344 = n31343 ^ n30700;
  assign n31335 = n29421 ^ n28669;
  assign n31336 = n30200 ^ n29421;
  assign n31337 = n31335 & n31336;
  assign n31338 = n31337 ^ n28669;
  assign n31345 = n31344 ^ n31338;
  assign n31351 = n29423 ^ n28686;
  assign n31352 = n30960 ^ n29423;
  assign n31353 = n31351 & n31352;
  assign n31354 = n31353 ^ n28686;
  assign n31346 = n30689 ^ n30688;
  assign n31347 = n31340 ^ n30689;
  assign n31348 = ~n31346 & ~n31347;
  assign n31349 = n31348 ^ n30688;
  assign n31350 = n31349 ^ n30742;
  assign n31355 = n31354 ^ n31350;
  assign n31357 = n29433 ^ n28683;
  assign n31358 = n30920 ^ n29433;
  assign n31359 = ~n31357 & ~n31358;
  assign n31360 = n31359 ^ n28683;
  assign n31356 = n31346 ^ n31340;
  assign n31361 = n31360 ^ n31356;
  assign n31369 = n30187 ^ n29465;
  assign n31370 = n30841 ^ n30187;
  assign n31371 = n31369 & ~n31370;
  assign n31372 = n31371 ^ n29465;
  assign n31362 = n30685 & n30714;
  assign n31363 = n30734 & ~n31362;
  assign n31364 = n31363 ^ n30702;
  assign n31365 = ~n30730 & ~n31364;
  assign n31366 = n31365 ^ n662;
  assign n31367 = n31366 ^ n30717;
  assign n31368 = n31367 ^ n30718;
  assign n31373 = n31372 ^ n31368;
  assign n31375 = n30047 ^ n29408;
  assign n31376 = n30796 ^ n30047;
  assign n31377 = n31375 & ~n31376;
  assign n31378 = n31377 ^ n29408;
  assign n31374 = n31363 ^ n30730;
  assign n31379 = n31378 ^ n31374;
  assign n31291 = n30707 ^ n30706;
  assign n31384 = n30707 ^ n30685;
  assign n31385 = ~n31291 & n31384;
  assign n31386 = n31385 ^ n30706;
  assign n31387 = n31386 ^ n30731;
  assign n31380 = n29972 ^ n29249;
  assign n31381 = n30764 ^ n29972;
  assign n31382 = n31380 & ~n31381;
  assign n31383 = n31382 ^ n29249;
  assign n31388 = n31387 ^ n31383;
  assign n31389 = n29868 ^ n29198;
  assign n31390 = n30542 ^ n29868;
  assign n31391 = n31389 & n31390;
  assign n31392 = n31391 ^ n29198;
  assign n31292 = n31291 ^ n30685;
  assign n31393 = n31392 ^ n31292;
  assign n31394 = n29790 ^ n29086;
  assign n31395 = n30529 ^ n29790;
  assign n31396 = ~n31394 & ~n31395;
  assign n31397 = n31396 ^ n29086;
  assign n31399 = n31398 ^ n31397;
  assign n31404 = n30679 ^ n30574;
  assign n31400 = n29797 ^ n28931;
  assign n31401 = n30468 ^ n29797;
  assign n31402 = ~n31400 & n31401;
  assign n31403 = n31402 ^ n28931;
  assign n31405 = n31404 ^ n31403;
  assign n31410 = n30575 ^ n2262;
  assign n31411 = n30673 ^ n30575;
  assign n31412 = n31410 & n31411;
  assign n31413 = n31412 ^ n2262;
  assign n31414 = n31413 ^ n30579;
  assign n31415 = n31414 ^ n30580;
  assign n31406 = n29804 ^ n28941;
  assign n31407 = n30331 ^ n29804;
  assign n31408 = n31406 & n31407;
  assign n31409 = n31408 ^ n28941;
  assign n31416 = n31415 ^ n31409;
  assign n31421 = n31410 ^ n30673;
  assign n31417 = n29945 ^ n28947;
  assign n31418 = n29945 ^ n29788;
  assign n31419 = ~n31417 & ~n31418;
  assign n31420 = n31419 ^ n28947;
  assign n31422 = n31421 ^ n31420;
  assign n31183 = n30583 ^ n2244;
  assign n31162 = n30658 & n30661;
  assign n31163 = n30599 & ~n31162;
  assign n31180 = n31163 ^ n30585;
  assign n31181 = n30586 & n31180;
  assign n31182 = n31181 ^ n2229;
  assign n31184 = n31183 ^ n31182;
  assign n31176 = n29894 ^ n29063;
  assign n31177 = n29894 ^ n29795;
  assign n31178 = ~n31176 & n31177;
  assign n31179 = n31178 ^ n29063;
  assign n31185 = n31184 ^ n31179;
  assign n31164 = n31163 ^ n30586;
  assign n31158 = n29811 ^ n28949;
  assign n31159 = n29811 ^ n29802;
  assign n31160 = ~n31158 & n31159;
  assign n31161 = n31160 ^ n28949;
  assign n31165 = n31164 ^ n31161;
  assign n31142 = n30658 ^ n30590;
  assign n31143 = n31122 & ~n31142;
  assign n31144 = n31143 ^ n30589;
  assign n31145 = n31144 ^ n30594;
  assign n31146 = n31145 ^ n30595;
  assign n31138 = n29818 ^ n28956;
  assign n31139 = n29818 ^ n29809;
  assign n31140 = n31138 & n31139;
  assign n31141 = n31140 ^ n28956;
  assign n31147 = n31146 ^ n31141;
  assign n31135 = n31127 ^ n31123;
  assign n31136 = n31124 & n31135;
  assign n31137 = n31136 ^ n31121;
  assign n31155 = n31146 ^ n31137;
  assign n31156 = ~n31147 & n31155;
  assign n31157 = n31156 ^ n31141;
  assign n31173 = n31164 ^ n31157;
  assign n31174 = ~n31165 & n31173;
  assign n31175 = n31174 ^ n31161;
  assign n31423 = n31184 ^ n31175;
  assign n31424 = ~n31185 & n31423;
  assign n31425 = n31424 ^ n31179;
  assign n31426 = n31425 ^ n31421;
  assign n31427 = ~n31422 & n31426;
  assign n31428 = n31427 ^ n31420;
  assign n31429 = n31428 ^ n31415;
  assign n31430 = n31416 & n31429;
  assign n31431 = n31430 ^ n31409;
  assign n31432 = n31431 ^ n31404;
  assign n31433 = n31405 & ~n31432;
  assign n31434 = n31433 ^ n31403;
  assign n31435 = n31434 ^ n31398;
  assign n31436 = n31399 & ~n31435;
  assign n31437 = n31436 ^ n31397;
  assign n31438 = n31437 ^ n31292;
  assign n31439 = n31393 & ~n31438;
  assign n31440 = n31439 ^ n31392;
  assign n31441 = n31440 ^ n31387;
  assign n31442 = n31388 & ~n31441;
  assign n31443 = n31442 ^ n31383;
  assign n31444 = n31443 ^ n31374;
  assign n31445 = ~n31379 & n31444;
  assign n31446 = n31445 ^ n31378;
  assign n31447 = n31446 ^ n31368;
  assign n31448 = ~n31373 & ~n31447;
  assign n31449 = n31448 ^ n31372;
  assign n31450 = n31449 ^ n31356;
  assign n31451 = n31361 & ~n31450;
  assign n31452 = n31451 ^ n31360;
  assign n31453 = n31452 ^ n31350;
  assign n31454 = n31355 & n31453;
  assign n31455 = n31454 ^ n31354;
  assign n31456 = n31455 ^ n31344;
  assign n31457 = ~n31345 & n31456;
  assign n31458 = n31457 ^ n31338;
  assign n31530 = n31465 ^ n31458;
  assign n31531 = n31466 & n31530;
  assign n31532 = n31531 ^ n31462;
  assign n31540 = n31539 ^ n31532;
  assign n31541 = n31540 ^ n28044;
  assign n31467 = n31466 ^ n31458;
  assign n31468 = n31467 ^ n28050;
  assign n31469 = n31455 ^ n31345;
  assign n31470 = n31469 ^ n28057;
  assign n31471 = n31452 ^ n31355;
  assign n31472 = n31471 ^ n28074;
  assign n31473 = n31449 ^ n31361;
  assign n31474 = n31473 ^ n28063;
  assign n31475 = n31446 ^ n31373;
  assign n31476 = n31475 ^ n28654;
  assign n31477 = n31443 ^ n31379;
  assign n31478 = n31477 ^ n28414;
  assign n31479 = n31440 ^ n31388;
  assign n31480 = n31479 ^ n28402;
  assign n31481 = n31437 ^ n31393;
  assign n31482 = n31481 ^ n28180;
  assign n31483 = n31434 ^ n31399;
  assign n31484 = n31483 ^ n27710;
  assign n31485 = n31431 ^ n31405;
  assign n31486 = n31485 ^ n27717;
  assign n31487 = n31428 ^ n31416;
  assign n31488 = n31487 ^ n27731;
  assign n31489 = n31425 ^ n31422;
  assign n31490 = n31489 ^ n27739;
  assign n31186 = n31185 ^ n31175;
  assign n31187 = n31186 ^ n27747;
  assign n31166 = n31165 ^ n31157;
  assign n31167 = n31166 ^ n27750;
  assign n31148 = n31147 ^ n31137;
  assign n31149 = n31148 ^ n27762;
  assign n31132 = n31128 ^ n31117;
  assign n31133 = ~n31129 & n31132;
  assign n31134 = n31133 ^ n28150;
  assign n31152 = n31148 ^ n31134;
  assign n31153 = ~n31149 & n31152;
  assign n31154 = n31153 ^ n27762;
  assign n31170 = n31166 ^ n31154;
  assign n31171 = ~n31167 & n31170;
  assign n31172 = n31171 ^ n27750;
  assign n31491 = n31186 ^ n31172;
  assign n31492 = n31187 & n31491;
  assign n31493 = n31492 ^ n27747;
  assign n31494 = n31493 ^ n31489;
  assign n31495 = ~n31490 & ~n31494;
  assign n31496 = n31495 ^ n27739;
  assign n31497 = n31496 ^ n31487;
  assign n31498 = n31488 & ~n31497;
  assign n31499 = n31498 ^ n27731;
  assign n31500 = n31499 ^ n31485;
  assign n31501 = ~n31486 & n31500;
  assign n31502 = n31501 ^ n27717;
  assign n31503 = n31502 ^ n31483;
  assign n31504 = n31484 & n31503;
  assign n31505 = n31504 ^ n27710;
  assign n31506 = n31505 ^ n31481;
  assign n31507 = n31482 & ~n31506;
  assign n31508 = n31507 ^ n28180;
  assign n31509 = n31508 ^ n31479;
  assign n31510 = ~n31480 & ~n31509;
  assign n31511 = n31510 ^ n28402;
  assign n31512 = n31511 ^ n31477;
  assign n31513 = ~n31478 & ~n31512;
  assign n31514 = n31513 ^ n28414;
  assign n31515 = n31514 ^ n31475;
  assign n31516 = n31476 & n31515;
  assign n31517 = n31516 ^ n28654;
  assign n31518 = n31517 ^ n31473;
  assign n31519 = n31474 & ~n31518;
  assign n31520 = n31519 ^ n28063;
  assign n31521 = n31520 ^ n31471;
  assign n31522 = ~n31472 & ~n31521;
  assign n31523 = n31522 ^ n28074;
  assign n31524 = n31523 ^ n31469;
  assign n31525 = ~n31470 & n31524;
  assign n31526 = n31525 ^ n28057;
  assign n31527 = n31526 ^ n31467;
  assign n31528 = n31468 & ~n31527;
  assign n31529 = n31528 ^ n28050;
  assign n31542 = n31541 ^ n31529;
  assign n31543 = n31523 ^ n31470;
  assign n31544 = n31505 ^ n31482;
  assign n31545 = n31499 ^ n31486;
  assign n31546 = n31496 ^ n31488;
  assign n31547 = n31493 ^ n31490;
  assign n31131 = n31114 & n31130;
  assign n31150 = n31149 ^ n31134;
  assign n31151 = ~n31131 & ~n31150;
  assign n31168 = n31167 ^ n31154;
  assign n31169 = ~n31151 & n31168;
  assign n31188 = n31187 ^ n31172;
  assign n31548 = n31169 & ~n31188;
  assign n31549 = ~n31547 & n31548;
  assign n31550 = n31546 & ~n31549;
  assign n31551 = n31545 & ~n31550;
  assign n31552 = n31502 ^ n31484;
  assign n31553 = n31551 & ~n31552;
  assign n31554 = ~n31544 & ~n31553;
  assign n31555 = n31508 ^ n31480;
  assign n31556 = n31554 & n31555;
  assign n31557 = n31511 ^ n31478;
  assign n31558 = n31556 & ~n31557;
  assign n31559 = n31514 ^ n31476;
  assign n31560 = ~n31558 & n31559;
  assign n31561 = n31517 ^ n31474;
  assign n31562 = n31560 & ~n31561;
  assign n31563 = n31520 ^ n31472;
  assign n31564 = n31562 & n31563;
  assign n31565 = ~n31543 & n31564;
  assign n31566 = n31526 ^ n31468;
  assign n31567 = ~n31565 & ~n31566;
  assign n31568 = ~n31542 & n31567;
  assign n31581 = n31538 ^ n31532;
  assign n31582 = ~n31539 & ~n31581;
  assign n31583 = n31582 ^ n31536;
  assign n31576 = n30753 ^ n30558;
  assign n31577 = ~n31537 & ~n31576;
  assign n31578 = n31577 ^ n1097;
  assign n31579 = n31578 ^ n30561;
  assign n31572 = n28920 ^ n28703;
  assign n31573 = n30199 ^ n28920;
  assign n31574 = ~n31572 & n31573;
  assign n31575 = n31574 ^ n28703;
  assign n31580 = n31579 ^ n31575;
  assign n31584 = n31583 ^ n31580;
  assign n31585 = n31584 ^ n28087;
  assign n31569 = n31540 ^ n31529;
  assign n31570 = n31541 & ~n31569;
  assign n31571 = n31570 ^ n28044;
  assign n31586 = n31585 ^ n31571;
  assign n31700 = n31568 & n31586;
  assign n31694 = n30757 ^ n1252;
  assign n31695 = n31694 ^ n30554;
  assign n31690 = n29482 ^ n28737;
  assign n31691 = n30197 ^ n29482;
  assign n31692 = ~n31690 & n31691;
  assign n31693 = n31692 ^ n28737;
  assign n31696 = n31695 ^ n31693;
  assign n31687 = n31583 ^ n31579;
  assign n31688 = n31580 & ~n31687;
  assign n31689 = n31688 ^ n31575;
  assign n31697 = n31696 ^ n31689;
  assign n31698 = n31697 ^ n27833;
  assign n31683 = n31571 ^ n28087;
  assign n31684 = n31584 ^ n31571;
  assign n31685 = ~n31683 & ~n31684;
  assign n31686 = n31685 ^ n28087;
  assign n31699 = n31698 ^ n31686;
  assign n31701 = n31700 ^ n31699;
  assign n2573 = n2568 ^ n2499;
  assign n2577 = n2576 ^ n2573;
  assign n2578 = n2577 ^ n2553;
  assign n31702 = n31701 ^ n2578;
  assign n31587 = n31586 ^ n31568;
  assign n31588 = n31587 ^ n2467;
  assign n31589 = n31567 ^ n31542;
  assign n2448 = n2417 ^ n2389;
  assign n2458 = n2457 ^ n2448;
  assign n2459 = n2458 ^ n2440;
  assign n31590 = n31589 ^ n2459;
  assign n31592 = n29264 ^ n2336;
  assign n31593 = n31592 ^ n25775;
  assign n31594 = n31593 ^ n2455;
  assign n31591 = n31566 ^ n31565;
  assign n31595 = n31594 ^ n31591;
  assign n31596 = n31564 ^ n31543;
  assign n1402 = n1359 ^ n1299;
  assign n1403 = n1402 ^ n1396;
  assign n1407 = n1406 ^ n1403;
  assign n31597 = n31596 ^ n1407;
  assign n31598 = n31563 ^ n31562;
  assign n1384 = n1344 ^ n1281;
  assign n1385 = n1384 ^ n1381;
  assign n1389 = n1388 ^ n1385;
  assign n31599 = n31598 ^ n1389;
  assign n31600 = n31561 ^ n31560;
  assign n31601 = n31600 ^ n1374;
  assign n31602 = n31559 ^ n31558;
  assign n31606 = n31605 ^ n31602;
  assign n31607 = n31557 ^ n31556;
  assign n31611 = n31610 ^ n31607;
  assign n31612 = n31555 ^ n31554;
  assign n31613 = n31612 ^ n833;
  assign n31615 = n29282 ^ n21845;
  assign n31616 = n31615 ^ n738;
  assign n31617 = n31616 ^ n823;
  assign n31614 = n31553 ^ n31544;
  assign n31618 = n31617 ^ n31614;
  assign n31619 = n31552 ^ n31551;
  assign n740 = n720 ^ n699;
  assign n750 = n749 ^ n740;
  assign n751 = n750 ^ n733;
  assign n31620 = n31619 ^ n751;
  assign n31622 = n29289 ^ n679;
  assign n31623 = n31622 ^ n25632;
  assign n31624 = n31623 ^ n747;
  assign n31621 = n31550 ^ n31545;
  assign n31625 = n31624 ^ n31621;
  assign n31627 = n29294 ^ n670;
  assign n31628 = n31627 ^ n25738;
  assign n31629 = n31628 ^ n20600;
  assign n31626 = n31549 ^ n31546;
  assign n31630 = n31629 ^ n31626;
  assign n31194 = n31168 ^ n31151;
  assign n31198 = n31197 ^ n31194;
  assign n31199 = n31150 ^ n31131;
  assign n31203 = n31202 ^ n31199;
  assign n31281 = n31280 ^ n31204;
  assign n31282 = ~n31208 & n31281;
  assign n31283 = n31282 ^ n31207;
  assign n31284 = n31283 ^ n31199;
  assign n31285 = n31203 & ~n31284;
  assign n31286 = n31285 ^ n31202;
  assign n31287 = n31286 ^ n31194;
  assign n31288 = n31198 & ~n31287;
  assign n31289 = n31288 ^ n31197;
  assign n31189 = n31188 ^ n31169;
  assign n31631 = ~n31189 & ~n31192;
  assign n31635 = n31548 ^ n31547;
  assign n31636 = ~n31634 & ~n31635;
  assign n31637 = ~n31631 & ~n31636;
  assign n31638 = n31289 & n31637;
  assign n31639 = n31189 & n31192;
  assign n31640 = n31635 ^ n31634;
  assign n31641 = ~n31639 & n31640;
  assign n31642 = n31641 ^ n31636;
  assign n31643 = ~n31638 & n31642;
  assign n31644 = n31643 ^ n31626;
  assign n31645 = ~n31630 & ~n31644;
  assign n31646 = n31645 ^ n31629;
  assign n31647 = n31646 ^ n31621;
  assign n31648 = n31625 & ~n31647;
  assign n31649 = n31648 ^ n31624;
  assign n31650 = n31649 ^ n31619;
  assign n31651 = n31620 & ~n31650;
  assign n31652 = n31651 ^ n751;
  assign n31653 = n31652 ^ n31614;
  assign n31654 = n31618 & ~n31653;
  assign n31655 = n31654 ^ n31617;
  assign n31656 = n31655 ^ n31612;
  assign n31657 = n31613 & ~n31656;
  assign n31658 = n31657 ^ n833;
  assign n31659 = n31658 ^ n31607;
  assign n31660 = ~n31611 & n31659;
  assign n31661 = n31660 ^ n31610;
  assign n31662 = n31661 ^ n31602;
  assign n31663 = n31606 & ~n31662;
  assign n31664 = n31663 ^ n31605;
  assign n31665 = n31664 ^ n31600;
  assign n31666 = n31601 & ~n31665;
  assign n31667 = n31666 ^ n1374;
  assign n31668 = n31667 ^ n31598;
  assign n31669 = ~n31599 & n31668;
  assign n31670 = n31669 ^ n1389;
  assign n31671 = n31670 ^ n31596;
  assign n31672 = n31597 & ~n31671;
  assign n31673 = n31672 ^ n1407;
  assign n31674 = n31673 ^ n31591;
  assign n31675 = n31595 & ~n31674;
  assign n31676 = n31675 ^ n31594;
  assign n31677 = n31676 ^ n31589;
  assign n31678 = ~n31590 & n31677;
  assign n31679 = n31678 ^ n2459;
  assign n31680 = n31679 ^ n31587;
  assign n31681 = n31588 & ~n31680;
  assign n31682 = n31681 ^ n2467;
  assign n31703 = n31702 ^ n31682;
  assign n31708 = n31707 ^ n31703;
  assign n31713 = n31679 ^ n31588;
  assign n31709 = n29844 ^ n28897;
  assign n31710 = n30907 ^ n29844;
  assign n31711 = ~n31709 & n31710;
  assign n31712 = n31711 ^ n28897;
  assign n31714 = n31713 ^ n31712;
  assign n31716 = n29851 ^ n28904;
  assign n31717 = n31009 ^ n29851;
  assign n31718 = ~n31716 & ~n31717;
  assign n31719 = n31718 ^ n28904;
  assign n31715 = n31676 ^ n31590;
  assign n31720 = n31719 ^ n31715;
  assign n31725 = n31673 ^ n31595;
  assign n31721 = n30257 ^ n28912;
  assign n31722 = n31002 ^ n30257;
  assign n31723 = n31721 & n31722;
  assign n31724 = n31723 ^ n28912;
  assign n31726 = n31725 ^ n31724;
  assign n31727 = n31670 ^ n31597;
  assign n31728 = n29861 ^ n28919;
  assign n31729 = n30913 ^ n29861;
  assign n31730 = n31728 & ~n31729;
  assign n31731 = n31730 ^ n28919;
  assign n31732 = n31727 & n31731;
  assign n31733 = n31732 ^ n31725;
  assign n31734 = ~n31726 & n31733;
  assign n31735 = n31734 ^ n31732;
  assign n31736 = n31735 ^ n31715;
  assign n31737 = ~n31720 & n31736;
  assign n31738 = n31737 ^ n31719;
  assign n31739 = n31738 ^ n31713;
  assign n31740 = ~n31714 & ~n31739;
  assign n31741 = n31740 ^ n31712;
  assign n31742 = n31741 ^ n31703;
  assign n31743 = n31708 & ~n31742;
  assign n31744 = n31743 ^ n31707;
  assign n31745 = n31744 ^ n31333;
  assign n31746 = ~n31334 & n31745;
  assign n31747 = n31746 ^ n31332;
  assign n31327 = n30876 ^ n30875;
  assign n31323 = n29826 ^ n28874;
  assign n31324 = n30881 ^ n29826;
  assign n31325 = ~n31323 & ~n31324;
  assign n31326 = n31325 ^ n28874;
  assign n31328 = n31327 ^ n31326;
  assign n31784 = n31747 ^ n31328;
  assign n31785 = n31784 ^ n28914;
  assign n31786 = n31744 ^ n31334;
  assign n31787 = n31786 ^ n28989;
  assign n31788 = n31741 ^ n31708;
  assign n31789 = n31788 ^ n28999;
  assign n31790 = n31738 ^ n31714;
  assign n31791 = n31790 ^ n28922;
  assign n31792 = n31735 ^ n31720;
  assign n31793 = n31792 ^ n28853;
  assign n31794 = n31731 ^ n31727;
  assign n31795 = ~n28752 & n31794;
  assign n31796 = n31795 ^ n28771;
  assign n31797 = n31732 ^ n31724;
  assign n31798 = n31797 ^ n31725;
  assign n31799 = n31798 ^ n31795;
  assign n31800 = ~n31796 & ~n31799;
  assign n31801 = n31800 ^ n28771;
  assign n31802 = n31801 ^ n31792;
  assign n31803 = ~n31793 & ~n31802;
  assign n31804 = n31803 ^ n28853;
  assign n31805 = n31804 ^ n31790;
  assign n31806 = ~n31791 & n31805;
  assign n31807 = n31806 ^ n28922;
  assign n31808 = n31807 ^ n31788;
  assign n31809 = n31789 & n31808;
  assign n31810 = n31809 ^ n28999;
  assign n31811 = n31810 ^ n31786;
  assign n31812 = ~n31787 & n31811;
  assign n31813 = n31812 ^ n28989;
  assign n31814 = n31813 ^ n31784;
  assign n31815 = n31785 & ~n31814;
  assign n31816 = n31815 ^ n28914;
  assign n31748 = n31747 ^ n31327;
  assign n31749 = n31328 & n31748;
  assign n31750 = n31749 ^ n31326;
  assign n31318 = n30281 ^ n28867;
  assign n31319 = n31035 ^ n30281;
  assign n31320 = n31318 & n31319;
  assign n31321 = n31320 ^ n28867;
  assign n30866 = n30865 ^ n30862;
  assign n30880 = n30879 ^ n30866;
  assign n31322 = n31321 ^ n30880;
  assign n31782 = n31750 ^ n31322;
  assign n31783 = n31782 ^ n28906;
  assign n31857 = n31816 ^ n31783;
  assign n31848 = n31807 ^ n31789;
  assign n31849 = n31801 ^ n31793;
  assign n31850 = n31804 ^ n31791;
  assign n31851 = ~n31849 & n31850;
  assign n31852 = ~n31848 & n31851;
  assign n31853 = n31810 ^ n31787;
  assign n31854 = ~n31852 & n31853;
  assign n31855 = n31813 ^ n31785;
  assign n31856 = ~n31854 & n31855;
  assign n31886 = n31857 ^ n31856;
  assign n31890 = n31889 ^ n31886;
  assign n31891 = n31855 ^ n31854;
  assign n31895 = n31894 ^ n31891;
  assign n31899 = n31853 ^ n31852;
  assign n31900 = n31899 ^ n31898;
  assign n31901 = n31851 ^ n31848;
  assign n1563 = n1562 ^ n1445;
  assign n1564 = n1563 ^ n1532;
  assign n1565 = n1564 ^ n1484;
  assign n31902 = n31901 ^ n1565;
  assign n31906 = n31850 ^ n31849;
  assign n31903 = n29671 ^ n22388;
  assign n31904 = n31903 ^ n26164;
  assign n31905 = n31904 ^ n1508;
  assign n31907 = n31906 ^ n31905;
  assign n31911 = n31910 ^ n31849;
  assign n31917 = n29674 ^ n22392;
  assign n31918 = n31917 ^ n25797;
  assign n31919 = n31918 ^ n20792;
  assign n31915 = n31794 ^ n28752;
  assign n31916 = n31914 & ~n31915;
  assign n31920 = n31919 ^ n31916;
  assign n31921 = n31798 ^ n31796;
  assign n31922 = n31921 ^ n31919;
  assign n31923 = n31920 & n31922;
  assign n31924 = n31923 ^ n31916;
  assign n31925 = n31924 ^ n31849;
  assign n31926 = ~n31911 & n31925;
  assign n31927 = n31926 ^ n31910;
  assign n31928 = n31927 ^ n31906;
  assign n31929 = n31907 & ~n31928;
  assign n31930 = n31929 ^ n31905;
  assign n31931 = n31930 ^ n31901;
  assign n31932 = n31902 & ~n31931;
  assign n31933 = n31932 ^ n1565;
  assign n31934 = n31933 ^ n31899;
  assign n31935 = ~n31900 & n31934;
  assign n31936 = n31935 ^ n31898;
  assign n31937 = n31936 ^ n31891;
  assign n31938 = n31895 & ~n31937;
  assign n31939 = n31938 ^ n31894;
  assign n31940 = n31939 ^ n31886;
  assign n31941 = ~n31890 & n31940;
  assign n31942 = n31941 ^ n31889;
  assign n31882 = n29656 ^ n1872;
  assign n31883 = n31882 ^ n26137;
  assign n31884 = n31883 ^ n2032;
  assign n31817 = n31816 ^ n31782;
  assign n31818 = n31783 & n31817;
  assign n31819 = n31818 ^ n28906;
  assign n31751 = n31750 ^ n30880;
  assign n31752 = n31322 & n31751;
  assign n31753 = n31752 ^ n31321;
  assign n31313 = n30290 ^ n29591;
  assign n31314 = n31123 ^ n30290;
  assign n31315 = n31313 & n31314;
  assign n31316 = n31315 ^ n29591;
  assign n31312 = n31250 ^ n31246;
  assign n31317 = n31316 ^ n31312;
  assign n31780 = n31753 ^ n31317;
  assign n31781 = n31780 ^ n28899;
  assign n31859 = n31819 ^ n31781;
  assign n31858 = n31856 & n31857;
  assign n31881 = n31859 ^ n31858;
  assign n31885 = n31884 ^ n31881;
  assign n32877 = n31942 ^ n31885;
  assign n32921 = ~n32876 & ~n32877;
  assign n31996 = n31915 ^ n31914;
  assign n31992 = n31035 ^ n29833;
  assign n31304 = n31256 ^ n31236;
  assign n31993 = n31304 ^ n31035;
  assign n31994 = n31992 & ~n31993;
  assign n31995 = n31994 ^ n29833;
  assign n31997 = n31996 ^ n31995;
  assign n32536 = n2600 ^ n2539;
  assign n32537 = n32536 ^ n26569;
  assign n32538 = n32537 ^ n21357;
  assign n32361 = n31664 ^ n31601;
  assign n32357 = n30235 ^ n28920;
  assign n32358 = n30984 ^ n30235;
  assign n32359 = ~n32357 & ~n32358;
  assign n32360 = n32359 ^ n28920;
  assign n32362 = n32361 ^ n32360;
  assign n32009 = n31271 ^ n31220;
  assign n32005 = n29811 ^ n29788;
  assign n32006 = n31398 ^ n29788;
  assign n32007 = n32005 & ~n32006;
  assign n32008 = n32007 ^ n29811;
  assign n32010 = n32009 ^ n32008;
  assign n31968 = n29818 ^ n29795;
  assign n31969 = n31404 ^ n29795;
  assign n31970 = n31968 & n31969;
  assign n31971 = n31970 ^ n29818;
  assign n31967 = n31268 ^ n31222;
  assign n31972 = n31971 ^ n31967;
  assign n31839 = n29896 ^ n29802;
  assign n31840 = n31415 ^ n29802;
  assign n31841 = ~n31839 & n31840;
  assign n31842 = n31841 ^ n29896;
  assign n31838 = n31265 ^ n31224;
  assign n31843 = n31842 ^ n31838;
  assign n31767 = n29897 ^ n29809;
  assign n31768 = n31421 ^ n29809;
  assign n31769 = ~n31767 & ~n31768;
  assign n31770 = n31769 ^ n29897;
  assign n31766 = n31262 ^ n31226;
  assign n31771 = n31770 ^ n31766;
  assign n31298 = n31259 ^ n31231;
  assign n31294 = n30305 ^ n29828;
  assign n31295 = n31184 ^ n30305;
  assign n31296 = n31294 & n31295;
  assign n31297 = n31296 ^ n29828;
  assign n31299 = n31298 ^ n31297;
  assign n31300 = n29815 ^ n29781;
  assign n31301 = n31164 ^ n29815;
  assign n31302 = ~n31300 & n31301;
  assign n31303 = n31302 ^ n29781;
  assign n31305 = n31304 ^ n31303;
  assign n31310 = n31253 ^ n31241;
  assign n31306 = n29823 ^ n29742;
  assign n31307 = n31146 ^ n29823;
  assign n31308 = ~n31306 & n31307;
  assign n31309 = n31308 ^ n29742;
  assign n31311 = n31310 ^ n31309;
  assign n31754 = n31753 ^ n31312;
  assign n31755 = n31317 & ~n31754;
  assign n31756 = n31755 ^ n31316;
  assign n31757 = n31756 ^ n31310;
  assign n31758 = ~n31311 & n31757;
  assign n31759 = n31758 ^ n31309;
  assign n31760 = n31759 ^ n31304;
  assign n31761 = ~n31305 & n31760;
  assign n31762 = n31761 ^ n31303;
  assign n31763 = n31762 ^ n31298;
  assign n31764 = n31299 & n31763;
  assign n31765 = n31764 ^ n31297;
  assign n31835 = n31766 ^ n31765;
  assign n31836 = n31771 & ~n31835;
  assign n31837 = n31836 ^ n31770;
  assign n31964 = n31838 ^ n31837;
  assign n31965 = ~n31843 & ~n31964;
  assign n31966 = n31965 ^ n31842;
  assign n32002 = n31967 ^ n31966;
  assign n32003 = ~n31972 & ~n32002;
  assign n32004 = n32003 ^ n31971;
  assign n32040 = n32009 ^ n32004;
  assign n32041 = ~n32010 & ~n32040;
  assign n32042 = n32041 ^ n32008;
  assign n32020 = n30529 ^ n29804;
  assign n32021 = n31374 ^ n30529;
  assign n32022 = ~n32020 & ~n32021;
  assign n32023 = n32022 ^ n29804;
  assign n32084 = n32019 & n32023;
  assign n32031 = n30331 ^ n29894;
  assign n32032 = n31292 ^ n30331;
  assign n32033 = ~n32031 & n32032;
  assign n32034 = n32033 ^ n29894;
  assign n32035 = n31274 ^ n31215;
  assign n32043 = n32034 & ~n32035;
  assign n32025 = n31277 ^ n31213;
  assign n32026 = n30468 ^ n29945;
  assign n32027 = n31387 ^ n30468;
  assign n32028 = n32026 & ~n32027;
  assign n32029 = n32028 ^ n29945;
  assign n32044 = ~n32025 & n32029;
  assign n32045 = ~n32043 & ~n32044;
  assign n32059 = n31283 ^ n31203;
  assign n32060 = n30542 ^ n29797;
  assign n32061 = n31368 ^ n30542;
  assign n32062 = n32060 & n32061;
  assign n32063 = n32062 ^ n29797;
  assign n32085 = ~n32059 & ~n32063;
  assign n32086 = n32045 & ~n32085;
  assign n32087 = ~n32084 & n32086;
  assign n31193 = n31192 ^ n31189;
  assign n32105 = n31289 ^ n31189;
  assign n32106 = n31193 & ~n32105;
  assign n32107 = n32106 ^ n31192;
  assign n32108 = n32107 ^ n31640;
  assign n32109 = n30841 ^ n29972;
  assign n32110 = n31344 ^ n30841;
  assign n32111 = ~n32109 & ~n32110;
  assign n32112 = n32111 ^ n29972;
  assign n32113 = ~n32108 & n32112;
  assign n32072 = n30764 ^ n29790;
  assign n32073 = n31356 ^ n30764;
  assign n32074 = ~n32072 & n32073;
  assign n32075 = n32074 ^ n29790;
  assign n32076 = n31286 ^ n31198;
  assign n32090 = ~n32075 & ~n32076;
  assign n31290 = n31289 ^ n31193;
  assign n32093 = n30796 ^ n29868;
  assign n32094 = n31350 ^ n30796;
  assign n32095 = n32093 & ~n32094;
  assign n32096 = n32095 ^ n29868;
  assign n32101 = ~n31290 & n32096;
  assign n32125 = n30920 ^ n30047;
  assign n32126 = n31465 ^ n30920;
  assign n32127 = n32125 & n32126;
  assign n32128 = n32127 ^ n30047;
  assign n32129 = n31643 ^ n31630;
  assign n32172 = n32128 & ~n32129;
  assign n32173 = ~n32101 & ~n32172;
  assign n32174 = ~n32090 & n32173;
  assign n32175 = ~n32113 & n32174;
  assign n32176 = n32087 & n32175;
  assign n32177 = ~n32042 & n32176;
  assign n32064 = n32063 ^ n32059;
  assign n32024 = n32023 ^ n32019;
  assign n32030 = n32029 ^ n32025;
  assign n32036 = ~n32034 & n32035;
  assign n32037 = n32036 ^ n32029;
  assign n32038 = n32030 & ~n32037;
  assign n32039 = n32038 ^ n32036;
  assign n32078 = n32039 ^ n32019;
  assign n32079 = n32024 & n32078;
  assign n32080 = n32079 ^ n32023;
  assign n32081 = n32080 ^ n32063;
  assign n32082 = n32064 & n32081;
  assign n32083 = n32082 ^ n32059;
  assign n32178 = n32083 & n32175;
  assign n32130 = n32129 ^ n32128;
  assign n32077 = n32075 & n32076;
  assign n32097 = n32096 ^ n31290;
  assign n32100 = ~n32077 & ~n32097;
  assign n32102 = n32101 ^ n32100;
  assign n32114 = n32108 & ~n32112;
  assign n32115 = ~n32113 & ~n32114;
  assign n32179 = ~n32102 & n32115;
  assign n32180 = n32179 ^ n32114;
  assign n32181 = n32180 ^ n32129;
  assign n32182 = ~n32130 & n32181;
  assign n32183 = n32182 ^ n32129;
  assign n32184 = ~n32178 & ~n32183;
  assign n32185 = ~n32177 & n32184;
  assign n32205 = n31652 ^ n31618;
  assign n32206 = n30211 ^ n29423;
  assign n32207 = n31695 ^ n30211;
  assign n32208 = n32206 & n32207;
  assign n32209 = n32208 ^ n29423;
  assign n32210 = ~n32205 & n32209;
  assign n32166 = n30960 ^ n30187;
  assign n32167 = n31538 ^ n30960;
  assign n32168 = n32166 & ~n32167;
  assign n32169 = n32168 ^ n30187;
  assign n32170 = n31646 ^ n31625;
  assign n32189 = ~n32169 & ~n32170;
  assign n32192 = n30200 ^ n29433;
  assign n32193 = n31579 ^ n30200;
  assign n32194 = ~n32192 & n32193;
  assign n32195 = n32194 ^ n29433;
  assign n32196 = n31649 ^ n31620;
  assign n32201 = n32195 & ~n32196;
  assign n32219 = n30220 ^ n29421;
  assign n32220 = n30778 ^ n30220;
  assign n32221 = n32219 & ~n32220;
  assign n32222 = n32221 ^ n29421;
  assign n32223 = n31655 ^ n31613;
  assign n32246 = n32222 & ~n32223;
  assign n32247 = ~n32201 & ~n32246;
  assign n32248 = ~n32189 & n32247;
  assign n32249 = ~n32210 & n32248;
  assign n32250 = ~n32185 & n32249;
  assign n32224 = n32223 ^ n32222;
  assign n32188 = n32169 & n32170;
  assign n32197 = n32196 ^ n32195;
  assign n32200 = ~n32188 & ~n32197;
  assign n32202 = n32201 ^ n32200;
  assign n32211 = n32205 & ~n32209;
  assign n32212 = ~n32210 & ~n32211;
  assign n32251 = ~n32202 & n32212;
  assign n32252 = n32251 ^ n32211;
  assign n32253 = n32252 ^ n32222;
  assign n32254 = ~n32224 & n32253;
  assign n32255 = n32254 ^ n32223;
  assign n32256 = ~n32250 & ~n32255;
  assign n32257 = n31658 ^ n31611;
  assign n32259 = n30199 ^ n29415;
  assign n32260 = n30817 ^ n30199;
  assign n32261 = ~n32259 & ~n32260;
  assign n32262 = n32261 ^ n29415;
  assign n32348 = n32257 & ~n32262;
  assign n32270 = n30197 ^ n29470;
  assign n32271 = n30854 ^ n30197;
  assign n32272 = ~n32270 & n32271;
  assign n32273 = n32272 ^ n29470;
  assign n32274 = n31661 ^ n31606;
  assign n32349 = ~n32273 & ~n32274;
  assign n32350 = ~n32348 & ~n32349;
  assign n32351 = ~n32256 & n32350;
  assign n32275 = n32274 ^ n32273;
  assign n32352 = ~n32257 & n32262;
  assign n32353 = n32352 ^ n32274;
  assign n32354 = n32275 & ~n32353;
  assign n32355 = n32354 ^ n32273;
  assign n32356 = ~n32351 & ~n32355;
  assign n32529 = n32361 ^ n32356;
  assign n32530 = n32362 & n32529;
  assign n32531 = n32530 ^ n32360;
  assign n32527 = n31667 ^ n31599;
  assign n32523 = n30244 ^ n29482;
  assign n32524 = n30978 ^ n30244;
  assign n32525 = n32523 & ~n32524;
  assign n32526 = n32525 ^ n29482;
  assign n32528 = n32527 ^ n32526;
  assign n32532 = n32531 ^ n32528;
  assign n32533 = n32532 ^ n28737;
  assign n32363 = n32362 ^ n32356;
  assign n32364 = n32363 ^ n28703;
  assign n32011 = n32010 ^ n32004;
  assign n32012 = n32011 ^ n28949;
  assign n31973 = n31972 ^ n31966;
  assign n31974 = n31973 ^ n28956;
  assign n31844 = n31843 ^ n31837;
  assign n31845 = n31844 ^ n28962;
  assign n31772 = n31771 ^ n31765;
  assign n31773 = n31772 ^ n28870;
  assign n31774 = n31762 ^ n31299;
  assign n31775 = n31774 ^ n28876;
  assign n31776 = n31759 ^ n31305;
  assign n31777 = n31776 ^ n28885;
  assign n31778 = n31756 ^ n31311;
  assign n31779 = n31778 ^ n28891;
  assign n31820 = n31819 ^ n31780;
  assign n31821 = ~n31781 & n31820;
  assign n31822 = n31821 ^ n28899;
  assign n31823 = n31822 ^ n31778;
  assign n31824 = ~n31779 & ~n31823;
  assign n31825 = n31824 ^ n28891;
  assign n31826 = n31825 ^ n31776;
  assign n31827 = ~n31777 & n31826;
  assign n31828 = n31827 ^ n28885;
  assign n31829 = n31828 ^ n31774;
  assign n31830 = ~n31775 & ~n31829;
  assign n31831 = n31830 ^ n28876;
  assign n31832 = n31831 ^ n31772;
  assign n31833 = ~n31773 & ~n31832;
  assign n31834 = n31833 ^ n28870;
  assign n31961 = n31844 ^ n31834;
  assign n31962 = ~n31845 & ~n31961;
  assign n31963 = n31962 ^ n28962;
  assign n32013 = n31973 ^ n31963;
  assign n32014 = n31974 & ~n32013;
  assign n32015 = n32014 ^ n28956;
  assign n32016 = n32015 ^ n32011;
  assign n32017 = ~n32012 & n32016;
  assign n32018 = n32017 ^ n28949;
  assign n32046 = ~n32042 & n32045;
  assign n32047 = ~n32039 & ~n32046;
  assign n32048 = n32047 ^ n32024;
  assign n32049 = n28941 & n32048;
  assign n32050 = n32035 ^ n32034;
  assign n32051 = n32042 ^ n32035;
  assign n32052 = ~n32050 & n32051;
  assign n32053 = n32052 ^ n32034;
  assign n32054 = n32053 ^ n32030;
  assign n32055 = ~n28947 & ~n32054;
  assign n32056 = n32050 ^ n32042;
  assign n32057 = ~n29063 & ~n32056;
  assign n32058 = ~n32055 & ~n32057;
  assign n32065 = n32047 ^ n32019;
  assign n32066 = n32024 & ~n32065;
  assign n32067 = n32066 ^ n32023;
  assign n32068 = n32067 ^ n32064;
  assign n32069 = n28931 & n32068;
  assign n32070 = n32058 & ~n32069;
  assign n32071 = ~n32049 & n32070;
  assign n32088 = ~n32042 & n32087;
  assign n32089 = ~n32083 & ~n32088;
  assign n32091 = ~n32089 & ~n32090;
  assign n32092 = ~n32077 & ~n32091;
  assign n32098 = n32097 ^ n32092;
  assign n32099 = n29198 & ~n32098;
  assign n32103 = n32091 & ~n32101;
  assign n32104 = n32102 & ~n32103;
  assign n32116 = n32115 ^ n32104;
  assign n32117 = n29249 & n32116;
  assign n32118 = n32076 ^ n32075;
  assign n32119 = n32118 ^ n32089;
  assign n32120 = n29086 & n32119;
  assign n32121 = n32112 ^ n32108;
  assign n32122 = n32108 ^ n32104;
  assign n32123 = ~n32121 & n32122;
  assign n32124 = n32123 ^ n32112;
  assign n32131 = n32130 ^ n32124;
  assign n32132 = n29408 & ~n32131;
  assign n32133 = ~n32120 & ~n32132;
  assign n32134 = ~n32117 & n32133;
  assign n32135 = ~n32099 & n32134;
  assign n32136 = n32071 & n32135;
  assign n32137 = n32018 & n32136;
  assign n32138 = n32068 ^ n28931;
  assign n32139 = n32048 ^ n28941;
  assign n32140 = n32054 ^ n28947;
  assign n32141 = n29063 & n32056;
  assign n32142 = n32140 & ~n32141;
  assign n32143 = n32142 ^ n32055;
  assign n32144 = n32143 ^ n32048;
  assign n32145 = n32139 & ~n32144;
  assign n32146 = n32145 ^ n28941;
  assign n32147 = n32146 ^ n32068;
  assign n32148 = n32138 & ~n32147;
  assign n32149 = n32148 ^ n28931;
  assign n32150 = n32135 & ~n32149;
  assign n32151 = n32131 ^ n29408;
  assign n32152 = n32116 ^ n29249;
  assign n32153 = n32098 ^ n29198;
  assign n32154 = ~n29086 & ~n32119;
  assign n32155 = n32154 ^ n32098;
  assign n32156 = ~n32153 & ~n32155;
  assign n32157 = n32156 ^ n29198;
  assign n32158 = n32157 ^ n32116;
  assign n32159 = n32152 & ~n32158;
  assign n32160 = n32159 ^ n29249;
  assign n32161 = n32160 ^ n32131;
  assign n32162 = ~n32151 & ~n32161;
  assign n32163 = n32162 ^ n32131;
  assign n32164 = ~n32150 & ~n32163;
  assign n32165 = ~n32137 & n32164;
  assign n32171 = n32170 ^ n32169;
  assign n32186 = n32185 ^ n32171;
  assign n32187 = ~n29465 & n32186;
  assign n32190 = ~n32185 & ~n32189;
  assign n32191 = ~n32188 & ~n32190;
  assign n32198 = n32197 ^ n32191;
  assign n32199 = ~n28683 & ~n32198;
  assign n32203 = n32190 & ~n32201;
  assign n32204 = n32202 & ~n32203;
  assign n32213 = n32212 ^ n32204;
  assign n32214 = n28686 & n32213;
  assign n32215 = n32209 ^ n32205;
  assign n32216 = n32205 ^ n32204;
  assign n32217 = ~n32215 & n32216;
  assign n32218 = n32217 ^ n32209;
  assign n32225 = n32224 ^ n32218;
  assign n32226 = n28669 & ~n32225;
  assign n32227 = ~n32214 & ~n32226;
  assign n32228 = ~n32199 & n32227;
  assign n32229 = ~n32187 & n32228;
  assign n32230 = ~n32165 & n32229;
  assign n32231 = n32225 ^ n28669;
  assign n32232 = n32213 ^ n28686;
  assign n32233 = n32198 ^ n28683;
  assign n32234 = n29465 & ~n32186;
  assign n32235 = n32234 ^ n32198;
  assign n32236 = n32233 & ~n32235;
  assign n32237 = n32236 ^ n28683;
  assign n32238 = n32237 ^ n32213;
  assign n32239 = n32232 & n32238;
  assign n32240 = n32239 ^ n28686;
  assign n32241 = n32240 ^ n32225;
  assign n32242 = ~n32231 & n32241;
  assign n32243 = n32242 ^ n28669;
  assign n32244 = ~n32230 & n32243;
  assign n32258 = n32257 ^ n32256;
  assign n32263 = n32262 ^ n32258;
  assign n32339 = ~n28663 & ~n32263;
  assign n32267 = n32262 ^ n32257;
  assign n32268 = ~n32258 & ~n32267;
  assign n32269 = n32268 ^ n32262;
  assign n32276 = n32275 ^ n32269;
  assign n32340 = n28661 & ~n32276;
  assign n32341 = ~n32339 & ~n32340;
  assign n32342 = ~n32244 & n32341;
  assign n32277 = n32276 ^ n28661;
  assign n32343 = n28663 & n32263;
  assign n32344 = n32343 ^ n32276;
  assign n32345 = ~n32277 & ~n32344;
  assign n32346 = n32345 ^ n28661;
  assign n32347 = ~n32342 & n32346;
  assign n32520 = n32363 ^ n32347;
  assign n32521 = n32364 & ~n32520;
  assign n32522 = n32521 ^ n28703;
  assign n32534 = n32533 ^ n32522;
  assign n32365 = n32364 ^ n32347;
  assign n32245 = n32244 ^ n28663;
  assign n32264 = n32263 ^ n32244;
  assign n32265 = ~n32245 & n32264;
  assign n32266 = n32265 ^ n28663;
  assign n32278 = n32277 ^ n32266;
  assign n32279 = n32263 ^ n28663;
  assign n32280 = n32279 ^ n32244;
  assign n32512 = ~n32278 & ~n32280;
  assign n32293 = n32018 & n32071;
  assign n32294 = n32149 & ~n32293;
  assign n32295 = ~n32120 & ~n32294;
  assign n32296 = ~n32099 & n32295;
  assign n32297 = n32157 & ~n32296;
  assign n32298 = n32297 ^ n32152;
  assign n32299 = ~n32154 & ~n32295;
  assign n32300 = n32299 ^ n32153;
  assign n32301 = n32297 ^ n32116;
  assign n32302 = n32152 & ~n32301;
  assign n32303 = n32302 ^ n29249;
  assign n32304 = n32303 ^ n32151;
  assign n32305 = n32300 & n32304;
  assign n32306 = ~n32298 & n32305;
  assign n32307 = n32119 ^ n29086;
  assign n32308 = n32307 ^ n32294;
  assign n32309 = n32018 & n32058;
  assign n32310 = n32143 & ~n32309;
  assign n32311 = n32310 ^ n32048;
  assign n32312 = n32139 & ~n32311;
  assign n32313 = n32312 ^ n28941;
  assign n32314 = n32313 ^ n32138;
  assign n32315 = n32310 ^ n32139;
  assign n32316 = n32056 ^ n29063;
  assign n32317 = n32056 ^ n32018;
  assign n32318 = n32316 & ~n32317;
  assign n32319 = n32318 ^ n29063;
  assign n32320 = n32319 ^ n32140;
  assign n32321 = n32316 ^ n32018;
  assign n32322 = ~n32320 & ~n32321;
  assign n32323 = ~n32315 & ~n32322;
  assign n32324 = n32314 & ~n32323;
  assign n32325 = n32308 & n32324;
  assign n32326 = n32306 & ~n32325;
  assign n32327 = n32015 ^ n32012;
  assign n31975 = n31974 ^ n31963;
  assign n31846 = n31845 ^ n31834;
  assign n31847 = n31822 ^ n31779;
  assign n31860 = ~n31858 & ~n31859;
  assign n31861 = ~n31847 & n31860;
  assign n31862 = n31825 ^ n31777;
  assign n31863 = ~n31861 & ~n31862;
  assign n31864 = n31828 ^ n31775;
  assign n31865 = n31863 & ~n31864;
  assign n31866 = n31831 ^ n31773;
  assign n31867 = n31865 & n31866;
  assign n31976 = ~n31846 & n31867;
  assign n32328 = n31975 & ~n31976;
  assign n32329 = n32327 & ~n32328;
  assign n32330 = n32306 & ~n32315;
  assign n32331 = ~n32329 & n32330;
  assign n32281 = ~n32165 & ~n32187;
  assign n32282 = ~n32199 & n32281;
  assign n32283 = ~n32237 & ~n32282;
  assign n32288 = n32283 ^ n32232;
  assign n32284 = n32283 ^ n32213;
  assign n32285 = n32232 & ~n32284;
  assign n32286 = n32285 ^ n28686;
  assign n32287 = n32286 ^ n32231;
  assign n32289 = ~n32234 & ~n32281;
  assign n32290 = n32289 ^ n32233;
  assign n32291 = n32186 ^ n29465;
  assign n32292 = n32291 ^ n32165;
  assign n32513 = n32290 & ~n32292;
  assign n32514 = ~n32287 & n32513;
  assign n32515 = n32288 & n32514;
  assign n32516 = ~n32331 & n32515;
  assign n32517 = ~n32326 & n32516;
  assign n32518 = n32512 & ~n32517;
  assign n32519 = ~n32365 & n32518;
  assign n32535 = n32534 ^ n32519;
  assign n32539 = n32538 ^ n32535;
  assign n32367 = n30091 ^ n2523;
  assign n32368 = n32367 ^ n26480;
  assign n32369 = n32368 ^ n21328;
  assign n32332 = ~n32326 & ~n32331;
  assign n32333 = ~n32292 & n32332;
  assign n32334 = n32290 & n32333;
  assign n32335 = n32288 & n32334;
  assign n32336 = ~n32287 & n32335;
  assign n32337 = ~n32280 & ~n32336;
  assign n32338 = ~n32278 & n32337;
  assign n32366 = n32365 ^ n32338;
  assign n32370 = n32369 ^ n32366;
  assign n32371 = n32328 ^ n32327;
  assign n32375 = n32374 ^ n32371;
  assign n31977 = n31976 ^ n31975;
  assign n31981 = n31980 ^ n31977;
  assign n31868 = n31867 ^ n31846;
  assign n31872 = n31871 ^ n31868;
  assign n31873 = n31866 ^ n31865;
  assign n31874 = n31873 ^ n2215;
  assign n31875 = n31864 ^ n31863;
  assign n31876 = n31875 ^ n2200;
  assign n31877 = n31862 ^ n31861;
  assign n31878 = n31877 ^ n2054;
  assign n31879 = n31860 ^ n31847;
  assign n2025 = n1949 ^ n1890;
  assign n2035 = n2034 ^ n2025;
  assign n2039 = n2038 ^ n2035;
  assign n31880 = n31879 ^ n2039;
  assign n31943 = n31942 ^ n31881;
  assign n31944 = n31885 & ~n31943;
  assign n31945 = n31944 ^ n31884;
  assign n31946 = n31945 ^ n31879;
  assign n31947 = ~n31880 & n31946;
  assign n31948 = n31947 ^ n2039;
  assign n31949 = n31948 ^ n31877;
  assign n31950 = ~n31878 & n31949;
  assign n31951 = n31950 ^ n2054;
  assign n31952 = n31951 ^ n31875;
  assign n31953 = n31876 & ~n31952;
  assign n31954 = n31953 ^ n2200;
  assign n31955 = n31954 ^ n31873;
  assign n31956 = ~n31874 & n31955;
  assign n31957 = n31956 ^ n2215;
  assign n31958 = n31957 ^ n31868;
  assign n31959 = n31872 & ~n31958;
  assign n31960 = n31959 ^ n31871;
  assign n32376 = n31977 ^ n31960;
  assign n32377 = ~n31981 & n32376;
  assign n32378 = n32377 ^ n31980;
  assign n32379 = n32378 ^ n32371;
  assign n32380 = n32375 & ~n32379;
  assign n32381 = n32380 ^ n32374;
  assign n32382 = ~n32321 & n32329;
  assign n32383 = ~n32320 & n32382;
  assign n32384 = n32383 ^ n32315;
  assign n32385 = n29768 ^ n22363;
  assign n32386 = n32385 ^ n26243;
  assign n32387 = n32386 ^ n539;
  assign n32388 = ~n32384 & ~n32387;
  assign n32389 = n29636 ^ n22463;
  assign n32390 = n32389 ^ n26217;
  assign n32391 = n32390 ^ n621;
  assign n32392 = n32329 ^ n32321;
  assign n32393 = ~n32391 & ~n32392;
  assign n32394 = n32382 ^ n32320;
  assign n32395 = n29762 ^ n22368;
  assign n32396 = n32395 ^ n626;
  assign n32397 = n32396 ^ n21143;
  assign n32398 = ~n32394 & ~n32397;
  assign n32399 = ~n32393 & ~n32398;
  assign n32400 = ~n32315 & ~n32383;
  assign n32401 = n32400 ^ n32314;
  assign n32405 = ~n32401 & ~n32404;
  assign n32406 = n32399 & ~n32405;
  assign n32407 = ~n32388 & n32406;
  assign n921 = n882 ^ n853;
  assign n931 = n930 ^ n921;
  assign n932 = n931 ^ n914;
  assign n32408 = n32314 & ~n32400;
  assign n32409 = n32308 & n32408;
  assign n32410 = n32300 & ~n32409;
  assign n32411 = n32410 ^ n32298;
  assign n32412 = ~n932 & n32411;
  assign n32416 = n32409 ^ n32300;
  assign n32417 = ~n32415 & n32416;
  assign n32418 = n30137 ^ n788;
  assign n32419 = n32418 ^ n26505;
  assign n32420 = n32419 ^ n21215;
  assign n32421 = n32408 ^ n32308;
  assign n32422 = ~n32420 & n32421;
  assign n32423 = ~n32417 & ~n32422;
  assign n935 = n897 ^ n868;
  assign n936 = n935 ^ n919;
  assign n940 = n939 ^ n936;
  assign n32424 = ~n32298 & n32410;
  assign n32425 = n32424 ^ n32304;
  assign n32426 = ~n940 & ~n32425;
  assign n32427 = n32423 & ~n32426;
  assign n32428 = ~n32412 & n32427;
  assign n32429 = n32407 & n32428;
  assign n32430 = n32381 & n32429;
  assign n32431 = n32404 ^ n32401;
  assign n32432 = n32387 ^ n32384;
  assign n32433 = n32397 ^ n32394;
  assign n32434 = n32391 & n32392;
  assign n32435 = n32434 ^ n32394;
  assign n32436 = n32433 & ~n32435;
  assign n32437 = n32436 ^ n32397;
  assign n32438 = n32437 ^ n32384;
  assign n32439 = n32432 & ~n32438;
  assign n32440 = n32439 ^ n32387;
  assign n32441 = n32440 ^ n32401;
  assign n32442 = n32431 & ~n32441;
  assign n32443 = n32442 ^ n32404;
  assign n32444 = n32428 & n32443;
  assign n32445 = n32425 ^ n940;
  assign n32446 = n32411 ^ n932;
  assign n32447 = n32416 ^ n32415;
  assign n32448 = n32420 & ~n32421;
  assign n32449 = n32448 ^ n32416;
  assign n32450 = ~n32447 & n32449;
  assign n32451 = n32450 ^ n32415;
  assign n32452 = n32451 ^ n32411;
  assign n32453 = ~n32446 & n32452;
  assign n32454 = n32453 ^ n932;
  assign n32455 = n32454 ^ n32425;
  assign n32456 = n32445 & n32455;
  assign n32457 = n32456 ^ n32425;
  assign n32458 = ~n32444 & ~n32457;
  assign n32459 = ~n32430 & n32458;
  assign n1215 = n1214 ^ n1130;
  assign n1225 = n1224 ^ n1215;
  assign n1229 = n1228 ^ n1225;
  assign n32460 = n32334 ^ n32288;
  assign n32461 = ~n1229 & n32460;
  assign n1058 = n1038 ^ n969;
  assign n1062 = n1061 ^ n1058;
  assign n1063 = n1062 ^ n1051;
  assign n32462 = n32332 ^ n32292;
  assign n32463 = ~n1063 & ~n32462;
  assign n32464 = n30108 ^ n22354;
  assign n32465 = n32464 ^ n1056;
  assign n32466 = n32465 ^ n1219;
  assign n32467 = n32333 ^ n32290;
  assign n32468 = ~n32466 & n32467;
  assign n32469 = ~n32463 & ~n32468;
  assign n32470 = n30163 ^ n22347;
  assign n32471 = n32470 ^ n26487;
  assign n32472 = n32471 ^ n2273;
  assign n32473 = n32335 ^ n32287;
  assign n32474 = ~n32472 & ~n32473;
  assign n32475 = n32469 & ~n32474;
  assign n32476 = ~n32461 & n32475;
  assign n32477 = ~n32459 & n32476;
  assign n32478 = n32473 ^ n32472;
  assign n32479 = n32460 ^ n1229;
  assign n32480 = n32467 ^ n32466;
  assign n32481 = n1063 & n32462;
  assign n32482 = n32481 ^ n32467;
  assign n32483 = ~n32480 & n32482;
  assign n32484 = n32483 ^ n32466;
  assign n32485 = n32484 ^ n32460;
  assign n32486 = ~n32479 & n32485;
  assign n32487 = n32486 ^ n1229;
  assign n32488 = n32487 ^ n32473;
  assign n32489 = n32478 & ~n32488;
  assign n32490 = n32489 ^ n32472;
  assign n32491 = ~n32477 & ~n32490;
  assign n32492 = n30101 ^ n22528;
  assign n32493 = n32492 ^ n2282;
  assign n32494 = n32493 ^ n21278;
  assign n32495 = n32336 ^ n32280;
  assign n32496 = ~n32494 & ~n32495;
  assign n32497 = n30096 ^ n2511;
  assign n32498 = n32497 ^ n26543;
  assign n32499 = n32498 ^ n2363;
  assign n32500 = n32337 ^ n32278;
  assign n32501 = ~n32499 & n32500;
  assign n32502 = ~n32496 & ~n32501;
  assign n32503 = ~n32491 & n32502;
  assign n32504 = n32500 ^ n32499;
  assign n32505 = n32494 & n32495;
  assign n32506 = ~n32504 & ~n32505;
  assign n32507 = n32506 ^ n32501;
  assign n32508 = ~n32503 & n32507;
  assign n32509 = n32508 ^ n32366;
  assign n32510 = ~n32370 & ~n32509;
  assign n32511 = n32510 ^ n32369;
  assign n32540 = n32539 ^ n32511;
  assign n31998 = n30881 ^ n29834;
  assign n31999 = n31310 ^ n30881;
  assign n32000 = n31998 & n31999;
  assign n32001 = n32000 ^ n29834;
  assign n32541 = n32540 ^ n32001;
  assign n32546 = n32508 ^ n32370;
  assign n32542 = n30891 ^ n29844;
  assign n32543 = n31312 ^ n30891;
  assign n32544 = ~n32542 & ~n32543;
  assign n32545 = n32544 ^ n29844;
  assign n32547 = n32546 ^ n32545;
  assign n32552 = n32495 ^ n32494;
  assign n32553 = n32495 ^ n32491;
  assign n32554 = n32552 & n32553;
  assign n32555 = n32554 ^ n32494;
  assign n32556 = n32555 ^ n32504;
  assign n32548 = n30897 ^ n29851;
  assign n32549 = n30897 ^ n30880;
  assign n32550 = ~n32548 & n32549;
  assign n32551 = n32550 ^ n29851;
  assign n32557 = n32556 ^ n32551;
  assign n32562 = ~n32459 & n32469;
  assign n32563 = ~n32461 & n32562;
  assign n32564 = ~n32487 & ~n32563;
  assign n32565 = n32564 ^ n32478;
  assign n32566 = n31009 ^ n29861;
  assign n32567 = n31333 ^ n31009;
  assign n32568 = ~n32566 & n32567;
  assign n32569 = n32568 ^ n29861;
  assign n32570 = ~n32565 & n32569;
  assign n32558 = n31327 ^ n30907;
  assign n32559 = n30907 ^ n30257;
  assign n32560 = n32558 & ~n32559;
  assign n32561 = n32560 ^ n30257;
  assign n32571 = n32570 ^ n32561;
  assign n32572 = n32494 ^ n32491;
  assign n32573 = n32572 ^ n32495;
  assign n32574 = n32573 ^ n32561;
  assign n32575 = n32571 & n32574;
  assign n32576 = n32575 ^ n32570;
  assign n32577 = n32576 ^ n32556;
  assign n32578 = ~n32557 & ~n32577;
  assign n32579 = n32578 ^ n32576;
  assign n32580 = n32579 ^ n32546;
  assign n32581 = n32547 & ~n32580;
  assign n32582 = n32581 ^ n32545;
  assign n32583 = n32582 ^ n32540;
  assign n32584 = ~n32541 & ~n32583;
  assign n32585 = n32584 ^ n32001;
  assign n32586 = n32585 ^ n31996;
  assign n32587 = ~n31997 & ~n32586;
  assign n32588 = n32587 ^ n31995;
  assign n31986 = n31123 ^ n29826;
  assign n31987 = n31298 ^ n31123;
  assign n31988 = ~n31986 & ~n31987;
  assign n31989 = n31988 ^ n29826;
  assign n31990 = n31921 ^ n31920;
  assign n32652 = n31989 & n31990;
  assign n32624 = n31146 ^ n30281;
  assign n32625 = n31766 ^ n31146;
  assign n32626 = n32624 & n32625;
  assign n32627 = n32626 ^ n30281;
  assign n32628 = n31924 ^ n31911;
  assign n32653 = n32627 & n32628;
  assign n32654 = ~n32652 & ~n32653;
  assign n32655 = n32588 & n32654;
  assign n32629 = n32628 ^ n32627;
  assign n32656 = ~n31989 & ~n31990;
  assign n32657 = n32656 ^ n32627;
  assign n32658 = n32629 & n32657;
  assign n32659 = n32658 ^ n32628;
  assign n32660 = ~n32655 & n32659;
  assign n32735 = n31184 ^ n29823;
  assign n32736 = n31967 ^ n31184;
  assign n32737 = ~n32735 & ~n32736;
  assign n32738 = n32737 ^ n29823;
  assign n32739 = n31930 ^ n31902;
  assign n32893 = ~n32738 & ~n32739;
  assign n32646 = n31164 ^ n30290;
  assign n32647 = n31838 ^ n31164;
  assign n32648 = n32646 & n32647;
  assign n32649 = n32648 ^ n30290;
  assign n32650 = n31927 ^ n31907;
  assign n32894 = n32649 & ~n32650;
  assign n32895 = ~n32893 & ~n32894;
  assign n32767 = n31933 ^ n31900;
  assign n32896 = n31421 ^ n29815;
  assign n32897 = n32009 ^ n31421;
  assign n32898 = ~n32896 & n32897;
  assign n32899 = n32898 ^ n29815;
  assign n32900 = n32767 & ~n32899;
  assign n32901 = n32895 & ~n32900;
  assign n32759 = n31936 ^ n31895;
  assign n32902 = n31415 ^ n30305;
  assign n32903 = n32035 ^ n31415;
  assign n32904 = ~n32902 & n32903;
  assign n32905 = n32904 ^ n30305;
  assign n32906 = ~n32759 & ~n32905;
  assign n32907 = n32901 & ~n32906;
  assign n32752 = n31939 ^ n31890;
  assign n32879 = n31404 ^ n29809;
  assign n32880 = n32025 ^ n31404;
  assign n32881 = n32879 & n32880;
  assign n32882 = n32881 ^ n29809;
  assign n32923 = n32752 & n32882;
  assign n33029 = n32907 & ~n32923;
  assign n33030 = ~n32660 & n33029;
  assign n32909 = n32905 ^ n32759;
  assign n32910 = n32899 ^ n32767;
  assign n32740 = n32739 ^ n32738;
  assign n32911 = ~n32649 & n32650;
  assign n32912 = n32740 & ~n32911;
  assign n32913 = n32912 ^ n32893;
  assign n32914 = n32913 ^ n32767;
  assign n32915 = ~n32910 & ~n32914;
  assign n32916 = n32915 ^ n32899;
  assign n32917 = n32916 ^ n32759;
  assign n32918 = n32909 & ~n32917;
  assign n32919 = n32918 ^ n32905;
  assign n33028 = n32919 & ~n32923;
  assign n33031 = n33030 ^ n33028;
  assign n32878 = n32877 ^ n32876;
  assign n32883 = ~n32752 & ~n32882;
  assign n32884 = n32883 ^ n32876;
  assign n32885 = n32878 & ~n32884;
  assign n32886 = n32885 ^ n32877;
  assign n33032 = n33030 ^ n32886;
  assign n33033 = ~n33030 & n33032;
  assign n33034 = n33033 ^ n33030;
  assign n33035 = n33031 & ~n33034;
  assign n33036 = n33035 ^ n33033;
  assign n33037 = n33036 ^ n33030;
  assign n33038 = n33037 ^ n32886;
  assign n33039 = ~n32921 & n33038;
  assign n33040 = n33039 ^ n32886;
  assign n32871 = n31945 ^ n31880;
  assign n32867 = n31292 ^ n29795;
  assign n32868 = n32059 ^ n31292;
  assign n32869 = ~n32867 & n32868;
  assign n32870 = n32869 ^ n29795;
  assign n32872 = n32871 ^ n32870;
  assign n33046 = n33040 ^ n32872;
  assign n33047 = n33046 ^ n29818;
  assign n33048 = ~n32883 & ~n33028;
  assign n33049 = ~n33030 & n33048;
  assign n33050 = n33049 ^ n32878;
  assign n33051 = n33050 ^ n29896;
  assign n32908 = ~n32660 & n32907;
  assign n33053 = ~n32908 & ~n32919;
  assign n33052 = n32882 ^ n32752;
  assign n33054 = n33053 ^ n33052;
  assign n33055 = n33054 ^ n29897;
  assign n33056 = ~n32660 & n32901;
  assign n33057 = ~n32916 & ~n33056;
  assign n33058 = n33057 ^ n32909;
  assign n33059 = n33058 ^ n29828;
  assign n33060 = ~n32660 & n32895;
  assign n33061 = n32913 & ~n33060;
  assign n33062 = n33061 ^ n32910;
  assign n33063 = n33062 ^ n29781;
  assign n32651 = n32650 ^ n32649;
  assign n32732 = n32660 ^ n32650;
  assign n32733 = ~n32651 & n32732;
  assign n32734 = n32733 ^ n32649;
  assign n32741 = n32740 ^ n32734;
  assign n32742 = n32741 ^ n29742;
  assign n32661 = n32660 ^ n32651;
  assign n32662 = n32661 ^ n29591;
  assign n31991 = n31990 ^ n31989;
  assign n32621 = n32588 ^ n31990;
  assign n32622 = n31991 & n32621;
  assign n32623 = n32622 ^ n31989;
  assign n32630 = n32629 ^ n32623;
  assign n32631 = n32630 ^ n28867;
  assign n32589 = n32588 ^ n31991;
  assign n32590 = n32589 ^ n28874;
  assign n32591 = n32585 ^ n31997;
  assign n32592 = n32591 ^ n28882;
  assign n32593 = n32582 ^ n32541;
  assign n32594 = n32593 ^ n28895;
  assign n32595 = n32579 ^ n32547;
  assign n32596 = n32595 ^ n28897;
  assign n32597 = n32576 ^ n32557;
  assign n32598 = n32597 ^ n28904;
  assign n32599 = n32569 ^ n32565;
  assign n32600 = n28919 & ~n32599;
  assign n32601 = n32600 ^ n28912;
  assign n32602 = n32573 ^ n32571;
  assign n32603 = n32602 ^ n32600;
  assign n32604 = n32601 & n32603;
  assign n32605 = n32604 ^ n28912;
  assign n32606 = n32605 ^ n32597;
  assign n32607 = n32598 & ~n32606;
  assign n32608 = n32607 ^ n28904;
  assign n32609 = n32608 ^ n32595;
  assign n32610 = ~n32596 & ~n32609;
  assign n32611 = n32610 ^ n28897;
  assign n32612 = n32611 ^ n32593;
  assign n32613 = n32594 & ~n32612;
  assign n32614 = n32613 ^ n28895;
  assign n32615 = n32614 ^ n32591;
  assign n32616 = ~n32592 & n32615;
  assign n32617 = n32616 ^ n28882;
  assign n32618 = n32617 ^ n32589;
  assign n32619 = n32590 & n32618;
  assign n32620 = n32619 ^ n28874;
  assign n32643 = n32630 ^ n32620;
  assign n32644 = n32631 & n32643;
  assign n32645 = n32644 ^ n28867;
  assign n32729 = n32661 ^ n32645;
  assign n32730 = ~n32662 & n32729;
  assign n32731 = n32730 ^ n29591;
  assign n33064 = n32741 ^ n32731;
  assign n33065 = n32742 & ~n33064;
  assign n33066 = n33065 ^ n29742;
  assign n33067 = n33066 ^ n33062;
  assign n33068 = ~n33063 & n33067;
  assign n33069 = n33068 ^ n29781;
  assign n33070 = n33069 ^ n33058;
  assign n33071 = ~n33059 & ~n33070;
  assign n33072 = n33071 ^ n29828;
  assign n33073 = n33072 ^ n33054;
  assign n33074 = ~n33055 & n33073;
  assign n33075 = n33074 ^ n29897;
  assign n33076 = n33075 ^ n33050;
  assign n33077 = n33051 & n33076;
  assign n33078 = n33077 ^ n29896;
  assign n33079 = n33078 ^ n33046;
  assign n33080 = ~n33047 & ~n33079;
  assign n33081 = n33080 ^ n29818;
  assign n33041 = n33040 ^ n32871;
  assign n33042 = ~n32872 & n33041;
  assign n33043 = n33042 ^ n32870;
  assign n32865 = n31948 ^ n31878;
  assign n32861 = n31387 ^ n29788;
  assign n32862 = n32076 ^ n31387;
  assign n32863 = n32861 & n32862;
  assign n32864 = n32863 ^ n29788;
  assign n32866 = n32865 ^ n32864;
  assign n33044 = n33043 ^ n32866;
  assign n33045 = n33044 ^ n29811;
  assign n33132 = n33081 ^ n33045;
  assign n33133 = n33069 ^ n33059;
  assign n32632 = n32631 ^ n32620;
  assign n32633 = n32605 ^ n32598;
  assign n32634 = n32608 ^ n32596;
  assign n32635 = ~n32633 & n32634;
  assign n32636 = n32611 ^ n32594;
  assign n32637 = n32635 & n32636;
  assign n32638 = n32614 ^ n32592;
  assign n32639 = ~n32637 & n32638;
  assign n32640 = n32617 ^ n32590;
  assign n32641 = ~n32639 & n32640;
  assign n32642 = ~n32632 & n32641;
  assign n32663 = n32662 ^ n32645;
  assign n32728 = ~n32642 & n32663;
  assign n32743 = n32742 ^ n32731;
  assign n33134 = n32728 & ~n32743;
  assign n33135 = n33066 ^ n33063;
  assign n33136 = ~n33134 & ~n33135;
  assign n33137 = ~n33133 & n33136;
  assign n33138 = n33072 ^ n33055;
  assign n33139 = n33137 & n33138;
  assign n33140 = n33075 ^ n33051;
  assign n33141 = n33139 & ~n33140;
  assign n33142 = n33078 ^ n33047;
  assign n33143 = ~n33141 & n33142;
  assign n33144 = n33132 & ~n33143;
  assign n33082 = n33081 ^ n33044;
  assign n33083 = ~n33045 & ~n33082;
  assign n33084 = n33083 ^ n29811;
  assign n32941 = n31951 ^ n31876;
  assign n32937 = n31374 ^ n30331;
  assign n32938 = n31374 ^ n31290;
  assign n32939 = n32937 & ~n32938;
  assign n32940 = n32939 ^ n30331;
  assign n33020 = n32941 ^ n32940;
  assign n32887 = n32886 ^ n32870;
  assign n32888 = n32872 & n32887;
  assign n32889 = n32888 ^ n32886;
  assign n32890 = n32889 ^ n32865;
  assign n32891 = n32866 & n32890;
  assign n32892 = n32891 ^ n32864;
  assign n32920 = n32919 ^ n32908;
  assign n32922 = ~n32870 & n32871;
  assign n32924 = n32864 & n32865;
  assign n32925 = ~n32923 & ~n32924;
  assign n32926 = ~n32922 & n32925;
  assign n32927 = ~n32921 & n32926;
  assign n32928 = n32927 ^ n32908;
  assign n32929 = ~n32908 & ~n32928;
  assign n32930 = n32929 ^ n32908;
  assign n32931 = n32920 & ~n32930;
  assign n32932 = n32931 ^ n32929;
  assign n32933 = n32932 ^ n32908;
  assign n32934 = n32933 ^ n32927;
  assign n32935 = n32892 & ~n32934;
  assign n32936 = n32935 ^ n32892;
  assign n33026 = n33020 ^ n32936;
  assign n33027 = n33026 ^ n29894;
  assign n33131 = n33084 ^ n33027;
  assign n33261 = n33144 ^ n33131;
  assign n33295 = n33260 & ~n33261;
  assign n33197 = n33143 ^ n33132;
  assign n33201 = n33200 ^ n33197;
  assign n33202 = n33142 ^ n33141;
  assign n33206 = n33205 ^ n33202;
  assign n33210 = n33140 ^ n33139;
  assign n33207 = n23084 ^ n2262;
  assign n33208 = n33207 ^ n26945;
  assign n33209 = n33208 ^ n21543;
  assign n33211 = n33210 ^ n33209;
  assign n33212 = n33138 ^ n33137;
  assign n33216 = n33215 ^ n33212;
  assign n33217 = n33136 ^ n33133;
  assign n33221 = n33220 ^ n33217;
  assign n33223 = n30594 ^ n2131;
  assign n33224 = n33223 ^ n1910;
  assign n33225 = n33224 ^ n21607;
  assign n33222 = n33135 ^ n33134;
  assign n33226 = n33225 ^ n33222;
  assign n32744 = n32743 ^ n32728;
  assign n32748 = n32747 ^ n32744;
  assign n32664 = n32663 ^ n32642;
  assign n1761 = n1760 ^ n1709;
  assign n1771 = n1770 ^ n1761;
  assign n1775 = n1774 ^ n1771;
  assign n32665 = n32664 ^ n1775;
  assign n32669 = n32641 ^ n32632;
  assign n32670 = n32669 ^ n32668;
  assign n32671 = n32640 ^ n32639;
  assign n32672 = n32671 ^ n1677;
  assign n32676 = n32636 ^ n32635;
  assign n32677 = ~n32675 & n32676;
  assign n32678 = n30613 ^ n1591;
  assign n32679 = n32678 ^ n26989;
  assign n32680 = n32679 ^ n1667;
  assign n32681 = n32638 ^ n32637;
  assign n32682 = ~n32680 & n32681;
  assign n32683 = ~n32677 & ~n32682;
  assign n32684 = n32634 ^ n32633;
  assign n32688 = n32687 ^ n32684;
  assign n32692 = n32691 ^ n32633;
  assign n32698 = n30621 ^ n22537;
  assign n32699 = n32698 ^ n26967;
  assign n32700 = n32699 ^ n21568;
  assign n32693 = n32599 ^ n28919;
  assign n32694 = n23280 ^ n2570;
  assign n32695 = n32694 ^ n30976;
  assign n32696 = n32695 ^ n1550;
  assign n32697 = ~n32693 & n32696;
  assign n32701 = n32700 ^ n32697;
  assign n32702 = n32602 ^ n32601;
  assign n32703 = n32702 ^ n32700;
  assign n32704 = n32701 & n32703;
  assign n32705 = n32704 ^ n32697;
  assign n32706 = n32705 ^ n32633;
  assign n32707 = ~n32692 & n32706;
  assign n32708 = n32707 ^ n32691;
  assign n32709 = n32708 ^ n32684;
  assign n32710 = n32688 & ~n32709;
  assign n32711 = n32710 ^ n32687;
  assign n32712 = n32683 & n32711;
  assign n32713 = n32681 ^ n32680;
  assign n32714 = n32675 & ~n32676;
  assign n32715 = n32714 ^ n32681;
  assign n32716 = ~n32713 & n32715;
  assign n32717 = n32716 ^ n32680;
  assign n32718 = ~n32712 & ~n32717;
  assign n32719 = n32718 ^ n32671;
  assign n32720 = n32672 & n32719;
  assign n32721 = n32720 ^ n1677;
  assign n32722 = n32721 ^ n32669;
  assign n32723 = n32670 & ~n32722;
  assign n32724 = n32723 ^ n32668;
  assign n32725 = n32724 ^ n32664;
  assign n32726 = ~n32665 & n32725;
  assign n32727 = n32726 ^ n1775;
  assign n33227 = n32744 ^ n32727;
  assign n33228 = ~n32748 & n33227;
  assign n33229 = n33228 ^ n32747;
  assign n33230 = n33229 ^ n33222;
  assign n33231 = ~n33226 & n33230;
  assign n33232 = n33231 ^ n33225;
  assign n33233 = n33232 ^ n33217;
  assign n33234 = n33221 & ~n33233;
  assign n33235 = n33234 ^ n33220;
  assign n33236 = n33235 ^ n33212;
  assign n33237 = ~n33216 & n33236;
  assign n33238 = n33237 ^ n33215;
  assign n33239 = n33238 ^ n33210;
  assign n33240 = n33211 & ~n33239;
  assign n33241 = n33240 ^ n33209;
  assign n33242 = n33241 ^ n33202;
  assign n33243 = ~n33206 & n33242;
  assign n33244 = n33243 ^ n33205;
  assign n33245 = n33244 ^ n33197;
  assign n33246 = n33201 & ~n33245;
  assign n33247 = n33246 ^ n33200;
  assign n33262 = ~n33260 & n33261;
  assign n33806 = n33247 & ~n33262;
  assign n33939 = ~n33295 & ~n33806;
  assign n33145 = n33131 & n33144;
  assign n33085 = n33084 ^ n33026;
  assign n33086 = n33027 & ~n33085;
  assign n33087 = n33086 ^ n29894;
  assign n33021 = n32941 ^ n32936;
  assign n33022 = n33020 & n33021;
  assign n33023 = n33022 ^ n32940;
  assign n32947 = n31954 ^ n31874;
  assign n32943 = n31368 ^ n30468;
  assign n32944 = n32108 ^ n31368;
  assign n32945 = n32943 & n32944;
  assign n32946 = n32945 ^ n30468;
  assign n32951 = n32947 ^ n32946;
  assign n33024 = n33023 ^ n32951;
  assign n33025 = n33024 ^ n29945;
  assign n33130 = n33087 ^ n33025;
  assign n33256 = n33145 ^ n33130;
  assign n33296 = n33256 ^ n33255;
  assign n33940 = n33939 ^ n33296;
  assign n32832 = n32392 ^ n32391;
  assign n32833 = n32392 ^ n32381;
  assign n32834 = n32832 & ~n32833;
  assign n32835 = n32834 ^ n32391;
  assign n32836 = n32835 ^ n32433;
  assign n35243 = n33940 ^ n32836;
  assign n32766 = n31766 ^ n31035;
  assign n32768 = n32767 ^ n31766;
  assign n32769 = n32766 & n32768;
  assign n32770 = n32769 ^ n31035;
  assign n32765 = n32696 ^ n32693;
  assign n32771 = n32770 ^ n32765;
  assign n32772 = n31298 ^ n30881;
  assign n32773 = n32739 ^ n31298;
  assign n32774 = ~n32772 & ~n32773;
  assign n32775 = n32774 ^ n30881;
  assign n33367 = n30939 ^ n23223;
  assign n33368 = n33367 ^ n27232;
  assign n33369 = n33368 ^ n2568;
  assign n32780 = n32381 & n32407;
  assign n32781 = ~n32443 & ~n32780;
  assign n32782 = n32423 & ~n32781;
  assign n32783 = ~n32451 & ~n32782;
  assign n32793 = n32783 ^ n32446;
  assign n32789 = n30854 ^ n30220;
  assign n32790 = n31727 ^ n30854;
  assign n32791 = ~n32789 & ~n32790;
  assign n32792 = n32791 ^ n30220;
  assign n32794 = n32793 ^ n32792;
  assign n32800 = n30817 ^ n30211;
  assign n32801 = n32527 ^ n30817;
  assign n32802 = n32800 & ~n32801;
  assign n32803 = n32802 ^ n30211;
  assign n32795 = n32421 ^ n32420;
  assign n32796 = n32781 ^ n32421;
  assign n32797 = ~n32795 & ~n32796;
  assign n32798 = n32797 ^ n32420;
  assign n32799 = n32798 ^ n32447;
  assign n32804 = n32803 ^ n32799;
  assign n32809 = n32795 ^ n32781;
  assign n32805 = n30778 ^ n30200;
  assign n32806 = n32361 ^ n30778;
  assign n32807 = ~n32805 & n32806;
  assign n32808 = n32807 ^ n30200;
  assign n32810 = n32809 ^ n32808;
  assign n32815 = n32381 & n32399;
  assign n32816 = ~n32437 & ~n32815;
  assign n32817 = n32816 ^ n32384;
  assign n32818 = n32432 & n32817;
  assign n32819 = n32818 ^ n32387;
  assign n32820 = n32819 ^ n32431;
  assign n32811 = n31695 ^ n30960;
  assign n32812 = n32274 ^ n31695;
  assign n32813 = n32811 & ~n32812;
  assign n32814 = n32813 ^ n30960;
  assign n32821 = n32820 ^ n32814;
  assign n32826 = n32816 ^ n32432;
  assign n32822 = n31579 ^ n30920;
  assign n32823 = n32257 ^ n31579;
  assign n32824 = n32822 & ~n32823;
  assign n32825 = n32824 ^ n30920;
  assign n32827 = n32826 ^ n32825;
  assign n32828 = n31538 ^ n30841;
  assign n32829 = n32223 ^ n31538;
  assign n32830 = n32828 & ~n32829;
  assign n32831 = n32830 ^ n30841;
  assign n32837 = n32836 ^ n32831;
  assign n32842 = n32832 ^ n32381;
  assign n32838 = n31465 ^ n30796;
  assign n32839 = n32205 ^ n31465;
  assign n32840 = ~n32838 & ~n32839;
  assign n32841 = n32840 ^ n30796;
  assign n32843 = n32842 ^ n32841;
  assign n32845 = n31344 ^ n30764;
  assign n32846 = n32196 ^ n31344;
  assign n32847 = ~n32845 & ~n32846;
  assign n32848 = n32847 ^ n30764;
  assign n32844 = n32378 ^ n32375;
  assign n32849 = n32848 ^ n32844;
  assign n32850 = n31350 ^ n30542;
  assign n32851 = n32170 ^ n31350;
  assign n32852 = ~n32850 & n32851;
  assign n32853 = n32852 ^ n30542;
  assign n31982 = n31981 ^ n31960;
  assign n32854 = n32853 ^ n31982;
  assign n32859 = n31957 ^ n31872;
  assign n32855 = n31356 ^ n30529;
  assign n32856 = n32129 ^ n31356;
  assign n32857 = n32855 & ~n32856;
  assign n32858 = n32857 ^ n30529;
  assign n32860 = n32859 ^ n32858;
  assign n32942 = ~n32940 & ~n32941;
  assign n32948 = n32946 & n32947;
  assign n32949 = ~n32942 & ~n32948;
  assign n32950 = ~n32936 & n32949;
  assign n32952 = n32940 & n32941;
  assign n32953 = n32951 & ~n32952;
  assign n32954 = n32953 ^ n32948;
  assign n32955 = ~n32950 & n32954;
  assign n32956 = n32955 ^ n32859;
  assign n32957 = n32860 & n32956;
  assign n32958 = n32957 ^ n32858;
  assign n32959 = n32958 ^ n31982;
  assign n32960 = ~n32854 & n32959;
  assign n32961 = n32960 ^ n32853;
  assign n32962 = n32961 ^ n32844;
  assign n32963 = ~n32849 & ~n32962;
  assign n32964 = n32963 ^ n32848;
  assign n32965 = n32964 ^ n32842;
  assign n32966 = ~n32843 & n32965;
  assign n32967 = n32966 ^ n32841;
  assign n32968 = n32967 ^ n32836;
  assign n32969 = n32837 & n32968;
  assign n32970 = n32969 ^ n32831;
  assign n32971 = n32970 ^ n32826;
  assign n32972 = n32827 & n32971;
  assign n32973 = n32972 ^ n32825;
  assign n32974 = n32973 ^ n32820;
  assign n32975 = n32821 & n32974;
  assign n32976 = n32975 ^ n32814;
  assign n32977 = n32976 ^ n32809;
  assign n32978 = n32810 & ~n32977;
  assign n32979 = n32978 ^ n32808;
  assign n32980 = n32979 ^ n32799;
  assign n32981 = n32804 & n32980;
  assign n32982 = n32981 ^ n32803;
  assign n32983 = n32982 ^ n32793;
  assign n32984 = ~n32794 & n32983;
  assign n32985 = n32984 ^ n32792;
  assign n32784 = n32783 ^ n32411;
  assign n32785 = ~n32446 & ~n32784;
  assign n32786 = n32785 ^ n932;
  assign n32787 = n32786 ^ n32445;
  assign n32776 = n30984 ^ n30199;
  assign n32777 = n31725 ^ n30984;
  assign n32778 = n32776 & n32777;
  assign n32779 = n32778 ^ n30199;
  assign n32788 = n32787 ^ n32779;
  assign n32998 = n32985 ^ n32788;
  assign n32999 = n32998 ^ n29415;
  assign n33000 = n32982 ^ n32794;
  assign n33001 = n33000 ^ n29421;
  assign n33002 = n32979 ^ n32804;
  assign n33003 = n33002 ^ n29423;
  assign n33004 = n32976 ^ n32810;
  assign n33005 = n33004 ^ n29433;
  assign n33006 = n32973 ^ n32821;
  assign n33007 = n33006 ^ n30187;
  assign n33008 = n32970 ^ n32827;
  assign n33009 = n33008 ^ n30047;
  assign n33010 = n32967 ^ n32837;
  assign n33011 = n33010 ^ n29972;
  assign n33012 = n32964 ^ n32843;
  assign n33013 = n33012 ^ n29868;
  assign n33014 = n32961 ^ n32849;
  assign n33015 = n33014 ^ n29790;
  assign n33016 = n32958 ^ n32854;
  assign n33017 = n33016 ^ n29797;
  assign n33018 = n32955 ^ n32860;
  assign n33019 = n33018 ^ n29804;
  assign n33088 = n33087 ^ n33024;
  assign n33089 = ~n33025 & n33088;
  assign n33090 = n33089 ^ n29945;
  assign n33091 = n33090 ^ n33018;
  assign n33092 = n33019 & ~n33091;
  assign n33093 = n33092 ^ n29804;
  assign n33094 = n33093 ^ n33016;
  assign n33095 = ~n33017 & ~n33094;
  assign n33096 = n33095 ^ n29797;
  assign n33097 = n33096 ^ n33014;
  assign n33098 = ~n33015 & n33097;
  assign n33099 = n33098 ^ n29790;
  assign n33100 = n33099 ^ n33012;
  assign n33101 = ~n33013 & ~n33100;
  assign n33102 = n33101 ^ n29868;
  assign n33103 = n33102 ^ n33010;
  assign n33104 = n33011 & ~n33103;
  assign n33105 = n33104 ^ n29972;
  assign n33106 = n33105 ^ n33008;
  assign n33107 = ~n33009 & n33106;
  assign n33108 = n33107 ^ n30047;
  assign n33109 = n33108 ^ n33006;
  assign n33110 = ~n33007 & ~n33109;
  assign n33111 = n33110 ^ n30187;
  assign n33112 = n33111 ^ n33004;
  assign n33113 = ~n33005 & ~n33112;
  assign n33114 = n33113 ^ n29433;
  assign n33115 = n33114 ^ n33002;
  assign n33116 = ~n33003 & n33115;
  assign n33117 = n33116 ^ n29423;
  assign n33118 = n33117 ^ n33000;
  assign n33119 = ~n33001 & n33118;
  assign n33120 = n33119 ^ n29421;
  assign n33121 = n33120 ^ n32998;
  assign n33122 = n32999 & n33121;
  assign n33123 = n33122 ^ n29415;
  assign n32991 = n30978 ^ n30197;
  assign n32992 = n31715 ^ n30978;
  assign n32993 = ~n32991 & n32992;
  assign n32994 = n32993 ^ n30197;
  assign n32989 = n32459 ^ n1063;
  assign n32990 = n32989 ^ n32462;
  assign n32995 = n32994 ^ n32990;
  assign n32986 = n32985 ^ n32787;
  assign n32987 = ~n32788 & n32986;
  assign n32988 = n32987 ^ n32779;
  assign n32996 = n32995 ^ n32988;
  assign n32997 = n32996 ^ n29470;
  assign n33124 = n33123 ^ n32997;
  assign n33125 = n33117 ^ n33001;
  assign n33126 = n33114 ^ n33003;
  assign n33127 = n33111 ^ n33005;
  assign n33128 = n33093 ^ n33017;
  assign n33129 = n33090 ^ n33019;
  assign n33146 = ~n33130 & n33145;
  assign n33147 = ~n33129 & ~n33146;
  assign n33148 = ~n33128 & ~n33147;
  assign n33149 = n33096 ^ n33015;
  assign n33150 = n33148 & n33149;
  assign n33151 = n33099 ^ n33013;
  assign n33152 = ~n33150 & ~n33151;
  assign n33153 = n33102 ^ n33011;
  assign n33154 = n33152 & ~n33153;
  assign n33155 = n33105 ^ n33009;
  assign n33156 = n33154 & n33155;
  assign n33157 = n33108 ^ n33007;
  assign n33158 = ~n33156 & ~n33157;
  assign n33159 = n33127 & n33158;
  assign n33160 = ~n33126 & n33159;
  assign n33161 = ~n33125 & n33160;
  assign n33162 = n33120 ^ n32999;
  assign n33163 = ~n33161 & ~n33162;
  assign n33164 = ~n33124 & n33163;
  assign n33178 = n32990 ^ n32988;
  assign n33179 = n32995 & ~n33178;
  assign n33180 = n33179 ^ n32994;
  assign n33172 = n32462 ^ n1063;
  assign n33173 = n32462 ^ n32459;
  assign n33174 = n33172 & n33173;
  assign n33175 = n33174 ^ n1063;
  assign n33176 = n33175 ^ n32480;
  assign n33168 = n30913 ^ n30235;
  assign n33169 = n31713 ^ n30913;
  assign n33170 = ~n33168 & ~n33169;
  assign n33171 = n33170 ^ n30235;
  assign n33177 = n33176 ^ n33171;
  assign n33181 = n33180 ^ n33177;
  assign n33182 = n33181 ^ n28920;
  assign n33165 = n33123 ^ n32996;
  assign n33166 = ~n32997 & n33165;
  assign n33167 = n33166 ^ n29470;
  assign n33183 = n33182 ^ n33167;
  assign n33365 = n33164 & ~n33183;
  assign n33359 = ~n32484 & ~n32562;
  assign n33360 = n33359 ^ n32479;
  assign n33355 = n31002 ^ n30244;
  assign n33356 = n31703 ^ n31002;
  assign n33357 = ~n33355 & ~n33356;
  assign n33358 = n33357 ^ n30244;
  assign n33361 = n33360 ^ n33358;
  assign n33352 = n33180 ^ n33176;
  assign n33353 = n33177 & ~n33352;
  assign n33354 = n33353 ^ n33171;
  assign n33362 = n33361 ^ n33354;
  assign n33363 = n33362 ^ n29482;
  assign n33348 = n33167 ^ n28920;
  assign n33349 = n33181 ^ n33167;
  assign n33350 = n33348 & n33349;
  assign n33351 = n33350 ^ n28920;
  assign n33364 = n33363 ^ n33351;
  assign n33366 = n33365 ^ n33364;
  assign n33370 = n33369 ^ n33366;
  assign n33184 = n33183 ^ n33164;
  assign n2430 = n2429 ^ n2369;
  assign n2431 = n2430 ^ n2423;
  assign n2432 = n2431 ^ n2411;
  assign n33185 = n33184 ^ n2432;
  assign n33187 = n30805 ^ n23044;
  assign n33188 = n33187 ^ n2344;
  assign n33189 = n33188 ^ n2417;
  assign n33186 = n33163 ^ n33124;
  assign n33190 = n33189 ^ n33186;
  assign n33191 = n33162 ^ n33161;
  assign n2326 = n2315 ^ n2302;
  assign n2333 = n2332 ^ n2326;
  assign n2337 = n2336 ^ n2333;
  assign n33192 = n33191 ^ n2337;
  assign n33193 = n33160 ^ n33125;
  assign n1355 = n1336 ^ n1252;
  assign n1356 = n1355 ^ n1352;
  assign n1360 = n1359 ^ n1356;
  assign n33194 = n33193 ^ n1360;
  assign n33195 = n33159 ^ n33126;
  assign n1340 = n1324 ^ n1237;
  assign n1341 = n1340 ^ n1197;
  assign n1345 = n1344 ^ n1341;
  assign n33196 = n33195 ^ n1345;
  assign n33248 = n30712 ^ n23067;
  assign n33249 = n33248 ^ n26925;
  assign n33250 = n33249 ^ n670;
  assign n33251 = n33146 ^ n33129;
  assign n33252 = ~n33250 & ~n33251;
  assign n33257 = ~n33255 & ~n33256;
  assign n663 = n662 ^ n554;
  assign n676 = n675 ^ n663;
  assign n680 = n679 ^ n676;
  assign n33263 = n33147 ^ n33128;
  assign n33264 = ~n680 & n33263;
  assign n33265 = ~n33262 & ~n33264;
  assign n33266 = ~n33257 & n33265;
  assign n33267 = ~n33252 & n33266;
  assign n33271 = n33153 ^ n33152;
  assign n33272 = ~n33270 & n33271;
  assign n33276 = n33151 ^ n33150;
  assign n33277 = ~n33275 & ~n33276;
  assign n33278 = n30717 ^ n23062;
  assign n33279 = n33278 ^ n27055;
  assign n33280 = n33279 ^ n720;
  assign n33281 = n33149 ^ n33148;
  assign n33282 = ~n33280 & n33281;
  assign n33283 = ~n33277 & ~n33282;
  assign n33287 = n33155 ^ n33154;
  assign n33288 = ~n33286 & ~n33287;
  assign n33289 = n33283 & ~n33288;
  assign n33290 = ~n33272 & n33289;
  assign n33291 = n33267 & n33290;
  assign n33292 = n33247 & n33291;
  assign n33293 = n33263 ^ n680;
  assign n33294 = n33251 ^ n33250;
  assign n33297 = ~n33295 & n33296;
  assign n33298 = n33297 ^ n33257;
  assign n33299 = n33298 ^ n33251;
  assign n33300 = n33294 & n33299;
  assign n33301 = n33300 ^ n33250;
  assign n33302 = n33301 ^ n33263;
  assign n33303 = ~n33293 & n33302;
  assign n33304 = n33303 ^ n680;
  assign n33305 = n33290 & n33304;
  assign n33306 = n33287 ^ n33286;
  assign n33307 = n33271 ^ n33270;
  assign n33308 = n33276 ^ n33275;
  assign n33309 = n33280 & ~n33281;
  assign n33310 = n33309 ^ n33276;
  assign n33311 = n33308 & ~n33310;
  assign n33312 = n33311 ^ n33275;
  assign n33313 = n33312 ^ n33270;
  assign n33314 = ~n33307 & ~n33313;
  assign n33315 = n33314 ^ n33271;
  assign n33316 = n33315 ^ n33287;
  assign n33317 = n33306 & n33316;
  assign n33318 = n33317 ^ n33286;
  assign n33319 = ~n33305 & ~n33318;
  assign n33320 = ~n33292 & n33319;
  assign n1158 = n1089 ^ n1020;
  assign n1168 = n1167 ^ n1158;
  assign n1172 = n1171 ^ n1168;
  assign n33321 = n33157 ^ n33156;
  assign n33322 = ~n1172 & n33321;
  assign n33323 = n33158 ^ n33127;
  assign n33324 = ~n1187 & n33323;
  assign n33325 = ~n33322 & ~n33324;
  assign n33326 = ~n33320 & n33325;
  assign n33327 = n33323 ^ n1187;
  assign n33328 = n1172 & ~n33321;
  assign n33329 = n33328 ^ n33323;
  assign n33330 = ~n33327 & n33329;
  assign n33331 = n33330 ^ n1187;
  assign n33332 = ~n33326 & ~n33331;
  assign n33333 = n33332 ^ n33195;
  assign n33334 = n33196 & n33333;
  assign n33335 = n33334 ^ n1345;
  assign n33336 = n33335 ^ n33193;
  assign n33337 = n33194 & ~n33336;
  assign n33338 = n33337 ^ n1360;
  assign n33339 = n33338 ^ n33191;
  assign n33340 = n33192 & ~n33339;
  assign n33341 = n33340 ^ n2337;
  assign n33342 = n33341 ^ n33186;
  assign n33343 = ~n33190 & n33342;
  assign n33344 = n33343 ^ n33189;
  assign n33345 = n33344 ^ n33184;
  assign n33346 = ~n33185 & n33345;
  assign n33347 = n33346 ^ n2432;
  assign n33371 = n33370 ^ n33347;
  assign n33372 = ~n32775 & n33371;
  assign n33373 = n33372 ^ n32765;
  assign n33374 = n33373 ^ n32770;
  assign n33376 = n32650 ^ n31304;
  assign n33377 = n31304 ^ n30891;
  assign n33378 = ~n33376 & ~n33377;
  assign n33379 = n33378 ^ n30891;
  assign n33375 = n33344 ^ n33185;
  assign n33380 = n33379 ^ n33375;
  assign n33385 = n33341 ^ n33190;
  assign n33381 = n32628 ^ n31310;
  assign n33382 = n31310 ^ n30897;
  assign n33383 = n33381 & n33382;
  assign n33384 = n33383 ^ n30897;
  assign n33386 = n33385 ^ n33384;
  assign n33388 = n31312 ^ n30907;
  assign n33389 = n31990 ^ n31312;
  assign n33390 = n33388 & ~n33389;
  assign n33391 = n33390 ^ n30907;
  assign n33387 = n33338 ^ n33192;
  assign n33392 = n33391 ^ n33387;
  assign n33393 = n31009 ^ n30880;
  assign n33394 = n31996 ^ n30880;
  assign n33395 = n33393 & ~n33394;
  assign n33396 = n33395 ^ n31009;
  assign n33397 = n33335 ^ n33194;
  assign n33398 = ~n33396 & n33397;
  assign n33399 = n33398 ^ n33387;
  assign n33400 = n33392 & n33399;
  assign n33401 = n33400 ^ n33398;
  assign n33402 = n33401 ^ n33385;
  assign n33403 = ~n33386 & n33402;
  assign n33404 = n33403 ^ n33384;
  assign n33405 = n33404 ^ n33375;
  assign n33406 = n33380 & n33405;
  assign n33407 = n33406 ^ n33379;
  assign n33408 = n32775 & ~n33371;
  assign n33409 = ~n33407 & ~n33408;
  assign n33410 = n33409 ^ n32770;
  assign n33411 = n33410 ^ n32770;
  assign n33412 = ~n33374 & ~n33411;
  assign n33413 = n33412 ^ n32770;
  assign n33414 = ~n32771 & n33413;
  assign n33415 = n33414 ^ n32765;
  assign n32763 = n32702 ^ n32701;
  assign n32758 = n31838 ^ n31123;
  assign n32760 = n32759 ^ n31838;
  assign n32761 = n32758 & ~n32760;
  assign n32762 = n32761 ^ n31123;
  assign n32764 = n32763 ^ n32762;
  assign n33528 = n33415 ^ n32764;
  assign n33529 = n33528 ^ n29826;
  assign n33530 = n33371 ^ n32775;
  assign n33531 = n33407 ^ n33371;
  assign n33532 = ~n33530 & n33531;
  assign n33533 = n33532 ^ n32775;
  assign n33534 = n33533 ^ n32771;
  assign n33535 = n33534 ^ n29833;
  assign n33536 = n33530 ^ n33407;
  assign n33537 = n33536 ^ n29834;
  assign n33538 = n33404 ^ n33380;
  assign n33539 = n33538 ^ n29844;
  assign n33540 = n33401 ^ n33386;
  assign n33541 = n33540 ^ n29851;
  assign n33542 = n33397 ^ n33396;
  assign n33543 = n29861 & ~n33542;
  assign n33544 = n33543 ^ n30257;
  assign n33545 = n33398 ^ n33391;
  assign n33546 = n33545 ^ n33387;
  assign n33547 = n33546 ^ n33543;
  assign n33548 = n33544 & n33547;
  assign n33549 = n33548 ^ n30257;
  assign n33550 = n33549 ^ n33540;
  assign n33551 = n33541 & n33550;
  assign n33552 = n33551 ^ n29851;
  assign n33553 = n33552 ^ n33538;
  assign n33554 = n33539 & n33553;
  assign n33555 = n33554 ^ n29844;
  assign n33556 = n33555 ^ n33536;
  assign n33557 = ~n33537 & ~n33556;
  assign n33558 = n33557 ^ n29834;
  assign n33559 = n33558 ^ n33534;
  assign n33560 = n33535 & n33559;
  assign n33561 = n33560 ^ n29833;
  assign n33562 = n33561 ^ n33528;
  assign n33563 = ~n33529 & ~n33562;
  assign n33564 = n33563 ^ n29826;
  assign n33416 = n33415 ^ n32763;
  assign n33417 = ~n32764 & ~n33416;
  assign n33418 = n33417 ^ n32762;
  assign n32756 = n32705 ^ n32692;
  assign n32751 = n31967 ^ n31146;
  assign n32753 = n32752 ^ n31967;
  assign n32754 = n32751 & ~n32753;
  assign n32755 = n32754 ^ n31146;
  assign n32757 = n32756 ^ n32755;
  assign n33526 = n33418 ^ n32757;
  assign n33527 = n33526 ^ n30281;
  assign n33606 = n33564 ^ n33527;
  assign n33607 = n33561 ^ n33529;
  assign n33608 = n33549 ^ n33541;
  assign n33609 = n33552 ^ n33539;
  assign n33610 = ~n33608 & n33609;
  assign n33611 = n33555 ^ n33537;
  assign n33612 = n33610 & n33611;
  assign n33613 = n33558 ^ n33535;
  assign n33614 = ~n33612 & ~n33613;
  assign n33615 = n33607 & ~n33614;
  assign n33616 = ~n33606 & n33615;
  assign n33565 = n33564 ^ n33526;
  assign n33566 = ~n33527 & n33565;
  assign n33567 = n33566 ^ n30281;
  assign n33426 = n32708 ^ n32688;
  assign n33422 = n32009 ^ n31164;
  assign n33423 = n32877 ^ n32009;
  assign n33424 = ~n33422 & ~n33423;
  assign n33425 = n33424 ^ n31164;
  assign n33518 = n33426 ^ n33425;
  assign n33419 = n33418 ^ n32756;
  assign n33420 = n32757 & n33419;
  assign n33421 = n33420 ^ n32755;
  assign n33524 = n33518 ^ n33421;
  assign n33525 = n33524 ^ n30290;
  assign n33617 = n33567 ^ n33525;
  assign n33618 = ~n33616 & n33617;
  assign n33568 = n33567 ^ n33524;
  assign n33569 = ~n33525 & n33568;
  assign n33570 = n33569 ^ n30290;
  assign n33519 = n33426 ^ n33421;
  assign n33520 = ~n33518 & n33519;
  assign n33521 = n33520 ^ n33425;
  assign n33430 = n32035 ^ n31184;
  assign n33431 = n32871 ^ n32035;
  assign n33432 = ~n33430 & n33431;
  assign n33433 = n33432 ^ n31184;
  assign n33428 = n32676 ^ n32675;
  assign n33429 = n33428 ^ n32711;
  assign n33456 = n33433 ^ n33429;
  assign n33522 = n33521 ^ n33456;
  assign n33523 = n33522 ^ n29823;
  assign n33619 = n33570 ^ n33523;
  assign n33620 = n33618 & n33619;
  assign n33571 = n33570 ^ n33522;
  assign n33572 = ~n33523 & ~n33571;
  assign n33573 = n33572 ^ n29823;
  assign n33457 = ~n33425 & n33426;
  assign n33458 = n33457 ^ n33433;
  assign n33459 = n33456 & n33458;
  assign n33460 = n33459 ^ n33429;
  assign n33427 = n33425 & ~n33426;
  assign n33434 = n33429 & n33433;
  assign n33435 = ~n33427 & ~n33434;
  assign n33509 = ~n33421 & n33435;
  assign n33510 = n33460 & ~n33509;
  assign n33440 = n32711 ^ n32676;
  assign n33441 = ~n33428 & n33440;
  assign n33442 = n33441 ^ n32675;
  assign n33443 = n33442 ^ n32713;
  assign n33436 = n32025 ^ n31421;
  assign n33437 = n32865 ^ n32025;
  assign n33438 = ~n33436 & n33437;
  assign n33439 = n33438 ^ n31421;
  assign n33455 = n33443 ^ n33439;
  assign n33516 = n33510 ^ n33455;
  assign n33517 = n33516 ^ n29815;
  assign n33621 = n33573 ^ n33517;
  assign n33622 = ~n33620 & n33621;
  assign n33574 = n33573 ^ n33516;
  assign n33575 = ~n33517 & n33574;
  assign n33576 = n33575 ^ n29815;
  assign n33511 = n33510 ^ n33443;
  assign n33512 = n33455 & ~n33511;
  assign n33513 = n33512 ^ n33439;
  assign n33450 = n32718 ^ n32672;
  assign n33446 = n32019 ^ n31415;
  assign n33447 = n32941 ^ n32019;
  assign n33448 = n33446 & n33447;
  assign n33449 = n33448 ^ n31415;
  assign n33454 = n33450 ^ n33449;
  assign n33514 = n33513 ^ n33454;
  assign n33515 = n33514 ^ n30305;
  assign n33623 = n33576 ^ n33515;
  assign n33624 = n33622 & n33623;
  assign n33577 = n33576 ^ n33514;
  assign n33578 = ~n33515 & n33577;
  assign n33579 = n33578 ^ n30305;
  assign n33472 = n32721 ^ n32670;
  assign n33468 = n32059 ^ n31404;
  assign n33469 = n32947 ^ n32059;
  assign n33470 = ~n33468 & n33469;
  assign n33471 = n33470 ^ n31404;
  assign n33501 = n33472 ^ n33471;
  assign n33444 = n33439 & n33443;
  assign n33445 = n33435 & ~n33444;
  assign n33451 = n33449 & n33450;
  assign n33452 = n33445 & ~n33451;
  assign n33453 = ~n33421 & n33452;
  assign n33461 = n33460 ^ n33443;
  assign n33462 = n33455 & ~n33461;
  assign n33463 = n33462 ^ n33439;
  assign n33464 = n33463 ^ n33449;
  assign n33465 = n33454 & ~n33464;
  assign n33466 = n33465 ^ n33450;
  assign n33467 = ~n33453 & n33466;
  assign n33507 = n33501 ^ n33467;
  assign n33508 = n33507 ^ n29809;
  assign n33625 = n33579 ^ n33508;
  assign n33626 = n33624 & n33625;
  assign n33580 = n33579 ^ n33507;
  assign n33581 = ~n33508 & ~n33580;
  assign n33582 = n33581 ^ n29809;
  assign n33502 = n33472 ^ n33467;
  assign n33503 = ~n33501 & n33502;
  assign n33504 = n33503 ^ n33471;
  assign n33478 = n32724 ^ n32665;
  assign n33474 = n32076 ^ n31398;
  assign n33475 = n32859 ^ n32076;
  assign n33476 = ~n33474 & ~n33475;
  assign n33477 = n33476 ^ n31398;
  assign n33482 = n33478 ^ n33477;
  assign n33505 = n33504 ^ n33482;
  assign n33506 = n33505 ^ n29802;
  assign n33627 = n33582 ^ n33506;
  assign n33628 = n33626 & ~n33627;
  assign n33583 = n33582 ^ n33505;
  assign n33584 = ~n33506 & ~n33583;
  assign n33585 = n33584 ^ n29802;
  assign n33473 = n33471 & ~n33472;
  assign n33479 = n33477 & n33478;
  assign n33480 = ~n33473 & ~n33479;
  assign n33481 = ~n33467 & n33480;
  assign n33483 = ~n33471 & n33472;
  assign n33484 = n33483 ^ n33477;
  assign n33485 = n33482 & n33484;
  assign n33486 = n33485 ^ n33478;
  assign n33487 = ~n33481 & n33486;
  assign n32749 = n32748 ^ n32727;
  assign n31293 = n31292 ^ n31290;
  assign n31983 = n31982 ^ n31290;
  assign n31984 = ~n31293 & n31983;
  assign n31985 = n31984 ^ n31292;
  assign n32750 = n32749 ^ n31985;
  assign n33499 = n33487 ^ n32750;
  assign n33500 = n33499 ^ n29795;
  assign n33605 = n33585 ^ n33500;
  assign n33641 = n33628 ^ n33605;
  assign n33645 = n33644 ^ n33641;
  assign n1850 = n1834 ^ n1795;
  assign n1866 = n1865 ^ n1850;
  assign n1873 = n1872 ^ n1866;
  assign n33646 = n33617 ^ n33616;
  assign n33647 = ~n1873 & n33646;
  assign n33648 = n33619 ^ n33618;
  assign n33649 = ~n1891 & ~n33648;
  assign n33650 = ~n33647 & ~n33649;
  assign n1999 = n1995 ^ n1923;
  assign n2006 = n2005 ^ n1999;
  assign n2013 = n2012 ^ n2006;
  assign n33651 = n33621 ^ n33620;
  assign n33652 = ~n2013 & ~n33651;
  assign n33653 = n33650 & ~n33652;
  assign n33657 = n33623 ^ n33622;
  assign n33658 = ~n33656 & n33657;
  assign n33659 = n33653 & ~n33658;
  assign n33663 = n33615 ^ n33606;
  assign n33664 = n33663 ^ n33662;
  assign n33668 = n33614 ^ n33607;
  assign n33669 = n33668 ^ n33667;
  assign n33670 = n33613 ^ n33612;
  assign n33674 = n33673 ^ n33670;
  assign n33675 = n33611 ^ n33610;
  assign n33679 = n33678 ^ n33675;
  assign n33681 = n30865 ^ n23405;
  assign n33682 = n33681 ^ n1559;
  assign n33683 = n33682 ^ n22388;
  assign n33680 = n33609 ^ n33608;
  assign n33684 = n33683 ^ n33680;
  assign n33685 = n30874 ^ n23397;
  assign n33686 = n33685 ^ n27119;
  assign n33687 = n33686 ^ n1526;
  assign n33688 = n33687 ^ n33608;
  assign n33694 = n30869 ^ n2636;
  assign n33695 = n33694 ^ n1553;
  assign n33696 = n33695 ^ n22392;
  assign n33689 = n2648 ^ n2578;
  assign n33690 = n33689 ^ n28042;
  assign n33691 = n33690 ^ n2634;
  assign n33692 = n33542 ^ n29861;
  assign n33693 = n33691 & ~n33692;
  assign n33697 = n33696 ^ n33693;
  assign n33698 = n33546 ^ n33544;
  assign n33699 = n33698 ^ n33696;
  assign n33700 = n33697 & n33699;
  assign n33701 = n33700 ^ n33693;
  assign n33702 = n33701 ^ n33608;
  assign n33703 = ~n33688 & n33702;
  assign n33704 = n33703 ^ n33687;
  assign n33705 = n33704 ^ n33680;
  assign n33706 = n33684 & ~n33705;
  assign n33707 = n33706 ^ n33683;
  assign n33708 = n33707 ^ n33675;
  assign n33709 = ~n33679 & n33708;
  assign n33710 = n33709 ^ n33678;
  assign n33711 = n33710 ^ n33670;
  assign n33712 = n33674 & ~n33711;
  assign n33713 = n33712 ^ n33673;
  assign n33714 = n33713 ^ n33668;
  assign n33715 = n33669 & ~n33714;
  assign n33716 = n33715 ^ n33667;
  assign n33717 = n33716 ^ n33663;
  assign n33718 = n33664 & ~n33717;
  assign n33719 = n33718 ^ n33662;
  assign n33720 = n33659 & n33719;
  assign n33721 = n33657 ^ n33656;
  assign n33722 = n1873 & ~n33646;
  assign n33723 = n33648 ^ n1891;
  assign n33724 = ~n33722 & n33723;
  assign n33725 = n33724 ^ n33649;
  assign n33726 = n33651 ^ n2013;
  assign n33727 = n33725 & n33726;
  assign n33728 = n33727 ^ n33652;
  assign n33729 = n33728 ^ n33657;
  assign n33730 = ~n33721 & ~n33729;
  assign n33731 = n33730 ^ n33656;
  assign n33732 = ~n33720 & ~n33731;
  assign n33733 = n33625 ^ n33624;
  assign n33734 = ~n2192 & n33733;
  assign n33738 = n33627 ^ n33626;
  assign n33739 = ~n33737 & ~n33738;
  assign n33740 = ~n33734 & ~n33739;
  assign n33741 = ~n33732 & n33740;
  assign n33742 = n2192 & ~n33733;
  assign n33743 = n33738 ^ n33737;
  assign n33744 = ~n33742 & n33743;
  assign n33745 = n33744 ^ n33739;
  assign n33746 = ~n33741 & n33745;
  assign n33747 = n33746 ^ n33641;
  assign n33748 = n33645 & n33747;
  assign n33749 = n33748 ^ n33644;
  assign n33629 = ~n33605 & ~n33628;
  assign n33586 = n33585 ^ n33499;
  assign n33587 = ~n33500 & n33586;
  assign n33588 = n33587 ^ n29795;
  assign n33495 = n33229 ^ n33226;
  assign n33491 = n32108 ^ n31387;
  assign n33492 = n32844 ^ n32108;
  assign n33493 = ~n33491 & ~n33492;
  assign n33494 = n33493 ^ n31387;
  assign n33496 = n33495 ^ n33494;
  assign n33488 = n33487 ^ n32749;
  assign n33489 = n32750 & ~n33488;
  assign n33490 = n33489 ^ n31985;
  assign n33497 = n33496 ^ n33490;
  assign n33498 = n33497 ^ n29788;
  assign n33604 = n33588 ^ n33498;
  assign n33636 = n33629 ^ n33604;
  assign n33640 = n33639 ^ n33636;
  assign n33804 = n33749 ^ n33640;
  assign n35244 = n33940 ^ n33804;
  assign n35245 = ~n35243 & ~n35244;
  assign n35246 = n35245 ^ n32836;
  assign n34730 = n31884 ^ n1956;
  assign n34731 = n34730 ^ n28504;
  assign n34732 = n34731 ^ n2121;
  assign n34336 = n33704 ^ n33684;
  assign n34332 = n32865 ^ n32009;
  assign n34333 = n33478 ^ n32865;
  assign n34334 = ~n34332 & ~n34333;
  assign n34335 = n34334 ^ n32009;
  assign n34474 = n34336 ^ n34335;
  assign n33862 = n32871 ^ n31967;
  assign n33863 = n33472 ^ n32871;
  assign n33864 = n33862 & n33863;
  assign n33865 = n33864 ^ n31967;
  assign n33861 = n33701 ^ n33688;
  assign n33866 = n33865 ^ n33861;
  assign n33868 = n32877 ^ n31838;
  assign n33869 = n33450 ^ n32877;
  assign n33870 = n33868 & n33869;
  assign n33871 = n33870 ^ n31838;
  assign n33867 = n33698 ^ n33697;
  assign n33872 = n33871 ^ n33867;
  assign n33874 = n32752 ^ n31766;
  assign n33875 = n33443 ^ n32752;
  assign n33876 = ~n33874 & ~n33875;
  assign n33877 = n33876 ^ n31766;
  assign n33873 = n33692 ^ n33691;
  assign n33878 = n33877 ^ n33873;
  assign n34002 = n33320 ^ n1172;
  assign n34003 = n34002 ^ n33321;
  assign n33998 = n31703 ^ n30978;
  assign n33999 = n32556 ^ n31703;
  assign n34000 = ~n33998 & ~n33999;
  assign n34001 = n34000 ^ n30978;
  assign n34004 = n34003 ^ n34001;
  assign n33883 = n31713 ^ n30984;
  assign n33884 = n32573 ^ n31713;
  assign n33885 = ~n33883 & n33884;
  assign n33886 = n33885 ^ n30984;
  assign n33778 = n33247 & n33267;
  assign n33779 = ~n33304 & ~n33778;
  assign n33780 = n33283 & ~n33779;
  assign n33781 = ~n33312 & ~n33780;
  assign n33879 = n33781 ^ n33271;
  assign n33880 = ~n33307 & ~n33879;
  assign n33881 = n33880 ^ n33270;
  assign n33882 = n33881 ^ n33306;
  assign n33887 = n33886 ^ n33882;
  assign n33888 = n31715 ^ n30854;
  assign n33889 = n32565 ^ n31715;
  assign n33890 = ~n33888 & ~n33889;
  assign n33891 = n33890 ^ n30854;
  assign n33782 = n33781 ^ n33307;
  assign n33892 = n33891 ^ n33782;
  assign n33893 = n31725 ^ n30817;
  assign n33894 = n33360 ^ n31725;
  assign n33895 = ~n33893 & ~n33894;
  assign n33896 = n33895 ^ n30817;
  assign n33788 = n33281 ^ n33280;
  assign n33789 = n33779 ^ n33281;
  assign n33790 = ~n33788 & ~n33789;
  assign n33791 = n33790 ^ n33280;
  assign n33792 = n33791 ^ n33308;
  assign n33897 = n33896 ^ n33792;
  assign n33898 = n31727 ^ n30778;
  assign n33899 = n33176 ^ n31727;
  assign n33900 = ~n33898 & n33899;
  assign n33901 = n33900 ^ n30778;
  assign n33799 = n33788 ^ n33779;
  assign n33902 = n33901 ^ n33799;
  assign n33903 = n32527 ^ n31695;
  assign n33904 = n32990 ^ n32527;
  assign n33905 = ~n33903 & ~n33904;
  assign n33906 = n33905 ^ n31695;
  assign n33807 = ~n33257 & n33806;
  assign n33808 = n33298 & ~n33807;
  assign n33809 = n33808 ^ n33251;
  assign n33810 = n33294 & n33809;
  assign n33811 = n33810 ^ n33250;
  assign n33812 = n33811 ^ n33293;
  assign n33907 = n33906 ^ n33812;
  assign n33598 = n33495 ^ n33490;
  assign n33599 = n33496 & ~n33598;
  assign n33600 = n33599 ^ n33494;
  assign n33908 = n33238 ^ n33211;
  assign n33909 = n32196 ^ n31356;
  assign n33910 = n32826 ^ n32196;
  assign n33911 = n33909 & n33910;
  assign n33912 = n33911 ^ n31356;
  assign n33913 = ~n33908 & ~n33912;
  assign n33592 = n32129 ^ n31374;
  assign n33593 = n32842 ^ n32129;
  assign n33594 = n33592 & ~n33593;
  assign n33595 = n33594 ^ n31374;
  assign n33596 = n33232 ^ n33221;
  assign n33914 = ~n33595 & ~n33596;
  assign n33762 = n32170 ^ n31368;
  assign n33763 = n32836 ^ n32170;
  assign n33764 = ~n33762 & ~n33763;
  assign n33765 = n33764 ^ n31368;
  assign n33766 = n33235 ^ n33216;
  assign n33915 = n33765 & n33766;
  assign n33916 = ~n33914 & ~n33915;
  assign n33850 = n33241 ^ n33206;
  assign n33917 = n32205 ^ n31350;
  assign n33918 = n32820 ^ n32205;
  assign n33919 = ~n33917 & ~n33918;
  assign n33920 = n33919 ^ n31350;
  assign n33921 = n33850 & n33920;
  assign n33922 = n33916 & ~n33921;
  assign n33923 = ~n33913 & n33922;
  assign n33843 = n33244 ^ n33201;
  assign n33924 = n32223 ^ n31344;
  assign n33925 = n32809 ^ n32223;
  assign n33926 = n33924 & ~n33925;
  assign n33927 = n33926 ^ n31344;
  assign n33928 = ~n33843 & ~n33927;
  assign n33830 = n33261 ^ n33260;
  assign n33831 = n33830 ^ n33247;
  assign n33929 = n32257 ^ n31465;
  assign n33930 = n32799 ^ n32257;
  assign n33931 = ~n33929 & ~n33930;
  assign n33932 = n33931 ^ n31465;
  assign n33933 = n33831 & ~n33932;
  assign n33934 = ~n33928 & ~n33933;
  assign n33935 = n32274 ^ n31538;
  assign n33936 = n32793 ^ n32274;
  assign n33937 = n33935 & ~n33936;
  assign n33938 = n33937 ^ n31538;
  assign n33941 = ~n33938 & n33940;
  assign n33942 = n33934 & ~n33941;
  assign n33819 = n33808 ^ n33294;
  assign n33943 = n32361 ^ n31579;
  assign n33944 = n32787 ^ n32361;
  assign n33945 = ~n33943 & ~n33944;
  assign n33946 = n33945 ^ n31579;
  assign n33947 = n33819 & n33946;
  assign n33948 = n33942 & ~n33947;
  assign n33949 = n33923 & n33948;
  assign n33950 = ~n33600 & n33949;
  assign n33951 = n33946 ^ n33819;
  assign n33952 = n33920 ^ n33850;
  assign n33767 = n33766 ^ n33765;
  assign n33953 = n33595 & n33596;
  assign n33954 = n33953 ^ n33765;
  assign n33955 = n33767 & n33954;
  assign n33956 = n33955 ^ n33766;
  assign n33957 = n33908 & n33912;
  assign n33958 = ~n33913 & ~n33957;
  assign n33959 = ~n33956 & n33958;
  assign n33960 = n33959 ^ n33957;
  assign n33961 = n33960 ^ n33850;
  assign n33962 = n33952 & n33961;
  assign n33963 = n33962 ^ n33920;
  assign n33964 = n33942 & ~n33963;
  assign n33965 = n33964 ^ n33946;
  assign n33966 = n33965 ^ n33946;
  assign n33967 = n33932 ^ n33831;
  assign n33968 = n33843 & n33927;
  assign n33969 = n33968 ^ n33932;
  assign n33970 = ~n33967 & ~n33969;
  assign n33971 = n33970 ^ n33831;
  assign n33972 = n33938 & ~n33940;
  assign n33973 = ~n33941 & ~n33972;
  assign n33974 = ~n33971 & n33973;
  assign n33975 = n33974 ^ n33972;
  assign n33976 = n33975 ^ n33946;
  assign n33977 = n33976 ^ n33946;
  assign n33978 = ~n33966 & ~n33977;
  assign n33979 = n33978 ^ n33946;
  assign n33980 = n33951 & ~n33979;
  assign n33981 = n33980 ^ n33819;
  assign n33982 = ~n33950 & n33981;
  assign n33983 = n33982 ^ n33812;
  assign n33984 = ~n33907 & ~n33983;
  assign n33985 = n33984 ^ n33906;
  assign n33986 = n33985 ^ n33799;
  assign n33987 = ~n33902 & ~n33986;
  assign n33988 = n33987 ^ n33901;
  assign n33989 = n33988 ^ n33792;
  assign n33990 = ~n33897 & n33989;
  assign n33991 = n33990 ^ n33896;
  assign n33992 = n33991 ^ n33782;
  assign n33993 = n33892 & n33992;
  assign n33994 = n33993 ^ n33891;
  assign n33995 = n33994 ^ n33882;
  assign n33996 = ~n33887 & ~n33995;
  assign n33997 = n33996 ^ n33886;
  assign n34096 = n34003 ^ n33997;
  assign n34097 = n34004 & n34096;
  assign n34098 = n34097 ^ n34001;
  assign n34091 = n31333 ^ n30913;
  assign n34092 = n32546 ^ n31333;
  assign n34093 = n34091 & ~n34092;
  assign n34094 = n34093 ^ n30913;
  assign n34086 = n33321 ^ n1172;
  assign n34087 = n33321 ^ n33320;
  assign n34088 = ~n34086 & ~n34087;
  assign n34089 = n34088 ^ n1172;
  assign n34090 = n34089 ^ n33327;
  assign n34095 = n34094 ^ n34090;
  assign n34099 = n34098 ^ n34095;
  assign n34100 = n34099 ^ n30235;
  assign n34005 = n34004 ^ n33997;
  assign n34006 = n34005 ^ n30197;
  assign n34007 = n33994 ^ n33887;
  assign n34008 = n34007 ^ n30199;
  assign n34009 = n33991 ^ n33892;
  assign n34010 = n34009 ^ n30220;
  assign n34011 = n33988 ^ n33897;
  assign n34012 = n34011 ^ n30211;
  assign n34013 = n33985 ^ n33902;
  assign n34014 = n34013 ^ n30200;
  assign n34015 = n33982 ^ n33907;
  assign n34016 = n34015 ^ n30960;
  assign n34017 = n33940 ^ n33938;
  assign n34018 = ~n33600 & n33923;
  assign n34019 = n33963 & ~n34018;
  assign n34020 = n33934 & ~n34019;
  assign n34021 = n33971 & ~n34020;
  assign n34022 = n34021 ^ n33940;
  assign n34023 = ~n34017 & ~n34022;
  assign n34024 = n34023 ^ n33938;
  assign n34025 = n34024 ^ n33951;
  assign n34026 = n34025 ^ n30920;
  assign n34027 = n34021 ^ n33973;
  assign n34028 = n34027 ^ n30841;
  assign n34029 = n33927 ^ n33843;
  assign n34030 = n34019 ^ n33843;
  assign n34031 = n34029 & n34030;
  assign n34032 = n34031 ^ n33927;
  assign n34033 = n34032 ^ n33967;
  assign n34034 = n34033 ^ n30796;
  assign n34035 = n34029 ^ n34019;
  assign n34036 = n34035 ^ n30764;
  assign n34037 = n33912 ^ n33908;
  assign n34038 = ~n33600 & n33916;
  assign n34039 = n33956 & ~n34038;
  assign n34040 = n34039 ^ n33908;
  assign n34041 = n34037 & n34040;
  assign n34042 = n34041 ^ n33912;
  assign n34043 = n34042 ^ n33952;
  assign n34044 = n34043 ^ n30542;
  assign n34045 = n34039 ^ n33958;
  assign n34046 = n34045 ^ n30529;
  assign n33597 = n33596 ^ n33595;
  assign n33759 = n33600 ^ n33596;
  assign n33760 = n33597 & n33759;
  assign n33761 = n33760 ^ n33595;
  assign n33768 = n33767 ^ n33761;
  assign n33769 = n33768 ^ n30468;
  assign n33601 = n33600 ^ n33597;
  assign n33602 = n33601 ^ n30331;
  assign n33589 = n33588 ^ n33497;
  assign n33590 = n33498 & n33589;
  assign n33591 = n33590 ^ n29788;
  assign n33756 = n33601 ^ n33591;
  assign n33757 = ~n33602 & ~n33756;
  assign n33758 = n33757 ^ n30331;
  assign n34047 = n33768 ^ n33758;
  assign n34048 = ~n33769 & ~n34047;
  assign n34049 = n34048 ^ n30468;
  assign n34050 = n34049 ^ n34045;
  assign n34051 = ~n34046 & ~n34050;
  assign n34052 = n34051 ^ n30529;
  assign n34053 = n34052 ^ n34043;
  assign n34054 = n34044 & ~n34053;
  assign n34055 = n34054 ^ n30542;
  assign n34056 = n34055 ^ n34035;
  assign n34057 = n34036 & n34056;
  assign n34058 = n34057 ^ n30764;
  assign n34059 = n34058 ^ n34033;
  assign n34060 = n34034 & ~n34059;
  assign n34061 = n34060 ^ n30796;
  assign n34062 = n34061 ^ n34027;
  assign n34063 = ~n34028 & ~n34062;
  assign n34064 = n34063 ^ n30841;
  assign n34065 = n34064 ^ n34025;
  assign n34066 = ~n34026 & ~n34065;
  assign n34067 = n34066 ^ n30920;
  assign n34068 = n34067 ^ n34015;
  assign n34069 = n34016 & n34068;
  assign n34070 = n34069 ^ n30960;
  assign n34071 = n34070 ^ n34013;
  assign n34072 = ~n34014 & n34071;
  assign n34073 = n34072 ^ n30200;
  assign n34074 = n34073 ^ n34011;
  assign n34075 = ~n34012 & ~n34074;
  assign n34076 = n34075 ^ n30211;
  assign n34077 = n34076 ^ n34009;
  assign n34078 = n34010 & ~n34077;
  assign n34079 = n34078 ^ n30220;
  assign n34080 = n34079 ^ n34007;
  assign n34081 = n34008 & ~n34080;
  assign n34082 = n34081 ^ n30199;
  assign n34083 = n34082 ^ n34005;
  assign n34084 = n34006 & ~n34083;
  assign n34085 = n34084 ^ n30197;
  assign n34101 = n34100 ^ n34085;
  assign n34102 = n34082 ^ n34006;
  assign n34103 = n34079 ^ n34008;
  assign n34104 = n34076 ^ n34010;
  assign n34105 = n34070 ^ n34014;
  assign n34106 = n34067 ^ n34016;
  assign n34107 = n34064 ^ n34026;
  assign n34108 = n34061 ^ n34028;
  assign n34109 = n34055 ^ n34036;
  assign n33770 = n33769 ^ n33758;
  assign n33603 = n33602 ^ n33591;
  assign n33630 = ~n33604 & ~n33629;
  assign n33771 = ~n33603 & n33630;
  assign n34110 = n33770 & n33771;
  assign n34111 = n34049 ^ n34046;
  assign n34112 = ~n34110 & n34111;
  assign n34113 = n34052 ^ n34044;
  assign n34114 = ~n34112 & ~n34113;
  assign n34115 = ~n34109 & n34114;
  assign n34116 = n34058 ^ n34034;
  assign n34117 = ~n34115 & ~n34116;
  assign n34118 = n34108 & n34117;
  assign n34119 = ~n34107 & n34118;
  assign n34120 = n34106 & ~n34119;
  assign n34121 = n34105 & n34120;
  assign n34122 = n34073 ^ n34012;
  assign n34123 = n34121 & n34122;
  assign n34124 = n34104 & n34123;
  assign n34125 = ~n34103 & ~n34124;
  assign n34126 = ~n34102 & n34125;
  assign n34262 = ~n34101 & n34126;
  assign n34256 = n34098 ^ n34090;
  assign n34257 = ~n34095 & n34256;
  assign n34258 = n34257 ^ n34094;
  assign n34254 = n33332 ^ n33196;
  assign n34250 = n31327 ^ n31002;
  assign n34251 = n32540 ^ n31327;
  assign n34252 = ~n34250 & ~n34251;
  assign n34253 = n34252 ^ n31002;
  assign n34255 = n34254 ^ n34253;
  assign n34259 = n34258 ^ n34255;
  assign n34260 = n34259 ^ n30244;
  assign n34246 = n34085 ^ n30235;
  assign n34247 = n34099 ^ n34085;
  assign n34248 = n34246 & ~n34247;
  assign n34249 = n34248 ^ n30235;
  assign n34261 = n34260 ^ n34249;
  assign n34263 = n34262 ^ n34261;
  assign n34264 = n34263 ^ n2542;
  assign n34127 = n34126 ^ n34101;
  assign n2504 = n2497 ^ n2459;
  assign n2517 = n2516 ^ n2504;
  assign n2524 = n2523 ^ n2517;
  assign n34128 = n34127 ^ n2524;
  assign n34130 = n31594 ^ n2396;
  assign n34131 = n34130 ^ n27973;
  assign n34132 = n34131 ^ n2511;
  assign n34129 = n34125 ^ n34102;
  assign n34133 = n34132 ^ n34129;
  assign n34137 = n34124 ^ n34103;
  assign n34134 = n22528 ^ n1407;
  assign n34135 = n34134 ^ n28011;
  assign n34136 = n34135 ^ n2384;
  assign n34138 = n34137 ^ n34136;
  assign n34140 = n23810 ^ n1389;
  assign n34141 = n34140 ^ n27978;
  assign n34142 = n34141 ^ n22347;
  assign n34139 = n34123 ^ n34104;
  assign n34143 = n34142 ^ n34139;
  assign n34145 = n1374 ^ n1288;
  assign n34146 = n34145 ^ n27983;
  assign n34147 = n34146 ^ n1214;
  assign n34144 = n34122 ^ n34121;
  assign n34148 = n34147 ^ n34144;
  assign n33750 = n33749 ^ n33636;
  assign n33751 = ~n33640 & n33750;
  assign n33752 = n33751 ^ n33639;
  assign n775 = n768 ^ n751;
  assign n794 = n793 ^ n775;
  assign n801 = n800 ^ n794;
  assign n34149 = n34116 ^ n34115;
  assign n34150 = ~n801 & ~n34149;
  assign n34151 = n34114 ^ n34109;
  assign n34152 = n31624 ^ n27579;
  assign n34153 = n34152 ^ n706;
  assign n34154 = n34153 ^ n788;
  assign n34155 = ~n34151 & ~n34154;
  assign n34156 = ~n34150 & ~n34155;
  assign n34160 = n34111 ^ n34110;
  assign n34161 = ~n34159 & n34160;
  assign n33631 = n33630 ^ n33603;
  assign n33632 = n31197 ^ n23876;
  assign n33633 = n33632 ^ n27599;
  assign n33634 = n33633 ^ n22463;
  assign n34162 = ~n33631 & ~n33634;
  assign n33772 = n33771 ^ n33770;
  assign n33773 = n31192 ^ n23837;
  assign n33774 = n33773 ^ n27594;
  assign n33775 = n33774 ^ n22368;
  assign n34163 = n33772 & ~n33775;
  assign n34164 = ~n34162 & ~n34163;
  assign n34165 = n31629 ^ n27584;
  assign n34166 = n34165 ^ n22477;
  assign n34167 = n34166 ^ n694;
  assign n34168 = n34113 ^ n34112;
  assign n34169 = ~n34167 & n34168;
  assign n34170 = n34164 & ~n34169;
  assign n34171 = ~n34161 & n34170;
  assign n34172 = n31617 ^ n23821;
  assign n34173 = n34172 ^ n808;
  assign n34174 = n34173 ^ n882;
  assign n34175 = n34117 ^ n34108;
  assign n34176 = ~n34174 & ~n34175;
  assign n34177 = n34118 ^ n34107;
  assign n34178 = ~n905 & n34177;
  assign n34179 = ~n34176 & ~n34178;
  assign n34180 = n34171 & n34179;
  assign n34181 = n34156 & n34180;
  assign n34182 = n33752 & n34181;
  assign n34183 = n34177 ^ n905;
  assign n34184 = n34149 ^ n801;
  assign n34185 = n34151 & n34154;
  assign n34186 = n34185 ^ n34149;
  assign n34187 = n34184 & ~n34186;
  assign n34188 = n34187 ^ n801;
  assign n34189 = n34168 ^ n34167;
  assign n34190 = n34160 ^ n34159;
  assign n33776 = n33775 ^ n33772;
  assign n34191 = n33631 & n33634;
  assign n34192 = n34191 ^ n33772;
  assign n34193 = ~n33776 & n34192;
  assign n34194 = n34193 ^ n33775;
  assign n34195 = n34194 ^ n34159;
  assign n34196 = ~n34190 & n34195;
  assign n34197 = n34196 ^ n34159;
  assign n34198 = ~n34189 & n34197;
  assign n34199 = n34198 ^ n34189;
  assign n34200 = n34199 ^ n34169;
  assign n34201 = n34156 & n34200;
  assign n34202 = n34174 & n34175;
  assign n34203 = ~n34201 & ~n34202;
  assign n34204 = ~n34188 & n34203;
  assign n34205 = n34204 ^ n34177;
  assign n34206 = n34205 ^ n34177;
  assign n34207 = n34177 ^ n34176;
  assign n34208 = n34207 ^ n34177;
  assign n34209 = ~n34206 & ~n34208;
  assign n34210 = n34209 ^ n34177;
  assign n34211 = ~n34183 & n34210;
  assign n34212 = n34211 ^ n905;
  assign n34213 = ~n34182 & ~n34212;
  assign n34217 = n34119 ^ n34106;
  assign n34218 = ~n34216 & ~n34217;
  assign n34222 = n34120 ^ n34105;
  assign n34223 = ~n34221 & n34222;
  assign n34224 = ~n34218 & ~n34223;
  assign n34225 = ~n34213 & n34224;
  assign n34226 = n34222 ^ n34221;
  assign n34227 = n34216 & n34217;
  assign n34228 = ~n34226 & ~n34227;
  assign n34229 = n34228 ^ n34223;
  assign n34230 = ~n34225 & n34229;
  assign n34231 = n34230 ^ n34144;
  assign n34232 = ~n34148 & ~n34231;
  assign n34233 = n34232 ^ n34147;
  assign n34234 = n34233 ^ n34139;
  assign n34235 = ~n34143 & n34234;
  assign n34236 = n34235 ^ n34142;
  assign n34237 = n34236 ^ n34137;
  assign n34238 = n34138 & ~n34237;
  assign n34239 = n34238 ^ n34136;
  assign n34240 = n34239 ^ n34129;
  assign n34241 = ~n34133 & n34240;
  assign n34242 = n34241 ^ n34132;
  assign n34243 = n34242 ^ n34127;
  assign n34244 = ~n34128 & n34243;
  assign n34245 = n34244 ^ n2524;
  assign n34265 = n34264 ^ n34245;
  assign n34266 = n32759 ^ n31298;
  assign n34267 = n33429 ^ n32759;
  assign n34268 = n34266 & n34267;
  assign n34269 = n34268 ^ n31298;
  assign n34270 = n34265 & n34269;
  assign n34271 = n34270 ^ n33873;
  assign n34272 = n34271 ^ n33877;
  assign n34273 = ~n34265 & ~n34269;
  assign n34278 = n34242 ^ n34128;
  assign n34274 = n32767 ^ n31304;
  assign n34275 = n33426 ^ n32767;
  assign n34276 = ~n34274 & n34275;
  assign n34277 = n34276 ^ n31304;
  assign n34279 = n34278 ^ n34277;
  assign n34284 = n34239 ^ n34133;
  assign n34280 = n32739 ^ n31310;
  assign n34281 = n32756 ^ n32739;
  assign n34282 = n34280 & n34281;
  assign n34283 = n34282 ^ n31310;
  assign n34285 = n34284 ^ n34283;
  assign n34290 = n34236 ^ n34138;
  assign n34286 = n32650 ^ n31312;
  assign n34287 = n32763 ^ n32650;
  assign n34288 = ~n34286 & n34287;
  assign n34289 = n34288 ^ n31312;
  assign n34291 = n34290 ^ n34289;
  assign n34292 = n34233 ^ n34143;
  assign n34293 = n32628 ^ n30880;
  assign n34294 = n32765 ^ n32628;
  assign n34295 = n34293 & ~n34294;
  assign n34296 = n34295 ^ n30880;
  assign n34297 = ~n34292 & ~n34296;
  assign n34298 = n34297 ^ n34290;
  assign n34299 = n34291 & n34298;
  assign n34300 = n34299 ^ n34297;
  assign n34301 = n34300 ^ n34283;
  assign n34302 = ~n34285 & ~n34301;
  assign n34303 = n34302 ^ n34284;
  assign n34304 = n34303 ^ n34277;
  assign n34305 = ~n34279 & n34304;
  assign n34306 = n34305 ^ n34278;
  assign n34307 = ~n34273 & ~n34306;
  assign n34308 = n34307 ^ n33877;
  assign n34309 = n34308 ^ n33877;
  assign n34310 = ~n34272 & ~n34309;
  assign n34311 = n34310 ^ n33877;
  assign n34312 = ~n33878 & n34311;
  assign n34313 = n34312 ^ n33873;
  assign n34314 = n34313 ^ n33867;
  assign n34315 = ~n33872 & ~n34314;
  assign n34316 = n34315 ^ n33871;
  assign n34317 = n34316 ^ n33865;
  assign n34318 = n33866 & n34317;
  assign n34319 = n34318 ^ n33861;
  assign n34480 = n34474 ^ n34319;
  assign n34481 = n34480 ^ n31164;
  assign n34518 = n34316 ^ n33866;
  assign n34482 = n34313 ^ n33872;
  assign n34483 = n34482 ^ n31123;
  assign n34484 = n34269 ^ n34265;
  assign n34485 = ~n34306 & n34484;
  assign n34486 = n34485 ^ n34270;
  assign n34487 = n34486 ^ n33878;
  assign n34488 = n34487 ^ n31035;
  assign n34489 = n34484 ^ n34306;
  assign n34490 = n34489 ^ n30881;
  assign n34491 = n34303 ^ n34279;
  assign n34492 = n34491 ^ n30891;
  assign n34493 = n34300 ^ n34285;
  assign n34494 = n34493 ^ n30897;
  assign n34495 = n34296 ^ n34292;
  assign n34496 = ~n31009 & n34495;
  assign n34497 = n34496 ^ n30907;
  assign n34498 = n34297 ^ n34289;
  assign n34499 = n34498 ^ n34290;
  assign n34500 = n34499 ^ n34496;
  assign n34501 = ~n34497 & n34500;
  assign n34502 = n34501 ^ n30907;
  assign n34503 = n34502 ^ n34493;
  assign n34504 = ~n34494 & ~n34503;
  assign n34505 = n34504 ^ n30897;
  assign n34506 = n34505 ^ n34491;
  assign n34507 = ~n34492 & ~n34506;
  assign n34508 = n34507 ^ n30891;
  assign n34509 = n34508 ^ n34489;
  assign n34510 = n34490 & ~n34509;
  assign n34511 = n34510 ^ n30881;
  assign n34512 = n34511 ^ n34487;
  assign n34513 = ~n34488 & ~n34512;
  assign n34514 = n34513 ^ n31035;
  assign n34515 = n34514 ^ n34482;
  assign n34516 = n34483 & ~n34515;
  assign n34517 = n34516 ^ n31123;
  assign n34519 = n34518 ^ n34517;
  assign n34520 = n34518 ^ n31146;
  assign n34521 = ~n34519 & ~n34520;
  assign n34522 = n34521 ^ n31146;
  assign n34523 = n34522 ^ n34480;
  assign n34524 = n34481 & ~n34523;
  assign n34525 = n34524 ^ n31164;
  assign n34616 = n34525 ^ n31184;
  assign n34475 = n34335 ^ n34319;
  assign n34476 = n34474 & n34475;
  assign n34477 = n34476 ^ n34336;
  assign n34330 = n33707 ^ n33679;
  assign n34326 = n32941 ^ n32035;
  assign n34327 = n32941 ^ n32749;
  assign n34328 = n34326 & n34327;
  assign n34329 = n34328 ^ n32035;
  assign n34349 = n34330 ^ n34329;
  assign n34478 = n34477 ^ n34349;
  assign n34617 = n34616 ^ n34478;
  assign n34602 = n34502 ^ n34494;
  assign n34603 = n34505 ^ n34492;
  assign n34604 = ~n34602 & n34603;
  assign n34605 = n34508 ^ n30881;
  assign n34606 = n34605 ^ n34489;
  assign n34607 = n34604 & n34606;
  assign n34608 = n34511 ^ n34488;
  assign n34609 = ~n34607 & n34608;
  assign n34610 = n34514 ^ n34483;
  assign n34611 = ~n34609 & ~n34610;
  assign n34612 = n34519 ^ n31146;
  assign n34613 = n34611 & n34612;
  assign n34614 = n34522 ^ n34481;
  assign n34615 = ~n34613 & ~n34614;
  assign n34729 = n34617 ^ n34615;
  assign n34733 = n34732 ^ n34729;
  assign n34734 = n34614 ^ n34613;
  assign n34738 = n34737 ^ n34734;
  assign n34740 = n31894 ^ n24182;
  assign n34741 = n34740 ^ n1658;
  assign n34742 = n34741 ^ n23100;
  assign n34739 = n34612 ^ n34611;
  assign n34743 = n34742 ^ n34739;
  assign n34747 = n34610 ^ n34609;
  assign n34744 = n31898 ^ n24188;
  assign n34745 = n34744 ^ n28510;
  assign n34746 = n34745 ^ n1653;
  assign n34748 = n34747 ^ n34746;
  assign n34749 = n34608 ^ n34607;
  assign n1566 = n1565 ^ n1460;
  assign n1585 = n1584 ^ n1566;
  assign n1592 = n1591 ^ n1585;
  assign n34750 = n34749 ^ n1592;
  assign n34754 = n34606 ^ n34604;
  assign n34751 = n28515 ^ n24195;
  assign n34752 = n34751 ^ n31905;
  assign n34753 = n34752 ^ n1579;
  assign n34755 = n34754 ^ n34753;
  assign n34759 = n34603 ^ n34602;
  assign n34760 = n34759 ^ n34758;
  assign n34761 = n31919 ^ n24199;
  assign n34762 = n34761 ^ n28525;
  assign n34763 = n34762 ^ n23108;
  assign n34764 = n34763 ^ n34602;
  assign n34765 = n32538 ^ n2617;
  assign n34766 = n34765 ^ n28640;
  assign n34767 = n34766 ^ n23280;
  assign n34768 = n34495 ^ n31009;
  assign n34769 = n34767 & ~n34768;
  assign n34773 = n34772 ^ n34769;
  assign n34774 = n34499 ^ n34497;
  assign n34775 = n34774 ^ n34772;
  assign n34776 = n34773 & ~n34775;
  assign n34777 = n34776 ^ n34769;
  assign n34778 = n34777 ^ n34602;
  assign n34779 = ~n34764 & n34778;
  assign n34780 = n34779 ^ n34763;
  assign n34781 = n34780 ^ n34759;
  assign n34782 = n34760 & ~n34781;
  assign n34783 = n34782 ^ n34758;
  assign n34784 = n34783 ^ n34754;
  assign n34785 = ~n34755 & n34784;
  assign n34786 = n34785 ^ n34753;
  assign n34787 = n34786 ^ n34749;
  assign n34788 = ~n34750 & n34787;
  assign n34789 = n34788 ^ n1592;
  assign n34790 = n34789 ^ n34747;
  assign n34791 = ~n34748 & n34790;
  assign n34792 = n34791 ^ n34746;
  assign n34793 = n34792 ^ n34739;
  assign n34794 = ~n34743 & n34793;
  assign n34795 = n34794 ^ n34742;
  assign n34796 = n34795 ^ n34734;
  assign n34797 = n34738 & ~n34796;
  assign n34798 = n34797 ^ n34737;
  assign n34799 = n34798 ^ n34729;
  assign n34800 = ~n34733 & n34799;
  assign n34801 = n34800 ^ n34732;
  assign n34618 = n34615 & ~n34617;
  assign n34479 = n34478 ^ n31184;
  assign n34526 = n34525 ^ n34478;
  assign n34527 = n34479 & ~n34526;
  assign n34528 = n34527 ^ n31184;
  assign n34350 = n34335 & n34336;
  assign n34351 = ~n34349 & ~n34350;
  assign n34331 = ~n34329 & n34330;
  assign n34352 = n34351 ^ n34331;
  assign n34337 = ~n34335 & ~n34336;
  assign n34338 = ~n34331 & ~n34337;
  assign n34465 = ~n34319 & n34338;
  assign n34466 = n34352 & ~n34465;
  assign n34324 = n33710 ^ n33674;
  assign n34320 = n32947 ^ n32025;
  assign n34321 = n33495 ^ n32947;
  assign n34322 = ~n34320 & ~n34321;
  assign n34323 = n34322 ^ n32025;
  assign n34353 = n34324 ^ n34323;
  assign n34472 = n34466 ^ n34353;
  assign n34473 = n34472 ^ n31421;
  assign n34601 = n34528 ^ n34473;
  assign n34727 = n34618 ^ n34601;
  assign n2115 = n2039 ^ n1974;
  assign n2125 = n2124 ^ n2115;
  assign n2132 = n2131 ^ n2125;
  assign n34728 = n34727 ^ n2132;
  assign n35113 = n34801 ^ n34728;
  assign n35247 = n35246 ^ n35113;
  assign n35248 = n33831 ^ n32842;
  assign n33817 = n33746 ^ n33645;
  assign n35249 = n33831 ^ n33817;
  assign n35250 = ~n35248 & ~n35249;
  assign n35251 = n35250 ^ n32842;
  assign n35121 = n34798 ^ n34732;
  assign n35122 = n35121 ^ n34729;
  assign n35252 = n35251 ^ n35122;
  assign n35253 = n33843 ^ n32844;
  assign n33824 = n33733 ^ n2192;
  assign n33825 = n33733 ^ n33732;
  assign n33826 = ~n33824 & ~n33825;
  assign n33827 = n33826 ^ n2192;
  assign n33828 = n33827 ^ n33743;
  assign n35254 = n33843 ^ n33828;
  assign n35255 = n35253 & ~n35254;
  assign n35256 = n35255 ^ n32844;
  assign n35128 = n34795 ^ n34738;
  assign n35257 = n35256 ^ n35128;
  assign n35258 = n33850 ^ n31982;
  assign n34387 = n33732 ^ n2192;
  assign n34388 = n34387 ^ n33733;
  assign n35259 = n34388 ^ n33850;
  assign n35260 = n35258 & n35259;
  assign n35261 = n35260 ^ n31982;
  assign n35136 = n34792 ^ n34742;
  assign n35137 = n35136 ^ n34739;
  assign n35262 = n35261 ^ n35137;
  assign n35267 = n34789 ^ n34748;
  assign n35263 = n33908 ^ n32859;
  assign n33836 = n33650 & n33719;
  assign n33837 = n33725 & ~n33836;
  assign n33838 = n33837 ^ n33651;
  assign n33839 = n33726 & n33838;
  assign n33840 = n33839 ^ n2013;
  assign n33841 = n33840 ^ n33721;
  assign n35264 = n33908 ^ n33841;
  assign n35265 = n35263 & n35264;
  assign n35266 = n35265 ^ n32859;
  assign n35268 = n35267 ^ n35266;
  assign n35269 = n33766 ^ n32947;
  assign n33848 = n33837 ^ n33726;
  assign n35270 = n33848 ^ n33766;
  assign n35271 = n35269 & ~n35270;
  assign n35272 = n35271 ^ n32947;
  assign n35144 = n34786 ^ n1592;
  assign n35145 = n35144 ^ n34749;
  assign n35273 = n35272 ^ n35145;
  assign n35278 = n34780 ^ n34758;
  assign n35279 = n35278 ^ n34759;
  assign n35274 = n33495 ^ n32865;
  assign n33855 = n33646 ^ n1873;
  assign n34365 = n33855 ^ n33719;
  assign n35275 = n34365 ^ n33495;
  assign n35276 = n35274 & ~n35275;
  assign n35277 = n35276 ^ n32865;
  assign n35280 = n35279 ^ n35277;
  assign n35282 = n32871 ^ n32749;
  assign n34359 = n33716 ^ n33664;
  assign n35283 = n34359 ^ n32749;
  assign n35284 = n35282 & n35283;
  assign n35285 = n35284 ^ n32871;
  assign n35281 = n34777 ^ n34764;
  assign n35286 = n35285 ^ n35281;
  assign n35288 = n33478 ^ n32877;
  assign n34343 = n33713 ^ n33669;
  assign n35289 = n34343 ^ n33478;
  assign n35290 = ~n35288 & n35289;
  assign n35291 = n35290 ^ n32877;
  assign n35287 = n34774 ^ n34773;
  assign n35292 = n35291 ^ n35287;
  assign n35104 = n34768 ^ n34767;
  assign n35099 = n33472 ^ n32752;
  assign n35100 = n34324 ^ n33472;
  assign n35101 = ~n35099 & ~n35100;
  assign n35102 = n35101 ^ n32752;
  assign n35293 = n35104 ^ n35102;
  assign n34993 = n34217 ^ n34216;
  assign n34994 = n34217 ^ n34213;
  assign n34995 = n34993 & n34994;
  assign n34996 = n34995 ^ n34216;
  assign n34997 = n34996 ^ n34226;
  assign n34988 = n31996 ^ n31333;
  assign n34989 = n33375 ^ n31996;
  assign n34990 = ~n34988 & ~n34989;
  assign n34991 = n34990 ^ n31333;
  assign n34954 = n34216 ^ n34213;
  assign n34955 = n34954 ^ n34217;
  assign n34949 = n32540 ^ n31703;
  assign n34950 = n33385 ^ n32540;
  assign n34951 = ~n34949 & n34950;
  assign n34952 = n34951 ^ n31703;
  assign n34984 = n34955 ^ n34952;
  assign n34871 = n34175 ^ n34174;
  assign n34583 = n33752 & n34171;
  assign n34584 = ~n34200 & ~n34583;
  assign n34869 = n34156 & ~n34584;
  assign n34870 = ~n34188 & ~n34869;
  assign n34902 = n34870 ^ n34175;
  assign n34903 = n34871 & n34902;
  assign n34904 = n34903 ^ n34174;
  assign n34905 = n34904 ^ n34183;
  assign n34897 = n32546 ^ n31713;
  assign n34898 = n33387 ^ n32546;
  assign n34899 = n34897 & ~n34898;
  assign n34900 = n34899 ^ n31713;
  assign n34945 = n34905 ^ n34900;
  assign n34872 = n34871 ^ n34870;
  assign n34865 = n32556 ^ n31715;
  assign n34866 = n33397 ^ n32556;
  assign n34867 = n34865 & n34866;
  assign n34868 = n34867 ^ n31715;
  assign n34873 = n34872 ^ n34868;
  assign n34582 = n34154 ^ n34151;
  assign n34656 = n34584 ^ n34151;
  assign n34657 = n34582 & n34656;
  assign n34658 = n34657 ^ n34154;
  assign n34659 = n34658 ^ n34184;
  assign n34652 = n32573 ^ n31725;
  assign n34653 = n34254 ^ n32573;
  assign n34654 = ~n34652 & ~n34653;
  assign n34655 = n34654 ^ n31725;
  assign n34660 = n34659 ^ n34655;
  assign n34585 = n34584 ^ n34582;
  assign n34578 = n32565 ^ n31727;
  assign n34579 = n34090 ^ n32565;
  assign n34580 = ~n34578 & ~n34579;
  assign n34581 = n34580 ^ n31727;
  assign n34586 = n34585 ^ n34581;
  assign n34412 = n33752 & n34164;
  assign n34413 = ~n34194 & ~n34412;
  assign n34427 = n34413 ^ n34160;
  assign n34428 = ~n34190 & ~n34427;
  assign n34429 = n34428 ^ n34159;
  assign n34430 = n34429 ^ n34189;
  assign n34423 = n33360 ^ n32527;
  assign n34424 = n34003 ^ n33360;
  assign n34425 = ~n34423 & ~n34424;
  assign n34426 = n34425 ^ n32527;
  assign n34431 = n34430 ^ n34426;
  assign n34414 = n34413 ^ n34190;
  assign n33783 = n33782 ^ n32990;
  assign n33784 = n32990 ^ n32274;
  assign n33785 = n33783 & ~n33784;
  assign n33786 = n33785 ^ n32274;
  assign n33635 = n33634 ^ n33631;
  assign n33753 = n33752 ^ n33631;
  assign n33754 = n33635 & ~n33753;
  assign n33755 = n33754 ^ n33634;
  assign n33777 = n33776 ^ n33755;
  assign n33787 = n33786 ^ n33777;
  assign n33797 = n33752 ^ n33635;
  assign n33793 = n33792 ^ n32787;
  assign n33794 = n32787 ^ n32257;
  assign n33795 = ~n33793 & ~n33794;
  assign n33796 = n33795 ^ n32257;
  assign n33798 = n33797 ^ n33796;
  assign n33800 = n33799 ^ n32793;
  assign n33801 = n32793 ^ n32223;
  assign n33802 = ~n33800 & n33801;
  assign n33803 = n33802 ^ n32223;
  assign n33805 = n33804 ^ n33803;
  assign n33813 = n33812 ^ n32799;
  assign n33814 = n32799 ^ n32205;
  assign n33815 = ~n33813 & ~n33814;
  assign n33816 = n33815 ^ n32205;
  assign n33818 = n33817 ^ n33816;
  assign n33820 = n33819 ^ n32809;
  assign n33821 = n32809 ^ n32196;
  assign n33822 = n33820 & n33821;
  assign n33823 = n33822 ^ n32196;
  assign n33829 = n33828 ^ n33823;
  assign n33832 = n33831 ^ n32826;
  assign n33833 = n32826 ^ n32129;
  assign n33834 = ~n33832 & ~n33833;
  assign n33835 = n33834 ^ n32129;
  assign n33842 = n33841 ^ n33835;
  assign n33844 = n33843 ^ n32836;
  assign n33845 = n32836 ^ n32108;
  assign n33846 = ~n33844 & n33845;
  assign n33847 = n33846 ^ n32108;
  assign n33849 = n33848 ^ n33847;
  assign n33856 = n33719 ^ n33646;
  assign n33857 = ~n33855 & n33856;
  assign n33858 = n33857 ^ n1873;
  assign n33859 = n33858 ^ n33723;
  assign n33851 = n33850 ^ n32842;
  assign n33852 = n32842 ^ n31290;
  assign n33853 = n33851 & n33852;
  assign n33854 = n33853 ^ n31290;
  assign n33860 = n33859 ^ n33854;
  assign n34325 = ~n34323 & ~n34324;
  assign n34339 = n32859 ^ n32019;
  assign n34340 = n33596 ^ n32859;
  assign n34341 = ~n34339 & ~n34340;
  assign n34342 = n34341 ^ n32019;
  assign n34344 = n34342 & ~n34343;
  assign n34345 = n34338 & ~n34344;
  assign n34346 = ~n34325 & n34345;
  assign n34347 = ~n34319 & n34346;
  assign n34348 = n34343 ^ n34342;
  assign n34354 = n34352 & n34353;
  assign n34355 = n34354 ^ n34325;
  assign n34356 = ~n34348 & n34355;
  assign n34357 = n34356 ^ n34344;
  assign n34358 = ~n34347 & n34357;
  assign n34360 = n33766 ^ n31982;
  assign n34361 = n32059 ^ n31982;
  assign n34362 = ~n34360 & ~n34361;
  assign n34363 = n34362 ^ n32059;
  assign n34364 = ~n34359 & ~n34363;
  assign n34366 = n32844 ^ n32076;
  assign n34367 = n33908 ^ n32844;
  assign n34368 = n34366 & ~n34367;
  assign n34369 = n34368 ^ n32076;
  assign n34370 = n34365 & ~n34369;
  assign n34371 = ~n34364 & ~n34370;
  assign n34372 = ~n34358 & n34371;
  assign n34373 = n34369 ^ n34365;
  assign n34374 = n34359 & n34363;
  assign n34375 = ~n34373 & ~n34374;
  assign n34376 = n34375 ^ n34370;
  assign n34377 = ~n34372 & n34376;
  assign n34378 = n34377 ^ n33859;
  assign n34379 = n33860 & n34378;
  assign n34380 = n34379 ^ n33854;
  assign n34381 = n34380 ^ n33848;
  assign n34382 = ~n33849 & n34381;
  assign n34383 = n34382 ^ n33847;
  assign n34384 = n34383 ^ n33841;
  assign n34385 = ~n33842 & n34384;
  assign n34386 = n34385 ^ n33835;
  assign n34389 = n34388 ^ n34386;
  assign n34390 = n33940 ^ n32820;
  assign n34391 = n32820 ^ n32170;
  assign n34392 = n34390 & n34391;
  assign n34393 = n34392 ^ n32170;
  assign n34394 = n34393 ^ n34388;
  assign n34395 = ~n34389 & n34394;
  assign n34396 = n34395 ^ n34393;
  assign n34397 = n34396 ^ n33828;
  assign n34398 = n33829 & ~n34397;
  assign n34399 = n34398 ^ n33823;
  assign n34400 = n34399 ^ n33817;
  assign n34401 = ~n33818 & n34400;
  assign n34402 = n34401 ^ n33816;
  assign n34403 = n34402 ^ n33804;
  assign n34404 = ~n33805 & n34403;
  assign n34405 = n34404 ^ n33803;
  assign n34406 = n34405 ^ n33797;
  assign n34407 = ~n33798 & ~n34406;
  assign n34408 = n34407 ^ n33796;
  assign n34409 = n34408 ^ n33777;
  assign n34410 = ~n33787 & ~n34409;
  assign n34411 = n34410 ^ n33786;
  assign n34415 = n34414 ^ n34411;
  assign n34416 = n33882 ^ n33176;
  assign n34417 = n33176 ^ n32361;
  assign n34418 = n34416 & ~n34417;
  assign n34419 = n34418 ^ n32361;
  assign n34420 = n34419 ^ n34414;
  assign n34421 = ~n34415 & n34420;
  assign n34422 = n34421 ^ n34419;
  assign n34575 = n34430 ^ n34422;
  assign n34576 = n34431 & n34575;
  assign n34577 = n34576 ^ n34426;
  assign n34649 = n34585 ^ n34577;
  assign n34650 = ~n34586 & ~n34649;
  assign n34651 = n34650 ^ n34581;
  assign n34862 = n34659 ^ n34651;
  assign n34863 = n34660 & ~n34862;
  assign n34864 = n34863 ^ n34655;
  assign n34894 = n34872 ^ n34864;
  assign n34895 = n34873 & n34894;
  assign n34896 = n34895 ^ n34868;
  assign n34946 = n34905 ^ n34896;
  assign n34947 = ~n34945 & ~n34946;
  assign n34948 = n34947 ^ n34900;
  assign n34985 = n34955 ^ n34948;
  assign n34986 = n34984 & n34985;
  assign n34987 = n34986 ^ n34952;
  assign n34992 = n34991 ^ n34987;
  assign n34998 = n34997 ^ n34992;
  assign n34953 = n34952 ^ n34948;
  assign n34956 = n34955 ^ n34953;
  assign n34979 = n34956 ^ n30978;
  assign n34901 = n34900 ^ n34896;
  assign n34906 = n34905 ^ n34901;
  assign n34907 = n34906 ^ n30984;
  assign n34874 = n34873 ^ n34864;
  assign n34890 = n34874 ^ n30854;
  assign n34661 = n34660 ^ n34651;
  assign n34662 = n34661 ^ n30817;
  assign n34587 = n34586 ^ n34577;
  assign n34645 = n34587 ^ n30778;
  assign n34432 = n34431 ^ n34422;
  assign n34433 = n34432 ^ n31695;
  assign n34434 = n34419 ^ n34415;
  assign n34435 = n34434 ^ n31579;
  assign n34436 = n34408 ^ n33786;
  assign n34437 = n34436 ^ n33777;
  assign n34438 = n34437 ^ n31538;
  assign n34439 = n34405 ^ n33798;
  assign n34440 = n34439 ^ n31465;
  assign n34441 = n34402 ^ n33805;
  assign n34442 = n34441 ^ n31344;
  assign n34443 = n34399 ^ n33818;
  assign n34444 = n34443 ^ n31350;
  assign n34445 = n34396 ^ n33829;
  assign n34446 = n34445 ^ n31356;
  assign n34447 = n34393 ^ n34389;
  assign n34448 = n34447 ^ n31368;
  assign n34449 = n34383 ^ n33835;
  assign n34450 = n34449 ^ n33841;
  assign n34451 = n34450 ^ n31374;
  assign n34452 = n34380 ^ n33847;
  assign n34453 = n34452 ^ n33848;
  assign n34454 = n34453 ^ n31387;
  assign n34455 = n34377 ^ n33860;
  assign n34456 = n34455 ^ n31292;
  assign n34457 = n34363 ^ n34359;
  assign n34458 = n34363 ^ n34358;
  assign n34459 = n34457 & n34458;
  assign n34460 = n34459 ^ n34359;
  assign n34461 = n34460 ^ n34373;
  assign n34462 = n34461 ^ n31398;
  assign n34463 = n34457 ^ n34358;
  assign n34464 = n34463 ^ n31404;
  assign n34467 = n34466 ^ n34323;
  assign n34468 = n34353 & n34467;
  assign n34469 = n34468 ^ n34324;
  assign n34470 = n34469 ^ n34348;
  assign n34471 = n34470 ^ n31415;
  assign n34529 = n34528 ^ n34472;
  assign n34530 = n34473 & ~n34529;
  assign n34531 = n34530 ^ n31421;
  assign n34532 = n34531 ^ n34470;
  assign n34533 = n34471 & ~n34532;
  assign n34534 = n34533 ^ n31415;
  assign n34535 = n34534 ^ n34463;
  assign n34536 = n34464 & ~n34535;
  assign n34537 = n34536 ^ n31404;
  assign n34538 = n34537 ^ n34461;
  assign n34539 = n34462 & ~n34538;
  assign n34540 = n34539 ^ n31398;
  assign n34541 = n34540 ^ n34455;
  assign n34542 = n34456 & ~n34541;
  assign n34543 = n34542 ^ n31292;
  assign n34544 = n34543 ^ n34453;
  assign n34545 = n34454 & ~n34544;
  assign n34546 = n34545 ^ n31387;
  assign n34547 = n34546 ^ n34450;
  assign n34548 = ~n34451 & ~n34547;
  assign n34549 = n34548 ^ n31374;
  assign n34550 = n34549 ^ n34447;
  assign n34551 = ~n34448 & ~n34550;
  assign n34552 = n34551 ^ n31368;
  assign n34553 = n34552 ^ n34445;
  assign n34554 = n34446 & n34553;
  assign n34555 = n34554 ^ n31356;
  assign n34556 = n34555 ^ n34443;
  assign n34557 = n34444 & n34556;
  assign n34558 = n34557 ^ n31350;
  assign n34559 = n34558 ^ n34441;
  assign n34560 = ~n34442 & ~n34559;
  assign n34561 = n34560 ^ n31344;
  assign n34562 = n34561 ^ n34439;
  assign n34563 = ~n34440 & n34562;
  assign n34564 = n34563 ^ n31465;
  assign n34565 = n34564 ^ n34437;
  assign n34566 = n34438 & ~n34565;
  assign n34567 = n34566 ^ n31538;
  assign n34568 = n34567 ^ n34434;
  assign n34569 = ~n34435 & ~n34568;
  assign n34570 = n34569 ^ n31579;
  assign n34571 = n34570 ^ n34432;
  assign n34572 = n34433 & n34571;
  assign n34573 = n34572 ^ n31695;
  assign n34646 = n34587 ^ n34573;
  assign n34647 = ~n34645 & ~n34646;
  assign n34648 = n34647 ^ n30778;
  assign n34858 = n34661 ^ n34648;
  assign n34859 = ~n34662 & n34858;
  assign n34860 = n34859 ^ n30817;
  assign n34891 = n34874 ^ n34860;
  assign n34892 = n34890 & n34891;
  assign n34893 = n34892 ^ n30854;
  assign n34941 = n34906 ^ n34893;
  assign n34942 = ~n34907 & ~n34941;
  assign n34943 = n34942 ^ n30984;
  assign n34980 = n34956 ^ n34943;
  assign n34981 = n34979 & n34980;
  assign n34982 = n34981 ^ n30978;
  assign n34983 = n34982 ^ n30913;
  assign n34999 = n34998 ^ n34983;
  assign n34944 = n34943 ^ n30978;
  assign n34957 = n34956 ^ n34944;
  assign n34908 = n34907 ^ n34893;
  assign n34861 = n34860 ^ n30854;
  assign n34875 = n34874 ^ n34861;
  assign n34574 = n34573 ^ n30778;
  assign n34588 = n34587 ^ n34574;
  assign n34589 = n34570 ^ n34433;
  assign n34590 = n34567 ^ n31579;
  assign n34591 = n34590 ^ n34434;
  assign n34592 = n34561 ^ n31465;
  assign n34593 = n34592 ^ n34439;
  assign n34594 = n34555 ^ n31350;
  assign n34595 = n34594 ^ n34443;
  assign n34596 = n34546 ^ n34451;
  assign n34597 = n34540 ^ n31292;
  assign n34598 = n34597 ^ n34455;
  assign n34599 = n34531 ^ n31415;
  assign n34600 = n34599 ^ n34470;
  assign n34619 = n34601 & ~n34618;
  assign n34620 = n34600 & n34619;
  assign n34621 = n34534 ^ n34464;
  assign n34622 = n34620 & n34621;
  assign n34623 = n34537 ^ n31398;
  assign n34624 = n34623 ^ n34461;
  assign n34625 = n34622 & n34624;
  assign n34626 = ~n34598 & ~n34625;
  assign n34627 = n34543 ^ n31387;
  assign n34628 = n34627 ^ n34453;
  assign n34629 = ~n34626 & n34628;
  assign n34630 = ~n34596 & n34629;
  assign n34631 = n34549 ^ n31368;
  assign n34632 = n34631 ^ n34447;
  assign n34633 = n34630 & n34632;
  assign n34634 = n34552 ^ n34446;
  assign n34635 = ~n34633 & ~n34634;
  assign n34636 = ~n34595 & ~n34635;
  assign n34637 = n34558 ^ n34442;
  assign n34638 = n34636 & ~n34637;
  assign n34639 = ~n34593 & ~n34638;
  assign n34640 = n34564 ^ n34438;
  assign n34641 = n34639 & n34640;
  assign n34642 = ~n34591 & n34641;
  assign n34643 = n34589 & ~n34642;
  assign n34644 = n34588 & n34643;
  assign n34663 = n34662 ^ n34648;
  assign n34876 = n34644 & ~n34663;
  assign n34909 = n34875 & n34876;
  assign n34958 = ~n34908 & ~n34909;
  assign n35000 = ~n34957 & n34958;
  assign n35047 = n34999 & n35000;
  assign n35041 = n34998 ^ n30913;
  assign n35042 = n34998 ^ n34982;
  assign n35043 = n35041 & ~n35042;
  assign n35044 = n35043 ^ n30913;
  assign n35045 = n35044 ^ n31002;
  assign n35039 = n34230 ^ n34148;
  assign n35034 = n31990 ^ n31327;
  assign n35035 = n33371 ^ n31990;
  assign n35036 = ~n35034 & n35035;
  assign n35037 = n35036 ^ n31327;
  assign n35030 = n34997 ^ n34991;
  assign n35031 = n34997 ^ n34987;
  assign n35032 = ~n35030 & ~n35031;
  assign n35033 = n35032 ^ n34991;
  assign n35038 = n35037 ^ n35033;
  assign n35040 = n35039 ^ n35038;
  assign n35046 = n35045 ^ n35040;
  assign n35048 = n35047 ^ n35046;
  assign n35026 = n32369 ^ n2590;
  assign n35027 = n35026 ^ n28433;
  assign n35028 = n35027 ^ n23223;
  assign n35002 = n32499 ^ n2598;
  assign n35003 = n35002 ^ n28438;
  assign n35004 = n35003 ^ n2429;
  assign n35001 = n35000 ^ n34999;
  assign n35005 = n35004 ^ n35001;
  assign n34959 = n34958 ^ n34957;
  assign n34937 = n32494 ^ n24538;
  assign n34938 = n34937 ^ n2324;
  assign n34939 = n34938 ^ n23044;
  assign n34975 = n34959 ^ n34939;
  assign n34911 = n32472 ^ n24543;
  assign n34912 = n34911 ^ n28625;
  assign n34913 = n34912 ^ n2315;
  assign n34910 = n34909 ^ n34908;
  assign n34914 = n34913 ^ n34910;
  assign n34877 = n34876 ^ n34875;
  assign n34665 = n32466 ^ n24550;
  assign n34666 = n34665 ^ n1153;
  assign n34667 = n34666 ^ n1324;
  assign n34664 = n34663 ^ n34644;
  assign n34668 = n34667 ^ n34664;
  assign n34669 = n34643 ^ n34588;
  assign n1132 = n1125 ^ n1063;
  assign n1139 = n1138 ^ n1132;
  assign n1146 = n1145 ^ n1139;
  assign n34670 = n34669 ^ n1146;
  assign n34671 = n34642 ^ n34589;
  assign n1013 = n976 ^ n940;
  assign n1014 = n1013 ^ n1010;
  assign n1021 = n1020 ^ n1014;
  assign n34672 = n34671 ^ n1021;
  assign n34673 = n34641 ^ n34591;
  assign n980 = n964 ^ n932;
  assign n996 = n995 ^ n980;
  assign n1003 = n1002 ^ n996;
  assign n34674 = n34673 ^ n1003;
  assign n34675 = n34640 ^ n34639;
  assign n34679 = n34678 ^ n34675;
  assign n34681 = n32420 ^ n848;
  assign n34682 = n34681 ^ n28460;
  assign n34683 = n34682 ^ n23057;
  assign n34680 = n34638 ^ n34593;
  assign n34684 = n34683 ^ n34680;
  assign n34688 = n34637 ^ n34636;
  assign n34689 = n34688 ^ n34687;
  assign n34693 = n34635 ^ n34595;
  assign n34690 = n32387 ^ n24290;
  assign n34691 = n34690 ^ n28470;
  assign n34692 = n34691 ^ n554;
  assign n34694 = n34693 ^ n34692;
  assign n34698 = n34634 ^ n34633;
  assign n34695 = n32397 ^ n24157;
  assign n34696 = n34695 ^ n644;
  assign n34697 = n34696 ^ n23067;
  assign n34699 = n34698 ^ n34697;
  assign n34701 = n32391 ^ n24266;
  assign n34702 = n34701 ^ n28477;
  assign n34703 = n34702 ^ n639;
  assign n34700 = n34632 ^ n34630;
  assign n34704 = n34703 ^ n34700;
  assign n34820 = n34629 ^ n34596;
  assign n34705 = n34628 ^ n34626;
  assign n34709 = n34708 ^ n34705;
  assign n34710 = n34625 ^ n34598;
  assign n34714 = n34713 ^ n34710;
  assign n34715 = n34624 ^ n34622;
  assign n34719 = n34718 ^ n34715;
  assign n34723 = n34621 ^ n34620;
  assign n34724 = n34723 ^ n34722;
  assign n34725 = n34619 ^ n34600;
  assign n34726 = n34725 ^ n2147;
  assign n34802 = n34801 ^ n34727;
  assign n34803 = n34728 & ~n34802;
  assign n34804 = n34803 ^ n2132;
  assign n34805 = n34804 ^ n34725;
  assign n34806 = ~n34726 & n34805;
  assign n34807 = n34806 ^ n2147;
  assign n34808 = n34807 ^ n34723;
  assign n34809 = ~n34724 & n34808;
  assign n34810 = n34809 ^ n34722;
  assign n34811 = n34810 ^ n34715;
  assign n34812 = ~n34719 & n34811;
  assign n34813 = n34812 ^ n34718;
  assign n34814 = n34813 ^ n34710;
  assign n34815 = n34714 & ~n34814;
  assign n34816 = n34815 ^ n34713;
  assign n34817 = n34816 ^ n34705;
  assign n34818 = n34709 & ~n34817;
  assign n34819 = n34818 ^ n34708;
  assign n34821 = n34820 ^ n34819;
  assign n34825 = n34824 ^ n34820;
  assign n34826 = ~n34821 & n34825;
  assign n34827 = n34826 ^ n34824;
  assign n34828 = n34827 ^ n34700;
  assign n34829 = ~n34704 & n34828;
  assign n34830 = n34829 ^ n34703;
  assign n34831 = n34830 ^ n34698;
  assign n34832 = n34699 & ~n34831;
  assign n34833 = n34832 ^ n34697;
  assign n34834 = n34833 ^ n34693;
  assign n34835 = ~n34694 & n34834;
  assign n34836 = n34835 ^ n34692;
  assign n34837 = n34836 ^ n34688;
  assign n34838 = n34689 & ~n34837;
  assign n34839 = n34838 ^ n34687;
  assign n34840 = n34839 ^ n34680;
  assign n34841 = n34684 & ~n34840;
  assign n34842 = n34841 ^ n34683;
  assign n34843 = n34842 ^ n34675;
  assign n34844 = n34679 & ~n34843;
  assign n34845 = n34844 ^ n34678;
  assign n34846 = n34845 ^ n34673;
  assign n34847 = ~n34674 & n34846;
  assign n34848 = n34847 ^ n1003;
  assign n34849 = n34848 ^ n34671;
  assign n34850 = n34672 & ~n34849;
  assign n34851 = n34850 ^ n1021;
  assign n34852 = n34851 ^ n34669;
  assign n34853 = ~n34670 & n34852;
  assign n34854 = n34853 ^ n1146;
  assign n34855 = n34854 ^ n34664;
  assign n34856 = n34668 & ~n34855;
  assign n34857 = n34856 ^ n34667;
  assign n34878 = n34877 ^ n34857;
  assign n1317 = n1316 ^ n1229;
  assign n1330 = n1329 ^ n1317;
  assign n1337 = n1336 ^ n1330;
  assign n34887 = n34877 ^ n1337;
  assign n34888 = n34878 & ~n34887;
  assign n34889 = n34888 ^ n1337;
  assign n34934 = n34910 ^ n34889;
  assign n34935 = n34914 & ~n34934;
  assign n34936 = n34935 ^ n34913;
  assign n34976 = n34959 ^ n34936;
  assign n34977 = ~n34975 & n34976;
  assign n34978 = n34977 ^ n34939;
  assign n35023 = n35001 ^ n34978;
  assign n35024 = n35005 & ~n35023;
  assign n35025 = n35024 ^ n35004;
  assign n35029 = n35028 ^ n35025;
  assign n35049 = n35048 ^ n35029;
  assign n35019 = n33450 ^ n32759;
  assign n35020 = n34330 ^ n33450;
  assign n35021 = ~n35019 & ~n35020;
  assign n35022 = n35021 ^ n32759;
  assign n35050 = n35049 ^ n35022;
  assign n35006 = n35005 ^ n34978;
  assign n34971 = n33443 ^ n32767;
  assign n34972 = n34336 ^ n33443;
  assign n34973 = n34971 & n34972;
  assign n34974 = n34973 ^ n32767;
  assign n35007 = n35006 ^ n34974;
  assign n34940 = n34939 ^ n34936;
  assign n34960 = n34959 ^ n34940;
  assign n34930 = n33429 ^ n32739;
  assign n34931 = n33861 ^ n33429;
  assign n34932 = ~n34930 & ~n34931;
  assign n34933 = n34932 ^ n32739;
  assign n34961 = n34960 ^ n34933;
  assign n34879 = n34878 ^ n1337;
  assign n34880 = n32756 ^ n32628;
  assign n34881 = n33873 ^ n32756;
  assign n34882 = n34880 & ~n34881;
  assign n34883 = n34882 ^ n32628;
  assign n34920 = ~n34879 & ~n34883;
  assign n34916 = n33426 ^ n32650;
  assign n34917 = n33867 ^ n33426;
  assign n34918 = n34916 & n34917;
  assign n34919 = n34918 ^ n32650;
  assign n34921 = n34920 ^ n34919;
  assign n34915 = n34914 ^ n34889;
  assign n34927 = n34919 ^ n34915;
  assign n34928 = n34921 & ~n34927;
  assign n34929 = n34928 ^ n34920;
  assign n34968 = n34960 ^ n34929;
  assign n34969 = ~n34961 & n34968;
  assign n34970 = n34969 ^ n34933;
  assign n35016 = n35006 ^ n34970;
  assign n35017 = ~n35007 & ~n35016;
  assign n35018 = n35017 ^ n34974;
  assign n35096 = n35049 ^ n35018;
  assign n35097 = n35050 & n35096;
  assign n35098 = n35097 ^ n35022;
  assign n35294 = n35104 ^ n35098;
  assign n35295 = n35293 & n35294;
  assign n35296 = n35295 ^ n35102;
  assign n35297 = n35296 ^ n35287;
  assign n35298 = n35292 & n35297;
  assign n35299 = n35298 ^ n35291;
  assign n35300 = n35299 ^ n35281;
  assign n35301 = n35286 & n35300;
  assign n35302 = n35301 ^ n35285;
  assign n35303 = n35302 ^ n35279;
  assign n35304 = ~n35280 & n35303;
  assign n35305 = n35304 ^ n35277;
  assign n35151 = n34783 ^ n34753;
  assign n35152 = n35151 ^ n34754;
  assign n35306 = n35305 ^ n35152;
  assign n35307 = n33596 ^ n32941;
  assign n35308 = n33859 ^ n33596;
  assign n35309 = n35307 & ~n35308;
  assign n35310 = n35309 ^ n32941;
  assign n35311 = n35310 ^ n35152;
  assign n35312 = ~n35306 & ~n35311;
  assign n35313 = n35312 ^ n35310;
  assign n35314 = n35313 ^ n35145;
  assign n35315 = n35273 & n35314;
  assign n35316 = n35315 ^ n35272;
  assign n35317 = n35316 ^ n35267;
  assign n35318 = ~n35268 & ~n35317;
  assign n35319 = n35318 ^ n35266;
  assign n35320 = n35319 ^ n35137;
  assign n35321 = n35262 & n35320;
  assign n35322 = n35321 ^ n35261;
  assign n35323 = n35322 ^ n35128;
  assign n35324 = n35257 & n35323;
  assign n35325 = n35324 ^ n35256;
  assign n35326 = n35325 ^ n35122;
  assign n35327 = ~n35252 & n35326;
  assign n35328 = n35327 ^ n35251;
  assign n35329 = n35328 ^ n35113;
  assign n35330 = n35247 & ~n35329;
  assign n35331 = n35330 ^ n35246;
  assign n35240 = n34804 ^ n2147;
  assign n35241 = n35240 ^ n34725;
  assign n35236 = n33819 ^ n32826;
  assign n35237 = n33819 ^ n33797;
  assign n35238 = n35236 & n35237;
  assign n35239 = n35238 ^ n32826;
  assign n35242 = n35241 ^ n35239;
  assign n35404 = n35331 ^ n35242;
  assign n35405 = n35404 ^ n32129;
  assign n35406 = n35328 ^ n35247;
  assign n35407 = n35406 ^ n32108;
  assign n35408 = n35325 ^ n35252;
  assign n35409 = n35408 ^ n31290;
  assign n35410 = n35322 ^ n35256;
  assign n35411 = n35410 ^ n35128;
  assign n35412 = n35411 ^ n32076;
  assign n35413 = n35319 ^ n35262;
  assign n35414 = n35413 ^ n32059;
  assign n35415 = n35316 ^ n35268;
  assign n35416 = n35415 ^ n32019;
  assign n35417 = n35313 ^ n35273;
  assign n35418 = n35417 ^ n32025;
  assign n35419 = n35310 ^ n35306;
  assign n35420 = n35419 ^ n32035;
  assign n35421 = n35302 ^ n35277;
  assign n35422 = n35421 ^ n35279;
  assign n35423 = n35422 ^ n32009;
  assign n35424 = n35299 ^ n35285;
  assign n35425 = n35424 ^ n35281;
  assign n35426 = n35425 ^ n31967;
  assign n35427 = n35296 ^ n35291;
  assign n35428 = n35427 ^ n35287;
  assign n35429 = n35428 ^ n31838;
  assign n35103 = n35102 ^ n35098;
  assign n35105 = n35104 ^ n35103;
  assign n35106 = n35105 ^ n31766;
  assign n35051 = n35050 ^ n35018;
  assign n35092 = n35051 ^ n31298;
  assign n35008 = n35007 ^ n34970;
  assign n35009 = n35008 ^ n31304;
  assign n34962 = n34961 ^ n34929;
  assign n34964 = n34962 ^ n31310;
  assign n34884 = n34883 ^ n34879;
  assign n34885 = ~n30880 & n34884;
  assign n34886 = n34885 ^ n31312;
  assign n34922 = n34921 ^ n34915;
  assign n34923 = n34922 ^ n34885;
  assign n34924 = ~n34886 & ~n34923;
  assign n34925 = n34924 ^ n31312;
  assign n34965 = n34962 ^ n34925;
  assign n34966 = ~n34964 & ~n34965;
  assign n34967 = n34966 ^ n31310;
  assign n35012 = n35008 ^ n34967;
  assign n35013 = ~n35009 & n35012;
  assign n35014 = n35013 ^ n31304;
  assign n35093 = n35051 ^ n35014;
  assign n35094 = ~n35092 & n35093;
  assign n35095 = n35094 ^ n31298;
  assign n35430 = n35105 ^ n35095;
  assign n35431 = n35106 & ~n35430;
  assign n35432 = n35431 ^ n31766;
  assign n35433 = n35432 ^ n35428;
  assign n35434 = ~n35429 & n35433;
  assign n35435 = n35434 ^ n31838;
  assign n35436 = n35435 ^ n35425;
  assign n35437 = ~n35426 & ~n35436;
  assign n35438 = n35437 ^ n31967;
  assign n35439 = n35438 ^ n35422;
  assign n35440 = n35423 & n35439;
  assign n35441 = n35440 ^ n32009;
  assign n35442 = n35441 ^ n35419;
  assign n35443 = n35420 & ~n35442;
  assign n35444 = n35443 ^ n32035;
  assign n35445 = n35444 ^ n35417;
  assign n35446 = n35418 & ~n35445;
  assign n35447 = n35446 ^ n32025;
  assign n35448 = n35447 ^ n35415;
  assign n35449 = ~n35416 & ~n35448;
  assign n35450 = n35449 ^ n32019;
  assign n35451 = n35450 ^ n35413;
  assign n35452 = n35414 & n35451;
  assign n35453 = n35452 ^ n32059;
  assign n35454 = n35453 ^ n35411;
  assign n35455 = ~n35412 & n35454;
  assign n35456 = n35455 ^ n32076;
  assign n35457 = n35456 ^ n35408;
  assign n35458 = ~n35409 & n35457;
  assign n35459 = n35458 ^ n31290;
  assign n35460 = n35459 ^ n35406;
  assign n35461 = n35407 & ~n35460;
  assign n35462 = n35461 ^ n32108;
  assign n35463 = n35462 ^ n35404;
  assign n35464 = n35405 & ~n35463;
  assign n35465 = n35464 ^ n32129;
  assign n35332 = n35331 ^ n35241;
  assign n35333 = n35242 & n35332;
  assign n35334 = n35333 ^ n35239;
  assign n35233 = n34807 ^ n34722;
  assign n35234 = n35233 ^ n34723;
  assign n35229 = n33812 ^ n32820;
  assign n35230 = n33812 ^ n33777;
  assign n35231 = ~n35229 & ~n35230;
  assign n35232 = n35231 ^ n32820;
  assign n35235 = n35234 ^ n35232;
  assign n35402 = n35334 ^ n35235;
  assign n35403 = n35402 ^ n32170;
  assign n35559 = n35465 ^ n35403;
  assign n35529 = n35453 ^ n35412;
  assign n35530 = n35450 ^ n32059;
  assign n35531 = n35530 ^ n35413;
  assign n35532 = n35435 ^ n31967;
  assign n35533 = n35532 ^ n35425;
  assign n35534 = n35432 ^ n31838;
  assign n35535 = n35534 ^ n35428;
  assign n35107 = n35106 ^ n35095;
  assign n34926 = n34925 ^ n31310;
  assign n34963 = n34962 ^ n34926;
  assign n35010 = n35009 ^ n34967;
  assign n35011 = ~n34963 & n35010;
  assign n35015 = n35014 ^ n31298;
  assign n35052 = n35051 ^ n35015;
  assign n35108 = n35011 & n35052;
  assign n35536 = n35107 & ~n35108;
  assign n35537 = n35535 & ~n35536;
  assign n35538 = n35533 & n35537;
  assign n35539 = n35438 ^ n32009;
  assign n35540 = n35539 ^ n35422;
  assign n35541 = ~n35538 & ~n35540;
  assign n35542 = n35441 ^ n32035;
  assign n35543 = n35542 ^ n35419;
  assign n35544 = n35541 & n35543;
  assign n35545 = n35444 ^ n32025;
  assign n35546 = n35545 ^ n35417;
  assign n35547 = ~n35544 & ~n35546;
  assign n35548 = n35447 ^ n35416;
  assign n35549 = n35547 & n35548;
  assign n35550 = n35531 & n35549;
  assign n35551 = n35529 & n35550;
  assign n35552 = n35456 ^ n31290;
  assign n35553 = n35552 ^ n35408;
  assign n35554 = ~n35551 & ~n35553;
  assign n35555 = n35459 ^ n35407;
  assign n35556 = ~n35554 & ~n35555;
  assign n35557 = n35462 ^ n35405;
  assign n35558 = n35556 & ~n35557;
  assign n35633 = n35559 ^ n35558;
  assign n35637 = n35636 ^ n35633;
  assign n35638 = n35557 ^ n35556;
  assign n35642 = n35641 ^ n35638;
  assign n35643 = n35555 ^ n35554;
  assign n35647 = n35646 ^ n35643;
  assign n35651 = n35553 ^ n35551;
  assign n35648 = n33209 ^ n24980;
  assign n35649 = n35648 ^ n29314;
  assign n35650 = n35649 ^ n23865;
  assign n35652 = n35651 ^ n35650;
  assign n35653 = n35550 ^ n35529;
  assign n35657 = n35656 ^ n35653;
  assign n35658 = n35549 ^ n35531;
  assign n35662 = n35661 ^ n35658;
  assign n35664 = n33225 ^ n2236;
  assign n35665 = n35664 ^ n1997;
  assign n35666 = n35665 ^ n23452;
  assign n35663 = n35548 ^ n35547;
  assign n35667 = n35666 ^ n35663;
  assign n35668 = n35546 ^ n35544;
  assign n35672 = n35671 ^ n35668;
  assign n35673 = n35543 ^ n35541;
  assign n1827 = n1826 ^ n1775;
  assign n1840 = n1839 ^ n1827;
  assign n1847 = n1846 ^ n1840;
  assign n35674 = n35673 ^ n1847;
  assign n35678 = n35540 ^ n35538;
  assign n35679 = n35678 ^ n35677;
  assign n35680 = n35537 ^ n35533;
  assign n35681 = n35680 ^ n1737;
  assign n35685 = n35536 ^ n35535;
  assign n35682 = n32680 ^ n1636;
  assign n35683 = n35682 ^ n28794;
  assign n35684 = n35683 ^ n1724;
  assign n35686 = n35685 ^ n35684;
  assign n35109 = n35108 ^ n35107;
  assign n35110 = n35109 ^ n35091;
  assign n35053 = n35052 ^ n35011;
  assign n35057 = n35056 ^ n35053;
  assign n35058 = n35010 ^ n34963;
  assign n35062 = n35061 ^ n35058;
  assign n35063 = n32700 ^ n25014;
  assign n35064 = n35063 ^ n28816;
  assign n35065 = n35064 ^ n23397;
  assign n35066 = n35065 ^ n34963;
  assign n35070 = n33369 ^ n25336;
  assign n35071 = n35070 ^ n29449;
  assign n35072 = n35071 ^ n2648;
  assign n35073 = n34884 ^ n30880;
  assign n35074 = n35072 & ~n35073;
  assign n35067 = n32696 ^ n25010;
  assign n35068 = n35067 ^ n28811;
  assign n35069 = n35068 ^ n1553;
  assign n35075 = n35074 ^ n35069;
  assign n35076 = n34922 ^ n34886;
  assign n35077 = n35076 ^ n35069;
  assign n35078 = n35075 & n35077;
  assign n35079 = n35078 ^ n35074;
  assign n35080 = n35079 ^ n34963;
  assign n35081 = ~n35066 & n35080;
  assign n35082 = n35081 ^ n35065;
  assign n35083 = n35082 ^ n35058;
  assign n35084 = n35062 & ~n35083;
  assign n35085 = n35084 ^ n35061;
  assign n35086 = n35085 ^ n35053;
  assign n35087 = ~n35057 & n35086;
  assign n35088 = n35087 ^ n35056;
  assign n35687 = n35109 ^ n35088;
  assign n35688 = ~n35110 & n35687;
  assign n35689 = n35688 ^ n35091;
  assign n35690 = n35689 ^ n35685;
  assign n35691 = n35686 & ~n35690;
  assign n35692 = n35691 ^ n35684;
  assign n35693 = n35692 ^ n35680;
  assign n35694 = ~n35681 & n35693;
  assign n35695 = n35694 ^ n1737;
  assign n35696 = n35695 ^ n35678;
  assign n35697 = n35679 & ~n35696;
  assign n35698 = n35697 ^ n35677;
  assign n35699 = n35698 ^ n35673;
  assign n35700 = n35674 & ~n35699;
  assign n35701 = n35700 ^ n1847;
  assign n35702 = n35701 ^ n35668;
  assign n35703 = ~n35672 & n35702;
  assign n35704 = n35703 ^ n35671;
  assign n35705 = n35704 ^ n35663;
  assign n35706 = ~n35667 & n35705;
  assign n35707 = n35706 ^ n35666;
  assign n35708 = n35707 ^ n35658;
  assign n35709 = ~n35662 & n35708;
  assign n35710 = n35709 ^ n35661;
  assign n35711 = n35710 ^ n35653;
  assign n35712 = ~n35657 & n35711;
  assign n35713 = n35712 ^ n35656;
  assign n35714 = n35713 ^ n35651;
  assign n35715 = n35652 & ~n35714;
  assign n35716 = n35715 ^ n35650;
  assign n35717 = n35716 ^ n35643;
  assign n35718 = ~n35647 & n35717;
  assign n35719 = n35718 ^ n35646;
  assign n35720 = n35719 ^ n35638;
  assign n35721 = n35642 & ~n35720;
  assign n35722 = n35721 ^ n35641;
  assign n35723 = n35722 ^ n35633;
  assign n35724 = n35637 & ~n35723;
  assign n35725 = n35724 ^ n35636;
  assign n35629 = n33255 ^ n657;
  assign n35630 = n35629 ^ n29294;
  assign n35631 = n35630 ^ n23832;
  assign n35466 = n35465 ^ n35402;
  assign n35467 = n35403 & ~n35466;
  assign n35468 = n35467 ^ n32170;
  assign n35561 = n35468 ^ n32196;
  assign n35335 = n35334 ^ n35234;
  assign n35336 = ~n35235 & ~n35335;
  assign n35337 = n35336 ^ n35232;
  assign n35226 = n34810 ^ n34718;
  assign n35227 = n35226 ^ n34715;
  assign n35222 = n33799 ^ n32809;
  assign n35223 = n34414 ^ n33799;
  assign n35224 = n35222 & ~n35223;
  assign n35225 = n35224 ^ n32809;
  assign n35228 = n35227 ^ n35225;
  assign n35400 = n35337 ^ n35228;
  assign n35562 = n35561 ^ n35400;
  assign n35560 = n35558 & ~n35559;
  assign n35628 = n35562 ^ n35560;
  assign n35632 = n35631 ^ n35628;
  assign n36146 = n35725 ^ n35632;
  assign n36142 = n34997 ^ n34090;
  assign n35158 = n34845 ^ n34674;
  assign n36143 = n35158 ^ n34997;
  assign n36144 = n36142 & ~n36143;
  assign n36145 = n36144 ^ n34090;
  assign n36147 = n36146 ^ n36145;
  assign n36152 = n35722 ^ n35637;
  assign n36148 = n34955 ^ n34003;
  assign n35164 = n34842 ^ n34678;
  assign n35165 = n35164 ^ n34675;
  assign n36149 = n35165 ^ n34955;
  assign n36150 = ~n36148 & n36149;
  assign n36151 = n36150 ^ n34003;
  assign n36153 = n36152 ^ n36151;
  assign n36220 = n35719 ^ n35642;
  assign n36158 = n35716 ^ n35646;
  assign n36159 = n36158 ^ n35643;
  assign n36154 = n34872 ^ n33782;
  assign n35177 = n34836 ^ n34687;
  assign n35178 = n35177 ^ n34688;
  assign n36155 = n35178 ^ n34872;
  assign n36156 = ~n36154 & n36155;
  assign n36157 = n36156 ^ n33782;
  assign n36160 = n36159 ^ n36157;
  assign n36165 = n35713 ^ n35652;
  assign n36161 = n34659 ^ n33792;
  assign n35184 = n34833 ^ n34692;
  assign n35185 = n35184 ^ n34693;
  assign n36162 = n35185 ^ n34659;
  assign n36163 = n36161 & n36162;
  assign n36164 = n36163 ^ n33792;
  assign n36166 = n36165 ^ n36164;
  assign n36167 = n34585 ^ n33799;
  assign n35191 = n34830 ^ n34699;
  assign n36168 = n35191 ^ n34585;
  assign n36169 = ~n36167 & n36168;
  assign n36170 = n36169 ^ n33799;
  assign n36061 = n35710 ^ n35656;
  assign n36062 = n36061 ^ n35653;
  assign n36171 = n36170 ^ n36062;
  assign n36176 = n35707 ^ n35662;
  assign n36172 = n34430 ^ n33812;
  assign n35197 = n34827 ^ n34704;
  assign n36173 = n35197 ^ n34430;
  assign n36174 = n36172 & ~n36173;
  assign n36175 = n36174 ^ n33812;
  assign n36177 = n36176 ^ n36175;
  assign n36182 = n35704 ^ n35666;
  assign n36183 = n36182 ^ n35663;
  assign n36178 = n34414 ^ n33819;
  assign n35203 = n34824 ^ n34821;
  assign n36179 = n35203 ^ n34414;
  assign n36180 = ~n36178 & ~n36179;
  assign n36181 = n36180 ^ n33819;
  assign n36184 = n36183 ^ n36181;
  assign n36185 = n33831 ^ n33797;
  assign n35220 = n34813 ^ n34714;
  assign n36186 = n35220 ^ n33797;
  assign n36187 = ~n36185 & ~n36186;
  assign n36188 = n36187 ^ n33831;
  assign n36073 = n35698 ^ n1847;
  assign n36074 = n36073 ^ n35673;
  assign n36189 = n36188 ^ n36074;
  assign n36054 = n35695 ^ n35679;
  assign n36049 = n33843 ^ n33804;
  assign n36050 = n35227 ^ n33804;
  assign n36051 = ~n36049 & ~n36050;
  assign n36052 = n36051 ^ n33843;
  assign n36190 = n36054 ^ n36052;
  assign n35921 = n35692 ^ n1737;
  assign n35922 = n35921 ^ n35680;
  assign n35917 = n33850 ^ n33817;
  assign n35918 = n35234 ^ n33817;
  assign n35919 = n35917 & ~n35918;
  assign n35920 = n35919 ^ n33850;
  assign n35923 = n35922 ^ n35920;
  assign n35852 = n35689 ^ n35686;
  assign n35848 = n33908 ^ n33828;
  assign n35849 = n35241 ^ n33828;
  assign n35850 = n35848 & n35849;
  assign n35851 = n35850 ^ n33908;
  assign n35853 = n35852 ^ n35851;
  assign n35112 = n34388 ^ n33766;
  assign n35114 = n35113 ^ n34388;
  assign n35115 = ~n35112 & ~n35114;
  assign n35116 = n35115 ^ n33766;
  assign n35111 = n35110 ^ n35088;
  assign n35117 = n35116 ^ n35111;
  assign n35120 = n33841 ^ n33596;
  assign n35123 = n35122 ^ n33841;
  assign n35124 = ~n35120 & ~n35123;
  assign n35125 = n35124 ^ n33596;
  assign n35118 = n35085 ^ n35056;
  assign n35119 = n35118 ^ n35053;
  assign n35126 = n35125 ^ n35119;
  assign n35132 = n35082 ^ n35062;
  assign n35127 = n33848 ^ n33495;
  assign n35129 = n35128 ^ n33848;
  assign n35130 = n35127 & n35129;
  assign n35131 = n35130 ^ n33495;
  assign n35133 = n35132 ^ n35131;
  assign n35135 = n33859 ^ n32749;
  assign n35138 = n35137 ^ n33859;
  assign n35139 = ~n35135 & n35138;
  assign n35140 = n35139 ^ n32749;
  assign n35134 = n35079 ^ n35066;
  assign n35141 = n35140 ^ n35134;
  assign n35827 = n35076 ^ n35075;
  assign n35143 = n34359 ^ n33472;
  assign n35146 = n35145 ^ n34359;
  assign n35147 = n35143 & n35146;
  assign n35148 = n35147 ^ n33472;
  assign n35142 = n35073 ^ n35072;
  assign n35149 = n35148 ^ n35142;
  assign n35514 = n34851 ^ n34670;
  assign n35371 = n33371 ^ n32540;
  assign n35372 = n34284 ^ n33371;
  assign n35373 = n35371 & n35372;
  assign n35374 = n35373 ^ n32540;
  assign n35156 = n34848 ^ n1021;
  assign n35157 = n35156 ^ n34671;
  assign n35510 = n35374 ^ n35157;
  assign n35159 = n33375 ^ n32546;
  assign n35160 = n34290 ^ n33375;
  assign n35161 = ~n35159 & n35160;
  assign n35162 = n35161 ^ n32546;
  assign n35163 = n35162 ^ n35158;
  assign n35166 = n33385 ^ n32556;
  assign n35167 = n34292 ^ n33385;
  assign n35168 = n35166 & ~n35167;
  assign n35169 = n35168 ^ n32556;
  assign n35170 = n35169 ^ n35165;
  assign n35175 = n34839 ^ n34684;
  assign n35171 = n33387 ^ n32573;
  assign n35172 = n35039 ^ n33387;
  assign n35173 = ~n35171 & ~n35172;
  assign n35174 = n35173 ^ n32573;
  assign n35176 = n35175 ^ n35174;
  assign n35179 = n33397 ^ n32565;
  assign n35180 = n34997 ^ n33397;
  assign n35181 = ~n35179 & n35180;
  assign n35182 = n35181 ^ n32565;
  assign n35183 = n35182 ^ n35178;
  assign n35186 = n34254 ^ n33360;
  assign n35187 = n34955 ^ n34254;
  assign n35188 = ~n35186 & ~n35187;
  assign n35189 = n35188 ^ n33360;
  assign n35190 = n35189 ^ n35185;
  assign n35192 = n34090 ^ n33176;
  assign n35193 = n34905 ^ n34090;
  assign n35194 = n35192 & ~n35193;
  assign n35195 = n35194 ^ n33176;
  assign n35196 = n35195 ^ n35191;
  assign n35198 = n34003 ^ n32990;
  assign n35199 = n34872 ^ n34003;
  assign n35200 = ~n35198 & n35199;
  assign n35201 = n35200 ^ n32990;
  assign n35202 = n35201 ^ n35197;
  assign n35204 = n33882 ^ n32787;
  assign n35205 = n34659 ^ n33882;
  assign n35206 = n35204 & ~n35205;
  assign n35207 = n35206 ^ n32787;
  assign n35208 = n35207 ^ n35203;
  assign n35211 = n33782 ^ n32793;
  assign n35212 = n34585 ^ n33782;
  assign n35213 = n35211 & n35212;
  assign n35214 = n35213 ^ n32793;
  assign n35209 = n34816 ^ n34708;
  assign n35210 = n35209 ^ n34705;
  assign n35215 = n35214 ^ n35210;
  assign n35216 = n33792 ^ n32799;
  assign n35217 = n34430 ^ n33792;
  assign n35218 = ~n35216 & n35217;
  assign n35219 = n35218 ^ n32799;
  assign n35221 = n35220 ^ n35219;
  assign n35338 = n35337 ^ n35227;
  assign n35339 = ~n35228 & n35338;
  assign n35340 = n35339 ^ n35225;
  assign n35341 = n35340 ^ n35220;
  assign n35342 = ~n35221 & ~n35341;
  assign n35343 = n35342 ^ n35219;
  assign n35344 = n35343 ^ n35210;
  assign n35345 = n35215 & n35344;
  assign n35346 = n35345 ^ n35214;
  assign n35347 = n35346 ^ n35203;
  assign n35348 = n35208 & ~n35347;
  assign n35349 = n35348 ^ n35207;
  assign n35350 = n35349 ^ n35197;
  assign n35351 = n35202 & n35350;
  assign n35352 = n35351 ^ n35201;
  assign n35353 = n35352 ^ n35191;
  assign n35354 = ~n35196 & n35353;
  assign n35355 = n35354 ^ n35195;
  assign n35356 = n35355 ^ n35185;
  assign n35357 = ~n35190 & ~n35356;
  assign n35358 = n35357 ^ n35189;
  assign n35359 = n35358 ^ n35178;
  assign n35360 = ~n35183 & ~n35359;
  assign n35361 = n35360 ^ n35182;
  assign n35362 = n35361 ^ n35175;
  assign n35363 = ~n35176 & n35362;
  assign n35364 = n35363 ^ n35174;
  assign n35365 = n35364 ^ n35165;
  assign n35366 = ~n35170 & n35365;
  assign n35367 = n35366 ^ n35169;
  assign n35368 = n35367 ^ n35158;
  assign n35369 = ~n35163 & ~n35368;
  assign n35370 = n35369 ^ n35162;
  assign n35511 = n35370 ^ n35157;
  assign n35512 = n35510 & ~n35511;
  assign n35513 = n35512 ^ n35374;
  assign n35515 = n35514 ^ n35513;
  assign n35506 = n32765 ^ n31996;
  assign n35507 = n34278 ^ n32765;
  assign n35508 = n35506 & ~n35507;
  assign n35509 = n35508 ^ n31996;
  assign n35516 = n35515 ^ n35509;
  assign n35375 = n35374 ^ n35370;
  assign n35376 = n35375 ^ n35157;
  assign n35377 = n35376 ^ n31703;
  assign n35378 = n35367 ^ n35162;
  assign n35379 = n35378 ^ n35158;
  assign n35380 = n35379 ^ n31713;
  assign n35381 = n35364 ^ n35169;
  assign n35382 = n35381 ^ n35165;
  assign n35383 = n35382 ^ n31715;
  assign n35384 = n35361 ^ n35176;
  assign n35385 = n35384 ^ n31725;
  assign n35386 = n35358 ^ n35183;
  assign n35387 = n35386 ^ n31727;
  assign n35388 = n35355 ^ n35190;
  assign n35389 = n35388 ^ n32527;
  assign n35390 = n35352 ^ n35196;
  assign n35391 = n35390 ^ n32361;
  assign n35392 = n35349 ^ n35202;
  assign n35393 = n35392 ^ n32274;
  assign n35394 = n35346 ^ n35208;
  assign n35395 = n35394 ^ n32257;
  assign n35396 = n35343 ^ n35215;
  assign n35397 = n35396 ^ n32223;
  assign n35398 = n35340 ^ n35221;
  assign n35399 = n35398 ^ n32205;
  assign n35401 = n35400 ^ n32196;
  assign n35469 = n35468 ^ n35400;
  assign n35470 = ~n35401 & n35469;
  assign n35471 = n35470 ^ n32196;
  assign n35472 = n35471 ^ n35398;
  assign n35473 = ~n35399 & n35472;
  assign n35474 = n35473 ^ n32205;
  assign n35475 = n35474 ^ n35396;
  assign n35476 = ~n35397 & n35475;
  assign n35477 = n35476 ^ n32223;
  assign n35478 = n35477 ^ n35394;
  assign n35479 = ~n35395 & ~n35478;
  assign n35480 = n35479 ^ n32257;
  assign n35481 = n35480 ^ n35392;
  assign n35482 = n35393 & n35481;
  assign n35483 = n35482 ^ n32274;
  assign n35484 = n35483 ^ n35390;
  assign n35485 = n35391 & ~n35484;
  assign n35486 = n35485 ^ n32361;
  assign n35487 = n35486 ^ n35388;
  assign n35488 = ~n35389 & ~n35487;
  assign n35489 = n35488 ^ n32527;
  assign n35490 = n35489 ^ n35386;
  assign n35491 = ~n35387 & ~n35490;
  assign n35492 = n35491 ^ n31727;
  assign n35493 = n35492 ^ n35384;
  assign n35494 = n35385 & ~n35493;
  assign n35495 = n35494 ^ n31725;
  assign n35496 = n35495 ^ n35382;
  assign n35497 = ~n35383 & ~n35496;
  assign n35498 = n35497 ^ n31715;
  assign n35499 = n35498 ^ n35379;
  assign n35500 = n35380 & n35499;
  assign n35501 = n35500 ^ n31713;
  assign n35502 = n35501 ^ n35376;
  assign n35503 = ~n35377 & ~n35502;
  assign n35504 = n35503 ^ n31703;
  assign n35505 = n35504 ^ n31333;
  assign n35517 = n35516 ^ n35505;
  assign n35518 = n35501 ^ n31703;
  assign n35519 = n35518 ^ n35376;
  assign n35520 = n35489 ^ n35387;
  assign n35521 = n35486 ^ n35389;
  assign n35522 = n35483 ^ n35391;
  assign n35523 = n35480 ^ n32274;
  assign n35524 = n35523 ^ n35392;
  assign n35525 = n35477 ^ n35395;
  assign n35526 = n35474 ^ n32223;
  assign n35527 = n35526 ^ n35396;
  assign n35528 = n35471 ^ n35399;
  assign n35563 = ~n35560 & ~n35562;
  assign n35564 = n35528 & ~n35563;
  assign n35565 = n35527 & n35564;
  assign n35566 = ~n35525 & ~n35565;
  assign n35567 = ~n35524 & n35566;
  assign n35568 = n35522 & n35567;
  assign n35569 = n35521 & ~n35568;
  assign n35570 = ~n35520 & n35569;
  assign n35571 = n35492 ^ n31725;
  assign n35572 = n35571 ^ n35384;
  assign n35573 = n35570 & ~n35572;
  assign n35574 = n35495 ^ n35383;
  assign n35575 = n35573 & n35574;
  assign n35576 = n35498 ^ n31713;
  assign n35577 = n35576 ^ n35379;
  assign n35578 = ~n35575 & ~n35577;
  assign n35579 = ~n35519 & n35578;
  assign n35782 = ~n35517 & n35579;
  assign n35779 = n34854 ^ n34668;
  assign n35774 = n32763 ^ n31990;
  assign n35775 = n34265 ^ n32763;
  assign n35776 = n35774 & n35775;
  assign n35777 = n35776 ^ n31990;
  assign n35771 = n35514 ^ n35509;
  assign n35772 = n35515 & n35771;
  assign n35773 = n35772 ^ n35509;
  assign n35778 = n35777 ^ n35773;
  assign n35780 = n35779 ^ n35778;
  assign n35766 = n35516 ^ n31333;
  assign n35767 = n35516 ^ n35504;
  assign n35768 = n35766 & n35767;
  assign n35769 = n35768 ^ n31333;
  assign n35770 = n35769 ^ n31327;
  assign n35781 = n35780 ^ n35770;
  assign n35783 = n35782 ^ n35781;
  assign n35581 = n33189 ^ n25211;
  assign n35582 = n35581 ^ n2404;
  assign n35583 = n35582 ^ n2497;
  assign n35580 = n35579 ^ n35517;
  assign n35584 = n35583 ^ n35580;
  assign n35585 = n35578 ^ n35519;
  assign n2371 = n2357 ^ n2337;
  assign n2390 = n2389 ^ n2371;
  assign n2397 = n2396 ^ n2390;
  assign n35586 = n35585 ^ n2397;
  assign n35588 = n2295 ^ n1360;
  assign n35589 = n35588 ^ n29264;
  assign n35590 = n35589 ^ n2384;
  assign n35587 = n35577 ^ n35575;
  assign n35591 = n35590 ^ n35587;
  assign n35593 = n2300 ^ n1345;
  assign n35594 = n35593 ^ n1299;
  assign n35595 = n35594 ^ n23810;
  assign n35592 = n35574 ^ n35573;
  assign n35596 = n35595 ^ n35592;
  assign n35597 = n35572 ^ n35570;
  assign n1284 = n1244 ^ n1187;
  assign n1285 = n1284 ^ n1281;
  assign n1289 = n1288 ^ n1285;
  assign n35598 = n35597 ^ n1289;
  assign n35599 = n35569 ^ n35520;
  assign n1257 = n1172 ^ n1106;
  assign n1267 = n1266 ^ n1257;
  assign n1274 = n1273 ^ n1267;
  assign n35600 = n35599 ^ n1274;
  assign n35601 = n35568 ^ n35521;
  assign n35605 = n35604 ^ n35601;
  assign n35606 = n35567 ^ n35522;
  assign n35610 = n35609 ^ n35606;
  assign n35614 = n35566 ^ n35524;
  assign n35615 = n35614 ^ n35613;
  assign n35617 = n33280 ^ n24958;
  assign n35618 = n35617 ^ n29282;
  assign n35619 = n35618 ^ n768;
  assign n35616 = n35565 ^ n35525;
  assign n35620 = n35619 ^ n35616;
  assign n35621 = n35564 ^ n35527;
  assign n681 = n680 ^ n569;
  assign n700 = n699 ^ n681;
  assign n707 = n706 ^ n700;
  assign n35622 = n35621 ^ n707;
  assign n35626 = n35563 ^ n35528;
  assign n35623 = n29289 ^ n25080;
  assign n35624 = n35623 ^ n33250;
  assign n35625 = n35624 ^ n694;
  assign n35627 = n35626 ^ n35625;
  assign n35726 = n35725 ^ n35628;
  assign n35727 = n35632 & ~n35726;
  assign n35728 = n35727 ^ n35631;
  assign n35729 = n35728 ^ n35626;
  assign n35730 = n35627 & ~n35729;
  assign n35731 = n35730 ^ n35625;
  assign n35732 = n35731 ^ n35621;
  assign n35733 = ~n35622 & n35732;
  assign n35734 = n35733 ^ n707;
  assign n35735 = n35734 ^ n35616;
  assign n35736 = n35620 & ~n35735;
  assign n35737 = n35736 ^ n35619;
  assign n35738 = n35737 ^ n35614;
  assign n35739 = ~n35615 & n35738;
  assign n35740 = n35739 ^ n35613;
  assign n35741 = n35740 ^ n35606;
  assign n35742 = n35610 & ~n35741;
  assign n35743 = n35742 ^ n35609;
  assign n35744 = n35743 ^ n35601;
  assign n35745 = n35605 & ~n35744;
  assign n35746 = n35745 ^ n35604;
  assign n35747 = n35746 ^ n35599;
  assign n35748 = n35600 & ~n35747;
  assign n35749 = n35748 ^ n1274;
  assign n35750 = n35749 ^ n35597;
  assign n35751 = n35598 & ~n35750;
  assign n35752 = n35751 ^ n1289;
  assign n35753 = n35752 ^ n35592;
  assign n35754 = ~n35596 & n35753;
  assign n35755 = n35754 ^ n35595;
  assign n35756 = n35755 ^ n35587;
  assign n35757 = n35591 & ~n35756;
  assign n35758 = n35757 ^ n35590;
  assign n35759 = n35758 ^ n35585;
  assign n35760 = ~n35586 & n35759;
  assign n35761 = n35760 ^ n2397;
  assign n35762 = n35761 ^ n35580;
  assign n35763 = ~n35584 & n35762;
  assign n35764 = n35763 ^ n35583;
  assign n2493 = n2492 ^ n2432;
  assign n2500 = n2499 ^ n2493;
  assign n2501 = n2500 ^ n2480;
  assign n35765 = n35764 ^ n2501;
  assign n35784 = n35783 ^ n35765;
  assign n35150 = n34343 ^ n33450;
  assign n35153 = n35152 ^ n34343;
  assign n35154 = ~n35150 & n35153;
  assign n35155 = n35154 ^ n33450;
  assign n35785 = n35784 ^ n35155;
  assign n35790 = n35761 ^ n35584;
  assign n35786 = n34324 ^ n33443;
  assign n35787 = n35279 ^ n34324;
  assign n35788 = ~n35786 & ~n35787;
  assign n35789 = n35788 ^ n33443;
  assign n35791 = n35790 ^ n35789;
  assign n35796 = n35758 ^ n2397;
  assign n35797 = n35796 ^ n35585;
  assign n35792 = n34330 ^ n33429;
  assign n35793 = n35281 ^ n34330;
  assign n35794 = n35792 & ~n35793;
  assign n35795 = n35794 ^ n33429;
  assign n35798 = n35797 ^ n35795;
  assign n35803 = n35755 ^ n35591;
  assign n35799 = n34336 ^ n33426;
  assign n35800 = n35287 ^ n34336;
  assign n35801 = n35799 & ~n35800;
  assign n35802 = n35801 ^ n33426;
  assign n35804 = n35803 ^ n35802;
  assign n35805 = n35752 ^ n35595;
  assign n35806 = n35805 ^ n35592;
  assign n35807 = n33861 ^ n32756;
  assign n35808 = n35104 ^ n33861;
  assign n35809 = n35807 & ~n35808;
  assign n35810 = n35809 ^ n32756;
  assign n35811 = ~n35806 & ~n35810;
  assign n35812 = n35811 ^ n35803;
  assign n35813 = ~n35804 & n35812;
  assign n35814 = n35813 ^ n35811;
  assign n35815 = n35814 ^ n35797;
  assign n35816 = n35798 & n35815;
  assign n35817 = n35816 ^ n35795;
  assign n35818 = n35817 ^ n35790;
  assign n35819 = n35791 & ~n35818;
  assign n35820 = n35819 ^ n35789;
  assign n35821 = n35820 ^ n35784;
  assign n35822 = n35785 & ~n35821;
  assign n35823 = n35822 ^ n35155;
  assign n35824 = n35823 ^ n35142;
  assign n35825 = ~n35149 & ~n35824;
  assign n35826 = n35825 ^ n35148;
  assign n35828 = n35827 ^ n35826;
  assign n35829 = n34365 ^ n33478;
  assign n35830 = n35267 ^ n34365;
  assign n35831 = n35829 & ~n35830;
  assign n35832 = n35831 ^ n33478;
  assign n35833 = n35832 ^ n35827;
  assign n35834 = n35828 & n35833;
  assign n35835 = n35834 ^ n35832;
  assign n35836 = n35835 ^ n35134;
  assign n35837 = n35141 & ~n35836;
  assign n35838 = n35837 ^ n35140;
  assign n35839 = n35838 ^ n35132;
  assign n35840 = ~n35133 & n35839;
  assign n35841 = n35840 ^ n35131;
  assign n35842 = n35841 ^ n35119;
  assign n35843 = ~n35126 & ~n35842;
  assign n35844 = n35843 ^ n35125;
  assign n35845 = n35844 ^ n35111;
  assign n35846 = n35117 & n35845;
  assign n35847 = n35846 ^ n35116;
  assign n35914 = n35852 ^ n35847;
  assign n35915 = n35853 & n35914;
  assign n35916 = n35915 ^ n35851;
  assign n36046 = n35922 ^ n35916;
  assign n36047 = n35923 & n36046;
  assign n36048 = n36047 ^ n35920;
  assign n36191 = n36054 ^ n36048;
  assign n36192 = n36190 & n36191;
  assign n36193 = n36192 ^ n36052;
  assign n36194 = n36193 ^ n36074;
  assign n36195 = ~n36189 & ~n36194;
  assign n36196 = n36195 ^ n36188;
  assign n36065 = n35701 ^ n35672;
  assign n36197 = n36196 ^ n36065;
  assign n36198 = n33940 ^ n33777;
  assign n36199 = n35210 ^ n33777;
  assign n36200 = n36198 & n36199;
  assign n36201 = n36200 ^ n33940;
  assign n36202 = n36201 ^ n36065;
  assign n36203 = ~n36197 & n36202;
  assign n36204 = n36203 ^ n36201;
  assign n36205 = n36204 ^ n36183;
  assign n36206 = n36184 & ~n36205;
  assign n36207 = n36206 ^ n36181;
  assign n36208 = n36207 ^ n36176;
  assign n36209 = n36177 & ~n36208;
  assign n36210 = n36209 ^ n36175;
  assign n36211 = n36210 ^ n36062;
  assign n36212 = ~n36171 & ~n36211;
  assign n36213 = n36212 ^ n36170;
  assign n36214 = n36213 ^ n36165;
  assign n36215 = n36166 & ~n36214;
  assign n36216 = n36215 ^ n36164;
  assign n36217 = n36216 ^ n36159;
  assign n36218 = ~n36160 & n36217;
  assign n36219 = n36218 ^ n36157;
  assign n36221 = n36220 ^ n36219;
  assign n36222 = n34905 ^ n33882;
  assign n36223 = n35175 ^ n34905;
  assign n36224 = ~n36222 & n36223;
  assign n36225 = n36224 ^ n33882;
  assign n36226 = n36225 ^ n36220;
  assign n36227 = ~n36221 & n36226;
  assign n36228 = n36227 ^ n36225;
  assign n36229 = n36228 ^ n36152;
  assign n36230 = n36153 & ~n36229;
  assign n36231 = n36230 ^ n36151;
  assign n36232 = n36231 ^ n36146;
  assign n36233 = ~n36147 & ~n36232;
  assign n36234 = n36233 ^ n36145;
  assign n36135 = n35039 ^ n34254;
  assign n36136 = n35157 ^ n35039;
  assign n36137 = ~n36135 & ~n36136;
  assign n36138 = n36137 ^ n34254;
  assign n36267 = n36234 ^ n36138;
  assign n36139 = n35728 ^ n35625;
  assign n36140 = n36139 ^ n35626;
  assign n36268 = n36267 ^ n36140;
  assign n36269 = n36268 ^ n33360;
  assign n36270 = n36231 ^ n36147;
  assign n36271 = n36270 ^ n33176;
  assign n36272 = n36228 ^ n36153;
  assign n36273 = n36272 ^ n32990;
  assign n36274 = n36225 ^ n36221;
  assign n36275 = n36274 ^ n32787;
  assign n36276 = n36216 ^ n36157;
  assign n36277 = n36276 ^ n36159;
  assign n36278 = n36277 ^ n32793;
  assign n36310 = n36213 ^ n36164;
  assign n36311 = n36310 ^ n36165;
  assign n36279 = n36210 ^ n36170;
  assign n36280 = n36279 ^ n36062;
  assign n36281 = n36280 ^ n32809;
  assign n36282 = n36207 ^ n36175;
  assign n36283 = n36282 ^ n36176;
  assign n36284 = n36283 ^ n32820;
  assign n36285 = n36204 ^ n36181;
  assign n36286 = n36285 ^ n36183;
  assign n36287 = n36286 ^ n32826;
  assign n36288 = n36201 ^ n36197;
  assign n36289 = n36288 ^ n32836;
  assign n36290 = n36193 ^ n36189;
  assign n36291 = n36290 ^ n32842;
  assign n36053 = n36052 ^ n36048;
  assign n36055 = n36054 ^ n36053;
  assign n36056 = n36055 ^ n32844;
  assign n35924 = n35923 ^ n35916;
  assign n36042 = n35924 ^ n31982;
  assign n35854 = n35853 ^ n35847;
  assign n35855 = n35854 ^ n32859;
  assign n35856 = n35844 ^ n35117;
  assign n35857 = n35856 ^ n32947;
  assign n35858 = n35841 ^ n35125;
  assign n35859 = n35858 ^ n35119;
  assign n35860 = n35859 ^ n32941;
  assign n35861 = n35838 ^ n35133;
  assign n35862 = n35861 ^ n32865;
  assign n35863 = n35835 ^ n35141;
  assign n35864 = n35863 ^ n32871;
  assign n35865 = n35832 ^ n35828;
  assign n35866 = n35865 ^ n32877;
  assign n35867 = n35823 ^ n35149;
  assign n35868 = n35867 ^ n32752;
  assign n35869 = n35820 ^ n35785;
  assign n35870 = n35869 ^ n32759;
  assign n35871 = n35817 ^ n35791;
  assign n35872 = n35871 ^ n32767;
  assign n35873 = n35814 ^ n35798;
  assign n35874 = n35873 ^ n32739;
  assign n35875 = n35810 ^ n35806;
  assign n35876 = ~n32628 & n35875;
  assign n35877 = n35876 ^ n32650;
  assign n35878 = n35811 ^ n35802;
  assign n35879 = n35878 ^ n35803;
  assign n35880 = n35879 ^ n35876;
  assign n35881 = n35877 & ~n35880;
  assign n35882 = n35881 ^ n32650;
  assign n35883 = n35882 ^ n35873;
  assign n35884 = n35874 & ~n35883;
  assign n35885 = n35884 ^ n32739;
  assign n35886 = n35885 ^ n35871;
  assign n35887 = n35872 & n35886;
  assign n35888 = n35887 ^ n32767;
  assign n35889 = n35888 ^ n35869;
  assign n35890 = ~n35870 & ~n35889;
  assign n35891 = n35890 ^ n32759;
  assign n35892 = n35891 ^ n35867;
  assign n35893 = ~n35868 & ~n35892;
  assign n35894 = n35893 ^ n32752;
  assign n35895 = n35894 ^ n35865;
  assign n35896 = n35866 & n35895;
  assign n35897 = n35896 ^ n32877;
  assign n35898 = n35897 ^ n35863;
  assign n35899 = n35864 & n35898;
  assign n35900 = n35899 ^ n32871;
  assign n35901 = n35900 ^ n35861;
  assign n35902 = ~n35862 & n35901;
  assign n35903 = n35902 ^ n32865;
  assign n35904 = n35903 ^ n35859;
  assign n35905 = n35860 & n35904;
  assign n35906 = n35905 ^ n32941;
  assign n35907 = n35906 ^ n35856;
  assign n35908 = ~n35857 & ~n35907;
  assign n35909 = n35908 ^ n32947;
  assign n35910 = n35909 ^ n35854;
  assign n35911 = ~n35855 & ~n35910;
  assign n35912 = n35911 ^ n32859;
  assign n36043 = n35924 ^ n35912;
  assign n36044 = ~n36042 & ~n36043;
  assign n36045 = n36044 ^ n31982;
  assign n36292 = n36055 ^ n36045;
  assign n36293 = ~n36056 & ~n36292;
  assign n36294 = n36293 ^ n32844;
  assign n36295 = n36294 ^ n36290;
  assign n36296 = ~n36291 & n36295;
  assign n36297 = n36296 ^ n32842;
  assign n36298 = n36297 ^ n36288;
  assign n36299 = ~n36289 & n36298;
  assign n36300 = n36299 ^ n32836;
  assign n36301 = n36300 ^ n36286;
  assign n36302 = n36287 & n36301;
  assign n36303 = n36302 ^ n32826;
  assign n36304 = n36303 ^ n36283;
  assign n36305 = ~n36284 & ~n36304;
  assign n36306 = n36305 ^ n32820;
  assign n36307 = n36306 ^ n36280;
  assign n36308 = n36281 & ~n36307;
  assign n36309 = n36308 ^ n32809;
  assign n36312 = n36311 ^ n36309;
  assign n36313 = n36311 ^ n32799;
  assign n36314 = ~n36312 & ~n36313;
  assign n36315 = n36314 ^ n32799;
  assign n36316 = n36315 ^ n36277;
  assign n36317 = ~n36278 & ~n36316;
  assign n36318 = n36317 ^ n32793;
  assign n36319 = n36318 ^ n36274;
  assign n36320 = n36275 & ~n36319;
  assign n36321 = n36320 ^ n32787;
  assign n36322 = n36321 ^ n36272;
  assign n36323 = ~n36273 & ~n36322;
  assign n36324 = n36323 ^ n32990;
  assign n36325 = n36324 ^ n36270;
  assign n36326 = n36271 & ~n36325;
  assign n36327 = n36326 ^ n33176;
  assign n36328 = n36327 ^ n36268;
  assign n36329 = n36269 & n36328;
  assign n36330 = n36329 ^ n33360;
  assign n36141 = n36140 ^ n36138;
  assign n36235 = n36234 ^ n36140;
  assign n36236 = ~n36141 & n36235;
  assign n36237 = n36236 ^ n36138;
  assign n36132 = n35731 ^ n707;
  assign n36133 = n36132 ^ n35621;
  assign n36128 = n34292 ^ n33397;
  assign n36129 = n35514 ^ n34292;
  assign n36130 = ~n36128 & ~n36129;
  assign n36131 = n36130 ^ n33397;
  assign n36134 = n36133 ^ n36131;
  assign n36265 = n36237 ^ n36134;
  assign n36266 = n36265 ^ n32565;
  assign n36364 = n36330 ^ n36266;
  assign n36365 = n36327 ^ n36269;
  assign n36366 = n36324 ^ n36271;
  assign n36367 = n36318 ^ n32787;
  assign n36368 = n36367 ^ n36274;
  assign n36369 = n36315 ^ n32793;
  assign n36370 = n36369 ^ n36277;
  assign n36371 = n36297 ^ n36289;
  assign n36057 = n36056 ^ n36045;
  assign n35913 = n35912 ^ n31982;
  assign n35925 = n35924 ^ n35913;
  assign n35926 = n35906 ^ n32947;
  assign n35927 = n35926 ^ n35856;
  assign n35928 = n35903 ^ n35860;
  assign n35929 = n35900 ^ n32865;
  assign n35930 = n35929 ^ n35861;
  assign n35931 = n35897 ^ n35864;
  assign n35932 = n35891 ^ n35868;
  assign n35933 = n35888 ^ n32759;
  assign n35934 = n35933 ^ n35869;
  assign n35935 = n35882 ^ n32739;
  assign n35936 = n35935 ^ n35873;
  assign n35937 = n35885 ^ n35872;
  assign n35938 = ~n35936 & ~n35937;
  assign n35939 = ~n35934 & n35938;
  assign n35940 = ~n35932 & ~n35939;
  assign n35941 = n35894 ^ n32877;
  assign n35942 = n35941 ^ n35865;
  assign n35943 = ~n35940 & n35942;
  assign n35944 = ~n35931 & n35943;
  assign n35945 = n35930 & ~n35944;
  assign n35946 = ~n35928 & n35945;
  assign n35947 = n35927 & ~n35946;
  assign n35948 = n35909 ^ n35855;
  assign n35949 = n35947 & ~n35948;
  assign n36058 = n35925 & n35949;
  assign n36372 = ~n36057 & n36058;
  assign n36373 = n36294 ^ n32842;
  assign n36374 = n36373 ^ n36290;
  assign n36375 = ~n36372 & ~n36374;
  assign n36376 = n36371 & ~n36375;
  assign n36377 = n36300 ^ n36287;
  assign n36378 = n36376 & ~n36377;
  assign n36379 = n36303 ^ n32820;
  assign n36380 = n36379 ^ n36283;
  assign n36381 = n36378 & ~n36380;
  assign n36382 = n36306 ^ n32809;
  assign n36383 = n36382 ^ n36280;
  assign n36384 = ~n36381 & n36383;
  assign n36385 = n36312 ^ n32799;
  assign n36386 = ~n36384 & n36385;
  assign n36387 = ~n36370 & n36386;
  assign n36388 = n36368 & ~n36387;
  assign n36389 = n36321 ^ n32990;
  assign n36390 = n36389 ^ n36272;
  assign n36391 = n36388 & ~n36390;
  assign n36392 = ~n36366 & n36391;
  assign n36393 = n36365 & ~n36392;
  assign n36394 = n36364 & n36393;
  assign n36331 = n36330 ^ n36265;
  assign n36332 = ~n36266 & ~n36331;
  assign n36333 = n36332 ^ n32565;
  assign n36362 = n36333 ^ n32573;
  assign n36238 = n36237 ^ n36133;
  assign n36239 = ~n36134 & ~n36238;
  assign n36240 = n36239 ^ n36131;
  assign n36126 = n35734 ^ n35620;
  assign n36122 = n34290 ^ n33387;
  assign n36123 = n35779 ^ n34290;
  assign n36124 = n36122 & ~n36123;
  assign n36125 = n36124 ^ n33387;
  assign n36127 = n36126 ^ n36125;
  assign n36263 = n36240 ^ n36127;
  assign n36363 = n36362 ^ n36263;
  assign n36421 = n36394 ^ n36363;
  assign n36425 = n36424 ^ n36421;
  assign n36426 = n36393 ^ n36364;
  assign n36430 = n36429 ^ n36426;
  assign n36431 = n36392 ^ n36365;
  assign n36432 = n36431 ^ n977;
  assign n36434 = n34174 ^ n25621;
  assign n36435 = n36434 ^ n868;
  assign n36436 = n36435 ^ n964;
  assign n36433 = n36391 ^ n36366;
  assign n36437 = n36436 ^ n36433;
  assign n36438 = n36390 ^ n36388;
  assign n835 = n828 ^ n801;
  assign n854 = n853 ^ n835;
  assign n861 = n860 ^ n854;
  assign n36439 = n36438 ^ n861;
  assign n36441 = n34154 ^ n738;
  assign n36442 = n36441 ^ n30119;
  assign n36443 = n36442 ^ n848;
  assign n36440 = n36387 ^ n36368;
  assign n36444 = n36443 ^ n36440;
  assign n36446 = n34167 ^ n749;
  assign n36447 = n36446 ^ n30137;
  assign n36448 = n36447 ^ n24563;
  assign n36445 = n36386 ^ n36370;
  assign n36449 = n36448 ^ n36445;
  assign n36450 = n36385 ^ n36384;
  assign n36454 = n36453 ^ n36450;
  assign n36456 = n33775 ^ n25738;
  assign n36457 = n36456 ^ n29768;
  assign n36458 = n36457 ^ n24157;
  assign n36455 = n36383 ^ n36381;
  assign n36459 = n36458 ^ n36455;
  assign n36461 = n33634 ^ n25637;
  assign n36462 = n36461 ^ n29762;
  assign n36463 = n36462 ^ n24266;
  assign n36460 = n36380 ^ n36378;
  assign n36464 = n36463 ^ n36460;
  assign n36485 = n36377 ^ n36376;
  assign n36465 = n36375 ^ n36371;
  assign n36469 = n36468 ^ n36465;
  assign n36470 = n36374 ^ n36372;
  assign n36474 = n36473 ^ n36470;
  assign n36059 = n36058 ^ n36057;
  assign n36475 = n36059 ^ n36040;
  assign n35950 = n35949 ^ n35925;
  assign n35954 = n35953 ^ n35950;
  assign n35955 = n35948 ^ n35947;
  assign n2089 = n2085 ^ n2013;
  assign n2096 = n2095 ^ n2089;
  assign n2103 = n2102 ^ n2096;
  assign n35956 = n35955 ^ n2103;
  assign n35957 = n35946 ^ n35927;
  assign n35958 = n35957 ^ n1975;
  assign n35959 = n35945 ^ n35928;
  assign n1934 = n1918 ^ n1873;
  assign n1950 = n1949 ^ n1934;
  assign n1957 = n1956 ^ n1950;
  assign n35960 = n35959 ^ n1957;
  assign n35964 = n35944 ^ n35930;
  assign n35961 = n33662 ^ n1802;
  assign n35962 = n35961 ^ n29656;
  assign n35963 = n35962 ^ n1944;
  assign n35965 = n35964 ^ n35963;
  assign n35967 = n33667 ^ n1790;
  assign n35968 = n35967 ^ n29704;
  assign n35969 = n35968 ^ n24182;
  assign n35966 = n35943 ^ n35931;
  assign n35970 = n35969 ^ n35966;
  assign n35971 = n35942 ^ n35940;
  assign n35975 = n35974 ^ n35971;
  assign n35976 = n35939 ^ n35932;
  assign n35980 = n35979 ^ n35976;
  assign n35982 = n33683 ^ n25651;
  assign n35983 = n35982 ^ n1562;
  assign n35984 = n35983 ^ n24195;
  assign n35981 = n35938 ^ n35934;
  assign n35985 = n35984 ^ n35981;
  assign n35989 = n35937 ^ n35936;
  assign n35986 = n33687 ^ n1529;
  assign n35987 = n35986 ^ n29671;
  assign n35988 = n35987 ^ n25181;
  assign n35990 = n35989 ^ n35988;
  assign n35991 = n33696 ^ n1556;
  assign n35992 = n35991 ^ n29679;
  assign n35993 = n35992 ^ n24199;
  assign n35994 = n35993 ^ n35936;
  assign n35997 = n33691 ^ n2654;
  assign n35998 = n35997 ^ n29674;
  assign n35999 = n35998 ^ n24202;
  assign n35995 = n35875 ^ n32628;
  assign n35996 = n2620 & ~n35995;
  assign n36000 = n35999 ^ n35996;
  assign n36001 = n35879 ^ n35877;
  assign n36002 = n36001 ^ n35999;
  assign n36003 = n36000 & ~n36002;
  assign n36004 = n36003 ^ n35996;
  assign n36005 = n36004 ^ n35936;
  assign n36006 = ~n35994 & n36005;
  assign n36007 = n36006 ^ n35993;
  assign n36008 = n36007 ^ n35989;
  assign n36009 = ~n35990 & n36008;
  assign n36010 = n36009 ^ n35988;
  assign n36011 = n36010 ^ n35981;
  assign n36012 = n35985 & ~n36011;
  assign n36013 = n36012 ^ n35984;
  assign n36014 = n36013 ^ n35976;
  assign n36015 = n35980 & ~n36014;
  assign n36016 = n36015 ^ n35979;
  assign n36017 = n36016 ^ n35971;
  assign n36018 = n35975 & ~n36017;
  assign n36019 = n36018 ^ n35974;
  assign n36020 = n36019 ^ n35966;
  assign n36021 = n35970 & ~n36020;
  assign n36022 = n36021 ^ n35969;
  assign n36023 = n36022 ^ n35964;
  assign n36024 = ~n35965 & n36023;
  assign n36025 = n36024 ^ n35963;
  assign n36026 = n36025 ^ n35959;
  assign n36027 = ~n35960 & n36026;
  assign n36028 = n36027 ^ n1957;
  assign n36029 = n36028 ^ n35957;
  assign n36030 = n35958 & ~n36029;
  assign n36031 = n36030 ^ n1975;
  assign n36032 = n36031 ^ n35955;
  assign n36033 = n35956 & ~n36032;
  assign n36034 = n36033 ^ n2103;
  assign n36035 = n36034 ^ n35950;
  assign n36036 = ~n35954 & n36035;
  assign n36037 = n36036 ^ n35953;
  assign n36476 = n36059 ^ n36037;
  assign n36477 = n36475 & ~n36476;
  assign n36478 = n36477 ^ n36040;
  assign n36479 = n36478 ^ n36470;
  assign n36480 = n36474 & ~n36479;
  assign n36481 = n36480 ^ n36473;
  assign n36482 = n36481 ^ n36465;
  assign n36483 = n36469 & ~n36482;
  assign n36484 = n36483 ^ n36468;
  assign n36486 = n36485 ^ n36484;
  assign n36490 = n36489 ^ n36485;
  assign n36491 = ~n36486 & n36490;
  assign n36492 = n36491 ^ n36489;
  assign n36493 = n36492 ^ n36460;
  assign n36494 = n36464 & ~n36493;
  assign n36495 = n36494 ^ n36463;
  assign n36496 = n36495 ^ n36455;
  assign n36497 = ~n36459 & n36496;
  assign n36498 = n36497 ^ n36458;
  assign n36499 = n36498 ^ n36450;
  assign n36500 = n36454 & ~n36499;
  assign n36501 = n36500 ^ n36453;
  assign n36502 = n36501 ^ n36445;
  assign n36503 = n36449 & ~n36502;
  assign n36504 = n36503 ^ n36448;
  assign n36505 = n36504 ^ n36440;
  assign n36506 = ~n36444 & n36505;
  assign n36507 = n36506 ^ n36443;
  assign n36508 = n36507 ^ n36438;
  assign n36509 = ~n36439 & n36508;
  assign n36510 = n36509 ^ n861;
  assign n36511 = n36510 ^ n36433;
  assign n36512 = ~n36437 & n36511;
  assign n36513 = n36512 ^ n36436;
  assign n36514 = n36513 ^ n36431;
  assign n36515 = n36432 & ~n36514;
  assign n36516 = n36515 ^ n977;
  assign n36517 = n36516 ^ n36426;
  assign n36518 = ~n36430 & n36517;
  assign n36519 = n36518 ^ n36429;
  assign n36520 = n36519 ^ n36421;
  assign n36521 = n36425 & ~n36520;
  assign n36522 = n36521 ^ n36424;
  assign n36417 = n34147 ^ n1396;
  assign n36418 = n36417 ^ n30163;
  assign n36419 = n36418 ^ n1316;
  assign n36575 = n36522 ^ n36419;
  assign n36395 = ~n36363 & n36394;
  assign n36264 = n36263 ^ n32573;
  assign n36334 = n36333 ^ n36263;
  assign n36335 = ~n36264 & n36334;
  assign n36336 = n36335 ^ n32573;
  assign n36241 = n36240 ^ n36126;
  assign n36242 = n36127 & ~n36241;
  assign n36243 = n36242 ^ n36125;
  assign n36117 = n34284 ^ n33385;
  assign n36118 = n34879 ^ n34284;
  assign n36119 = n36117 & ~n36118;
  assign n36120 = n36119 ^ n33385;
  assign n36116 = n35737 ^ n35615;
  assign n36121 = n36120 ^ n36116;
  assign n36261 = n36243 ^ n36121;
  assign n36262 = n36261 ^ n32556;
  assign n36361 = n36336 ^ n36262;
  assign n36416 = n36395 ^ n36361;
  assign n36576 = n36575 ^ n36416;
  assign n36577 = n35281 ^ n33861;
  assign n36578 = n35281 ^ n35142;
  assign n36579 = n36577 & ~n36578;
  assign n36580 = n36579 ^ n33861;
  assign n36581 = n36576 & ~n36580;
  assign n36569 = n35279 ^ n34336;
  assign n36570 = n35827 ^ n35279;
  assign n36571 = n36569 & n36570;
  assign n36572 = n36571 ^ n34336;
  assign n36632 = n36581 ^ n36572;
  assign n36420 = n36419 ^ n36416;
  assign n36523 = n36522 ^ n36416;
  assign n36524 = n36420 & ~n36523;
  assign n36525 = n36524 ^ n36419;
  assign n36412 = n34142 ^ n25775;
  assign n36413 = n36412 ^ n30101;
  assign n36414 = n36413 ^ n24543;
  assign n36396 = ~n36361 & n36395;
  assign n36337 = n36336 ^ n36261;
  assign n36338 = ~n36262 & n36337;
  assign n36339 = n36338 ^ n32556;
  assign n36359 = n36339 ^ n32546;
  assign n36244 = n36243 ^ n36116;
  assign n36245 = n36121 & n36244;
  assign n36246 = n36245 ^ n36120;
  assign n36111 = n34278 ^ n33375;
  assign n36112 = n34915 ^ n34278;
  assign n36113 = n36111 & n36112;
  assign n36114 = n36113 ^ n33375;
  assign n36110 = n35740 ^ n35610;
  assign n36115 = n36114 ^ n36110;
  assign n36259 = n36246 ^ n36115;
  assign n36360 = n36359 ^ n36259;
  assign n36411 = n36396 ^ n36360;
  assign n36415 = n36414 ^ n36411;
  assign n36573 = n36525 ^ n36415;
  assign n36633 = n36632 ^ n36573;
  assign n36629 = n36580 ^ n36576;
  assign n36630 = ~n32756 & ~n36629;
  assign n36631 = n36630 ^ n33426;
  assign n36722 = n36633 ^ n36631;
  assign n36718 = n34767 ^ n25797;
  assign n36719 = n36718 ^ n25010;
  assign n36720 = n36719 ^ n30621;
  assign n36713 = n35028 ^ n26590;
  assign n36714 = n36713 ^ n25336;
  assign n36715 = n36714 ^ n30976;
  assign n36716 = n36629 ^ n32756;
  assign n36717 = n36715 & n36716;
  assign n36721 = n36720 ^ n36717;
  assign n37414 = n36722 ^ n36721;
  assign n37409 = n36054 ^ n35128;
  assign n36775 = n36016 ^ n35975;
  assign n37410 = n36775 ^ n36054;
  assign n37411 = n37409 & ~n37410;
  assign n37412 = n37411 ^ n35128;
  assign n37345 = n36716 ^ n36715;
  assign n37340 = n35922 ^ n35137;
  assign n36069 = n36013 ^ n35979;
  assign n36070 = n36069 ^ n35976;
  assign n37341 = n36070 ^ n35922;
  assign n37342 = n37340 & n37341;
  assign n37343 = n37342 ^ n35137;
  assign n37405 = n37345 ^ n37343;
  assign n37244 = n36516 ^ n36430;
  assign n37095 = n36513 ^ n977;
  assign n37096 = n37095 ^ n36431;
  assign n37090 = n35049 ^ n34265;
  assign n37091 = n35797 ^ n35049;
  assign n37092 = n37090 & n37091;
  assign n37093 = n37092 ^ n34265;
  assign n37240 = n37096 ^ n37093;
  assign n37077 = n36510 ^ n36437;
  assign n37072 = n35006 ^ n34278;
  assign n37073 = n35803 ^ n35006;
  assign n37074 = ~n37072 & ~n37073;
  assign n37075 = n37074 ^ n34278;
  assign n37086 = n37077 ^ n37075;
  assign n37020 = n36507 ^ n861;
  assign n37021 = n37020 ^ n36438;
  assign n37015 = n34960 ^ n34284;
  assign n37016 = n35806 ^ n34960;
  assign n37017 = n37015 & ~n37016;
  assign n37018 = n37017 ^ n34284;
  assign n37068 = n37021 ^ n37018;
  assign n36928 = n36504 ^ n36443;
  assign n36929 = n36928 ^ n36440;
  assign n36924 = n34915 ^ n34290;
  assign n36544 = n35749 ^ n35598;
  assign n36925 = n36544 ^ n34915;
  assign n36926 = n36924 & ~n36925;
  assign n36927 = n36926 ^ n34290;
  assign n36930 = n36929 ^ n36927;
  assign n36794 = n36501 ^ n36448;
  assign n36795 = n36794 ^ n36445;
  assign n36790 = n34879 ^ n34292;
  assign n36355 = n35746 ^ n35600;
  assign n36791 = n36355 ^ n34879;
  assign n36792 = n36790 & n36791;
  assign n36793 = n36792 ^ n34292;
  assign n36796 = n36795 ^ n36793;
  assign n36801 = n36498 ^ n36453;
  assign n36802 = n36801 ^ n36450;
  assign n36797 = n35779 ^ n35039;
  assign n36255 = n35743 ^ n35604;
  assign n36256 = n36255 ^ n35601;
  assign n36798 = n36256 ^ n35779;
  assign n36799 = n36797 & ~n36798;
  assign n36800 = n36799 ^ n35039;
  assign n36803 = n36802 ^ n36800;
  assign n36808 = n36495 ^ n36459;
  assign n36804 = n35514 ^ n34997;
  assign n36805 = n36110 ^ n35514;
  assign n36806 = n36804 & n36805;
  assign n36807 = n36806 ^ n34997;
  assign n36809 = n36808 ^ n36807;
  assign n36811 = n35157 ^ n34955;
  assign n36812 = n36116 ^ n35157;
  assign n36813 = ~n36811 & n36812;
  assign n36814 = n36813 ^ n34955;
  assign n36810 = n36492 ^ n36464;
  assign n36815 = n36814 ^ n36810;
  assign n36817 = n35158 ^ n34905;
  assign n36818 = n36126 ^ n35158;
  assign n36819 = n36817 & n36818;
  assign n36820 = n36819 ^ n34905;
  assign n36816 = n36489 ^ n36486;
  assign n36821 = n36820 ^ n36816;
  assign n36824 = n35165 ^ n34872;
  assign n36825 = n36133 ^ n35165;
  assign n36826 = ~n36824 & n36825;
  assign n36827 = n36826 ^ n34872;
  assign n36822 = n36481 ^ n36468;
  assign n36823 = n36822 ^ n36465;
  assign n36828 = n36827 ^ n36823;
  assign n36833 = n36478 ^ n36474;
  assign n36829 = n35175 ^ n34659;
  assign n36830 = n36140 ^ n35175;
  assign n36831 = n36829 & ~n36830;
  assign n36832 = n36831 ^ n34659;
  assign n36834 = n36833 ^ n36832;
  assign n36835 = n35178 ^ n34585;
  assign n36836 = n36146 ^ n35178;
  assign n36837 = ~n36835 & ~n36836;
  assign n36838 = n36837 ^ n34585;
  assign n36041 = n36040 ^ n36037;
  assign n36060 = n36059 ^ n36041;
  assign n36839 = n36838 ^ n36060;
  assign n36841 = n35185 ^ n34430;
  assign n36842 = n36152 ^ n35185;
  assign n36843 = n36841 & n36842;
  assign n36844 = n36843 ^ n34430;
  assign n36840 = n36034 ^ n35954;
  assign n36845 = n36844 ^ n36840;
  assign n36848 = n35191 ^ n34414;
  assign n36849 = n36220 ^ n35191;
  assign n36850 = n36848 & ~n36849;
  assign n36851 = n36850 ^ n34414;
  assign n36846 = n36031 ^ n2103;
  assign n36847 = n36846 ^ n35955;
  assign n36852 = n36851 ^ n36847;
  assign n36854 = n35197 ^ n33777;
  assign n36855 = n36159 ^ n35197;
  assign n36856 = n36854 & ~n36855;
  assign n36857 = n36856 ^ n33777;
  assign n36853 = n36028 ^ n35958;
  assign n36858 = n36857 ^ n36853;
  assign n36861 = n35203 ^ n33797;
  assign n36862 = n36165 ^ n35203;
  assign n36863 = n36861 & ~n36862;
  assign n36864 = n36863 ^ n33797;
  assign n36859 = n36025 ^ n1957;
  assign n36860 = n36859 ^ n35959;
  assign n36865 = n36864 ^ n36860;
  assign n36867 = n35210 ^ n33804;
  assign n36868 = n36062 ^ n35210;
  assign n36869 = ~n36867 & n36868;
  assign n36870 = n36869 ^ n33804;
  assign n36866 = n36022 ^ n35965;
  assign n36871 = n36870 ^ n36866;
  assign n36876 = n36019 ^ n35969;
  assign n36877 = n36876 ^ n35966;
  assign n36872 = n35220 ^ n33817;
  assign n36873 = n36176 ^ n35220;
  assign n36874 = ~n36872 & n36873;
  assign n36875 = n36874 ^ n33817;
  assign n36878 = n36877 ^ n36875;
  assign n36771 = n35227 ^ n33828;
  assign n36772 = n36183 ^ n35227;
  assign n36773 = ~n36771 & ~n36772;
  assign n36774 = n36773 ^ n33828;
  assign n36776 = n36775 ^ n36774;
  assign n36078 = n36010 ^ n35984;
  assign n36079 = n36078 ^ n35981;
  assign n36072 = n35241 ^ n33841;
  assign n36075 = n36074 ^ n35241;
  assign n36076 = n36072 & n36075;
  assign n36077 = n36076 ^ n33841;
  assign n36080 = n36079 ^ n36077;
  assign n36085 = n36007 ^ n35988;
  assign n36086 = n36085 ^ n35989;
  assign n36081 = n35113 ^ n33848;
  assign n36082 = n36054 ^ n35113;
  assign n36083 = ~n36081 & ~n36082;
  assign n36084 = n36083 ^ n33848;
  assign n36087 = n36086 ^ n36084;
  assign n36089 = n35122 ^ n33859;
  assign n36090 = n35922 ^ n35122;
  assign n36091 = ~n36089 & ~n36090;
  assign n36092 = n36091 ^ n33859;
  assign n36088 = n36004 ^ n35994;
  assign n36093 = n36092 ^ n36088;
  assign n36098 = n36001 ^ n36000;
  assign n36094 = n35128 ^ n34365;
  assign n36095 = n35852 ^ n35128;
  assign n36096 = ~n36094 & ~n36095;
  assign n36097 = n36096 ^ n34365;
  assign n36099 = n36098 ^ n36097;
  assign n36104 = n35995 ^ n2620;
  assign n36100 = n35137 ^ n34359;
  assign n36101 = n35137 ^ n35111;
  assign n36102 = ~n36100 & ~n36101;
  assign n36103 = n36102 ^ n34359;
  assign n36105 = n36104 ^ n36103;
  assign n36250 = n34265 ^ n33371;
  assign n36251 = n34960 ^ n34265;
  assign n36252 = n36250 & n36251;
  assign n36253 = n36252 ^ n33371;
  assign n36351 = n36256 ^ n36253;
  assign n36247 = n36246 ^ n36110;
  assign n36248 = ~n36115 & n36247;
  assign n36249 = n36248 ^ n36114;
  assign n36352 = n36256 ^ n36249;
  assign n36353 = n36351 & n36352;
  assign n36354 = n36353 ^ n36253;
  assign n36356 = n36355 ^ n36354;
  assign n36347 = n33873 ^ n32765;
  assign n36348 = n35006 ^ n33873;
  assign n36349 = n36347 & n36348;
  assign n36350 = n36349 ^ n32765;
  assign n36357 = n36356 ^ n36350;
  assign n36254 = n36253 ^ n36249;
  assign n36257 = n36256 ^ n36254;
  assign n36258 = n36257 ^ n32540;
  assign n36260 = n36259 ^ n32546;
  assign n36340 = n36339 ^ n36259;
  assign n36341 = n36260 & n36340;
  assign n36342 = n36341 ^ n32546;
  assign n36343 = n36342 ^ n36257;
  assign n36344 = ~n36258 & n36343;
  assign n36345 = n36344 ^ n32540;
  assign n36346 = n36345 ^ n31996;
  assign n36358 = n36357 ^ n36346;
  assign n36397 = ~n36360 & ~n36396;
  assign n36398 = n36342 ^ n32540;
  assign n36399 = n36398 ^ n36257;
  assign n36400 = n36397 & ~n36399;
  assign n36552 = n36358 & n36400;
  assign n36545 = n33867 ^ n32763;
  assign n36546 = n35049 ^ n33867;
  assign n36547 = n36545 & n36546;
  assign n36548 = n36547 ^ n32763;
  assign n36549 = n36548 ^ n36544;
  assign n36541 = n36355 ^ n36350;
  assign n36542 = ~n36356 & ~n36541;
  assign n36543 = n36542 ^ n36350;
  assign n36550 = n36549 ^ n36543;
  assign n36536 = n36357 ^ n31996;
  assign n36537 = n36357 ^ n36345;
  assign n36538 = n36536 & n36537;
  assign n36539 = n36538 ^ n31996;
  assign n36540 = n36539 ^ n31990;
  assign n36551 = n36550 ^ n36540;
  assign n36553 = n36552 ^ n36551;
  assign n36402 = n34132 ^ n2446;
  assign n36403 = n36402 ^ n30091;
  assign n36404 = n36403 ^ n2598;
  assign n36401 = n36400 ^ n36358;
  assign n36405 = n36404 ^ n36401;
  assign n36409 = n36399 ^ n36397;
  assign n36406 = n34136 ^ n2457;
  assign n36407 = n36406 ^ n30096;
  assign n36408 = n36407 ^ n24538;
  assign n36410 = n36409 ^ n36408;
  assign n36526 = n36525 ^ n36411;
  assign n36527 = n36415 & ~n36526;
  assign n36528 = n36527 ^ n36414;
  assign n36529 = n36528 ^ n36409;
  assign n36530 = ~n36410 & n36529;
  assign n36531 = n36530 ^ n36408;
  assign n36532 = n36531 ^ n36401;
  assign n36533 = n36405 & ~n36532;
  assign n36534 = n36533 ^ n36404;
  assign n2591 = n2590 ^ n2524;
  assign n2601 = n2600 ^ n2591;
  assign n2602 = n2601 ^ n2576;
  assign n36535 = n36534 ^ n2602;
  assign n36554 = n36553 ^ n36535;
  assign n36106 = n35267 ^ n34343;
  assign n36107 = n35267 ^ n35119;
  assign n36108 = ~n36106 & ~n36107;
  assign n36109 = n36108 ^ n34343;
  assign n36555 = n36554 ^ n36109;
  assign n36560 = n36531 ^ n36405;
  assign n36556 = n35145 ^ n34324;
  assign n36557 = n35145 ^ n35132;
  assign n36558 = ~n36556 & n36557;
  assign n36559 = n36558 ^ n34324;
  assign n36561 = n36560 ^ n36559;
  assign n36566 = n36528 ^ n36408;
  assign n36567 = n36566 ^ n36409;
  assign n36562 = n35152 ^ n34330;
  assign n36563 = n35152 ^ n35134;
  assign n36564 = n36562 & ~n36563;
  assign n36565 = n36564 ^ n34330;
  assign n36568 = n36567 ^ n36565;
  assign n36574 = n36573 ^ n36572;
  assign n36582 = n36581 ^ n36573;
  assign n36583 = ~n36574 & n36582;
  assign n36584 = n36583 ^ n36581;
  assign n36585 = n36584 ^ n36567;
  assign n36586 = n36568 & n36585;
  assign n36587 = n36586 ^ n36565;
  assign n36588 = n36587 ^ n36560;
  assign n36589 = n36561 & n36588;
  assign n36590 = n36589 ^ n36559;
  assign n36591 = n36590 ^ n36554;
  assign n36592 = ~n36555 & n36591;
  assign n36593 = n36592 ^ n36109;
  assign n36594 = n36593 ^ n36104;
  assign n36595 = ~n36105 & n36594;
  assign n36596 = n36595 ^ n36103;
  assign n36597 = n36596 ^ n36098;
  assign n36598 = ~n36099 & ~n36597;
  assign n36599 = n36598 ^ n36097;
  assign n36600 = n36599 ^ n36088;
  assign n36601 = ~n36093 & ~n36600;
  assign n36602 = n36601 ^ n36092;
  assign n36603 = n36602 ^ n36086;
  assign n36604 = n36087 & n36603;
  assign n36605 = n36604 ^ n36084;
  assign n36606 = n36605 ^ n36079;
  assign n36607 = ~n36080 & n36606;
  assign n36608 = n36607 ^ n36077;
  assign n36767 = n36608 ^ n36070;
  assign n36064 = n35234 ^ n34388;
  assign n36066 = n36065 ^ n35234;
  assign n36067 = ~n36064 & ~n36066;
  assign n36068 = n36067 ^ n34388;
  assign n36768 = n36608 ^ n36068;
  assign n36769 = ~n36767 & n36768;
  assign n36770 = n36769 ^ n36070;
  assign n36879 = n36775 ^ n36770;
  assign n36880 = n36776 & ~n36879;
  assign n36881 = n36880 ^ n36774;
  assign n36882 = n36881 ^ n36877;
  assign n36883 = ~n36878 & ~n36882;
  assign n36884 = n36883 ^ n36875;
  assign n36885 = n36884 ^ n36866;
  assign n36886 = n36871 & ~n36885;
  assign n36887 = n36886 ^ n36870;
  assign n36888 = n36887 ^ n36860;
  assign n36889 = ~n36865 & ~n36888;
  assign n36890 = n36889 ^ n36864;
  assign n36891 = n36890 ^ n36853;
  assign n36892 = ~n36858 & ~n36891;
  assign n36893 = n36892 ^ n36857;
  assign n36894 = n36893 ^ n36847;
  assign n36895 = n36852 & n36894;
  assign n36896 = n36895 ^ n36851;
  assign n36897 = n36896 ^ n36840;
  assign n36898 = n36845 & n36897;
  assign n36899 = n36898 ^ n36844;
  assign n36900 = n36899 ^ n36060;
  assign n36901 = ~n36839 & n36900;
  assign n36902 = n36901 ^ n36838;
  assign n36903 = n36902 ^ n36833;
  assign n36904 = n36834 & n36903;
  assign n36905 = n36904 ^ n36832;
  assign n36906 = n36905 ^ n36823;
  assign n36907 = ~n36828 & ~n36906;
  assign n36908 = n36907 ^ n36827;
  assign n36909 = n36908 ^ n36816;
  assign n36910 = ~n36821 & n36909;
  assign n36911 = n36910 ^ n36820;
  assign n36912 = n36911 ^ n36810;
  assign n36913 = ~n36815 & n36912;
  assign n36914 = n36913 ^ n36814;
  assign n36915 = n36914 ^ n36808;
  assign n36916 = n36809 & ~n36915;
  assign n36917 = n36916 ^ n36807;
  assign n36918 = n36917 ^ n36802;
  assign n36919 = n36803 & n36918;
  assign n36920 = n36919 ^ n36800;
  assign n36921 = n36920 ^ n36795;
  assign n36922 = ~n36796 & ~n36921;
  assign n36923 = n36922 ^ n36793;
  assign n37012 = n36929 ^ n36923;
  assign n37013 = ~n36930 & ~n37012;
  assign n37014 = n37013 ^ n36927;
  assign n37069 = n37021 ^ n37014;
  assign n37070 = n37068 & n37069;
  assign n37071 = n37070 ^ n37018;
  assign n37087 = n37077 ^ n37071;
  assign n37088 = n37086 & ~n37087;
  assign n37089 = n37088 ^ n37075;
  assign n37241 = n37096 ^ n37089;
  assign n37242 = n37240 & n37241;
  assign n37243 = n37242 ^ n37093;
  assign n37245 = n37244 ^ n37243;
  assign n37236 = n35104 ^ n33873;
  assign n37237 = n35790 ^ n35104;
  assign n37238 = n37236 & ~n37237;
  assign n37239 = n37238 ^ n33873;
  assign n37246 = n37245 ^ n37239;
  assign n37094 = n37093 ^ n37089;
  assign n37097 = n37096 ^ n37094;
  assign n37231 = n37097 ^ n33371;
  assign n37076 = n37075 ^ n37071;
  assign n37078 = n37077 ^ n37076;
  assign n37081 = n37078 ^ n33375;
  assign n37019 = n37018 ^ n37014;
  assign n37022 = n37021 ^ n37019;
  assign n37023 = n37022 ^ n33385;
  assign n36931 = n36930 ^ n36923;
  assign n36932 = n36931 ^ n33387;
  assign n36933 = n36920 ^ n36796;
  assign n36934 = n36933 ^ n33397;
  assign n36935 = n36917 ^ n36800;
  assign n36936 = n36935 ^ n36802;
  assign n36937 = n36936 ^ n34254;
  assign n36938 = n36911 ^ n36815;
  assign n36939 = n36938 ^ n34003;
  assign n36940 = n36908 ^ n36821;
  assign n36941 = n36940 ^ n33882;
  assign n36942 = n36905 ^ n36828;
  assign n36943 = n36942 ^ n33782;
  assign n36944 = n36902 ^ n36832;
  assign n36945 = n36944 ^ n36833;
  assign n36946 = n36945 ^ n33792;
  assign n36947 = n36899 ^ n36839;
  assign n36948 = n36947 ^ n33799;
  assign n36949 = n36896 ^ n36845;
  assign n36950 = n36949 ^ n33812;
  assign n36951 = n36893 ^ n36852;
  assign n36952 = n36951 ^ n33819;
  assign n36953 = n36890 ^ n36858;
  assign n36954 = n36953 ^ n33940;
  assign n36955 = n36887 ^ n36865;
  assign n36956 = n36955 ^ n33831;
  assign n36957 = n36884 ^ n36871;
  assign n36958 = n36957 ^ n33843;
  assign n36959 = n36881 ^ n36875;
  assign n36960 = n36959 ^ n36877;
  assign n36961 = n36960 ^ n33850;
  assign n36777 = n36776 ^ n36770;
  assign n36778 = n36777 ^ n33908;
  assign n36610 = n36605 ^ n36080;
  assign n36611 = n36610 ^ n33596;
  assign n36612 = n36602 ^ n36084;
  assign n36613 = n36612 ^ n36086;
  assign n36614 = n36613 ^ n33495;
  assign n36615 = n36599 ^ n36093;
  assign n36616 = n36615 ^ n32749;
  assign n36617 = n36596 ^ n36097;
  assign n36618 = n36617 ^ n36098;
  assign n36619 = n36618 ^ n33478;
  assign n36620 = n36593 ^ n36105;
  assign n36621 = n36620 ^ n33472;
  assign n36622 = n36590 ^ n36555;
  assign n36623 = n36622 ^ n33450;
  assign n36624 = n36587 ^ n36559;
  assign n36625 = n36624 ^ n36560;
  assign n36626 = n36625 ^ n33443;
  assign n36627 = n36584 ^ n36568;
  assign n36628 = n36627 ^ n33429;
  assign n36634 = n36633 ^ n36630;
  assign n36635 = n36631 & ~n36634;
  assign n36636 = n36635 ^ n33426;
  assign n36637 = n36636 ^ n36627;
  assign n36638 = ~n36628 & ~n36637;
  assign n36639 = n36638 ^ n33429;
  assign n36640 = n36639 ^ n36625;
  assign n36641 = n36626 & ~n36640;
  assign n36642 = n36641 ^ n33443;
  assign n36643 = n36642 ^ n36622;
  assign n36644 = n36623 & ~n36643;
  assign n36645 = n36644 ^ n33450;
  assign n36646 = n36645 ^ n36620;
  assign n36647 = ~n36621 & ~n36646;
  assign n36648 = n36647 ^ n33472;
  assign n36649 = n36648 ^ n36618;
  assign n36650 = n36619 & n36649;
  assign n36651 = n36650 ^ n33478;
  assign n36652 = n36651 ^ n36615;
  assign n36653 = ~n36616 & n36652;
  assign n36654 = n36653 ^ n32749;
  assign n36655 = n36654 ^ n36613;
  assign n36656 = ~n36614 & n36655;
  assign n36657 = n36656 ^ n33495;
  assign n36658 = n36657 ^ n36610;
  assign n36659 = n36611 & n36658;
  assign n36660 = n36659 ^ n33596;
  assign n36661 = n36660 ^ n33766;
  assign n36071 = n36070 ^ n36068;
  assign n36609 = n36608 ^ n36071;
  assign n36764 = n36660 ^ n36609;
  assign n36765 = ~n36661 & n36764;
  assign n36766 = n36765 ^ n33766;
  assign n36962 = n36777 ^ n36766;
  assign n36963 = n36778 & n36962;
  assign n36964 = n36963 ^ n33908;
  assign n36965 = n36964 ^ n36960;
  assign n36966 = n36961 & n36965;
  assign n36967 = n36966 ^ n33850;
  assign n36968 = n36967 ^ n36957;
  assign n36969 = ~n36958 & ~n36968;
  assign n36970 = n36969 ^ n33843;
  assign n36971 = n36970 ^ n36955;
  assign n36972 = ~n36956 & ~n36971;
  assign n36973 = n36972 ^ n33831;
  assign n36974 = n36973 ^ n36953;
  assign n36975 = n36954 & ~n36974;
  assign n36976 = n36975 ^ n33940;
  assign n36977 = n36976 ^ n36951;
  assign n36978 = n36952 & ~n36977;
  assign n36979 = n36978 ^ n33819;
  assign n36980 = n36979 ^ n36949;
  assign n36981 = ~n36950 & n36980;
  assign n36982 = n36981 ^ n33812;
  assign n36983 = n36982 ^ n36947;
  assign n36984 = n36948 & n36983;
  assign n36985 = n36984 ^ n33799;
  assign n36986 = n36985 ^ n36945;
  assign n36987 = ~n36946 & n36986;
  assign n36988 = n36987 ^ n33792;
  assign n36989 = n36988 ^ n36942;
  assign n36990 = ~n36943 & n36989;
  assign n36991 = n36990 ^ n33782;
  assign n36992 = n36991 ^ n36940;
  assign n36993 = n36941 & ~n36992;
  assign n36994 = n36993 ^ n33882;
  assign n36995 = n36994 ^ n36938;
  assign n36996 = n36939 & ~n36995;
  assign n36997 = n36996 ^ n34003;
  assign n36998 = n36997 ^ n34090;
  assign n36999 = n36914 ^ n36809;
  assign n37000 = n36999 ^ n36997;
  assign n37001 = ~n36998 & n37000;
  assign n37002 = n37001 ^ n34090;
  assign n37003 = n37002 ^ n36936;
  assign n37004 = n36937 & ~n37003;
  assign n37005 = n37004 ^ n34254;
  assign n37006 = n37005 ^ n36933;
  assign n37007 = ~n36934 & ~n37006;
  assign n37008 = n37007 ^ n33397;
  assign n37009 = n37008 ^ n36931;
  assign n37010 = n36932 & ~n37009;
  assign n37011 = n37010 ^ n33387;
  assign n37064 = n37022 ^ n37011;
  assign n37065 = ~n37023 & ~n37064;
  assign n37066 = n37065 ^ n33385;
  assign n37082 = n37078 ^ n37066;
  assign n37083 = n37081 & ~n37082;
  assign n37084 = n37083 ^ n33375;
  assign n37232 = n37097 ^ n37084;
  assign n37233 = ~n37231 & ~n37232;
  assign n37234 = n37233 ^ n33371;
  assign n37235 = n37234 ^ n32765;
  assign n37247 = n37246 ^ n37235;
  assign n37024 = n37023 ^ n37011;
  assign n37025 = n37002 ^ n36937;
  assign n37026 = n36991 ^ n36941;
  assign n37027 = n36988 ^ n33782;
  assign n37028 = n37027 ^ n36942;
  assign n37029 = n36985 ^ n36946;
  assign n37030 = n36982 ^ n33799;
  assign n37031 = n37030 ^ n36947;
  assign n37032 = n36979 ^ n36950;
  assign n37033 = n36964 ^ n33850;
  assign n37034 = n37033 ^ n36960;
  assign n36662 = n36661 ^ n36609;
  assign n36663 = n36636 ^ n33429;
  assign n36664 = n36663 ^ n36627;
  assign n36665 = n36639 ^ n36626;
  assign n36666 = n36664 & n36665;
  assign n36667 = n36642 ^ n33450;
  assign n36668 = n36667 ^ n36622;
  assign n36669 = n36666 & n36668;
  assign n36670 = n36645 ^ n36621;
  assign n36671 = ~n36669 & n36670;
  assign n36672 = n36648 ^ n33478;
  assign n36673 = n36672 ^ n36618;
  assign n36674 = ~n36671 & ~n36673;
  assign n36675 = n36651 ^ n36616;
  assign n36676 = n36674 & ~n36675;
  assign n36677 = n36654 ^ n33495;
  assign n36678 = n36677 ^ n36613;
  assign n36679 = ~n36676 & n36678;
  assign n36680 = n36657 ^ n36611;
  assign n36681 = n36679 & ~n36680;
  assign n36763 = ~n36662 & ~n36681;
  assign n36779 = n36778 ^ n36766;
  assign n37035 = n36763 & n36779;
  assign n37036 = ~n37034 & n37035;
  assign n37037 = n36967 ^ n36958;
  assign n37038 = n37036 & ~n37037;
  assign n37039 = n36970 ^ n33831;
  assign n37040 = n37039 ^ n36955;
  assign n37041 = ~n37038 & ~n37040;
  assign n37042 = n36973 ^ n36954;
  assign n37043 = ~n37041 & n37042;
  assign n37044 = n36976 ^ n36952;
  assign n37045 = n37043 & n37044;
  assign n37046 = ~n37032 & n37045;
  assign n37047 = ~n37031 & ~n37046;
  assign n37048 = n37029 & ~n37047;
  assign n37049 = n37028 & n37048;
  assign n37050 = n37026 & ~n37049;
  assign n37051 = n36994 ^ n34003;
  assign n37052 = n37051 ^ n36938;
  assign n37053 = n37050 & n37052;
  assign n37054 = n36999 ^ n34090;
  assign n37055 = n37054 ^ n36997;
  assign n37056 = n37053 & n37055;
  assign n37057 = n37025 & ~n37056;
  assign n37058 = n37005 ^ n36934;
  assign n37059 = n37057 & ~n37058;
  assign n37060 = n37008 ^ n33387;
  assign n37061 = n37060 ^ n36931;
  assign n37062 = n37059 & ~n37061;
  assign n37063 = n37024 & n37062;
  assign n37067 = n37066 ^ n33375;
  assign n37079 = n37078 ^ n37067;
  assign n37080 = ~n37063 & ~n37079;
  assign n37085 = n37084 ^ n33371;
  assign n37098 = n37097 ^ n37085;
  assign n37248 = n37080 & n37098;
  assign n37310 = ~n37247 & n37248;
  assign n37307 = n36519 ^ n36425;
  assign n37302 = n35287 ^ n33867;
  assign n37303 = n35784 ^ n35287;
  assign n37304 = ~n37302 & n37303;
  assign n37305 = n37304 ^ n33867;
  assign n37299 = n37244 ^ n37239;
  assign n37300 = n37245 & n37299;
  assign n37301 = n37300 ^ n37239;
  assign n37306 = n37305 ^ n37301;
  assign n37308 = n37307 ^ n37306;
  assign n37294 = n37246 ^ n32765;
  assign n37295 = n37246 ^ n37234;
  assign n37296 = ~n37294 & ~n37295;
  assign n37297 = n37296 ^ n32765;
  assign n37298 = n37297 ^ n32763;
  assign n37309 = n37308 ^ n37298;
  assign n37311 = n37310 ^ n37309;
  assign n37290 = n35004 ^ n26569;
  assign n37291 = n37290 ^ n2492;
  assign n37292 = n37291 ^ n30939;
  assign n37250 = n34939 ^ n26480;
  assign n37251 = n37250 ^ n25211;
  assign n37252 = n37251 ^ n2369;
  assign n37249 = n37248 ^ n37247;
  assign n37253 = n37252 ^ n37249;
  assign n37100 = n34913 ^ n26543;
  assign n37101 = n37100 ^ n30805;
  assign n37102 = n37101 ^ n2357;
  assign n37099 = n37098 ^ n37080;
  assign n37103 = n37102 ^ n37099;
  assign n37223 = n37079 ^ n37063;
  assign n37105 = n34667 ^ n26487;
  assign n37106 = n37105 ^ n1252;
  assign n37107 = n37106 ^ n2300;
  assign n37104 = n37062 ^ n37024;
  assign n37108 = n37107 ^ n37104;
  assign n37109 = n37061 ^ n37059;
  assign n1231 = n1224 ^ n1146;
  assign n1238 = n1237 ^ n1231;
  assign n1245 = n1244 ^ n1238;
  assign n37110 = n37109 ^ n1245;
  assign n37111 = n37058 ^ n37057;
  assign n1100 = n1056 ^ n1021;
  assign n1107 = n1106 ^ n1100;
  assign n1108 = n1107 ^ n1097;
  assign n37112 = n37111 ^ n1108;
  assign n37113 = n37056 ^ n37025;
  assign n1067 = n1061 ^ n1003;
  assign n1077 = n1076 ^ n1067;
  assign n1090 = n1089 ^ n1077;
  assign n37114 = n37113 ^ n1090;
  assign n37115 = n37055 ^ n37053;
  assign n37119 = n37118 ^ n37115;
  assign n37121 = n34683 ^ n930;
  assign n37122 = n37121 ^ n30693;
  assign n37123 = n37122 ^ n25094;
  assign n37120 = n37052 ^ n37050;
  assign n37124 = n37123 ^ n37120;
  assign n37128 = n37049 ^ n37026;
  assign n37129 = n37128 ^ n37127;
  assign n37133 = n37048 ^ n37028;
  assign n37130 = n34692 ^ n26505;
  assign n37131 = n37130 ^ n30717;
  assign n37132 = n37131 ^ n569;
  assign n37134 = n37133 ^ n37132;
  assign n37138 = n37047 ^ n37029;
  assign n37135 = n34697 ^ n25808;
  assign n37136 = n37135 ^ n662;
  assign n37137 = n37136 ^ n25080;
  assign n37139 = n37138 ^ n37137;
  assign n37143 = n37046 ^ n37031;
  assign n37140 = n34703 ^ n26243;
  assign n37141 = n37140 ^ n30712;
  assign n37142 = n37141 ^ n657;
  assign n37144 = n37143 ^ n37142;
  assign n37145 = n37045 ^ n37032;
  assign n37149 = n37148 ^ n37145;
  assign n37182 = n37044 ^ n37043;
  assign n37150 = n37042 ^ n37041;
  assign n37154 = n37153 ^ n37150;
  assign n37171 = n37040 ^ n37038;
  assign n37158 = n37037 ^ n37036;
  assign n37155 = n34722 ^ n26203;
  assign n37156 = n37155 ^ n24985;
  assign n37157 = n37156 ^ n2262;
  assign n37159 = n37158 ^ n37157;
  assign n37163 = n37035 ^ n37034;
  assign n36780 = n36779 ^ n36763;
  assign n2220 = n2132 ^ n2064;
  assign n2230 = n2229 ^ n2220;
  assign n2237 = n2236 ^ n2230;
  assign n36781 = n36780 ^ n2237;
  assign n36683 = n34732 ^ n2046;
  assign n36684 = n36683 ^ n30594;
  assign n36685 = n36684 ^ n2226;
  assign n36682 = n36681 ^ n36662;
  assign n36686 = n36685 ^ n36682;
  assign n36687 = n36680 ^ n36679;
  assign n36691 = n36690 ^ n36687;
  assign n36749 = n36678 ^ n36676;
  assign n36695 = n36675 ^ n36674;
  assign n36692 = n34746 ^ n26142;
  assign n36693 = n36692 ^ n30608;
  assign n36694 = n36693 ^ n1704;
  assign n36696 = n36695 ^ n36694;
  assign n36697 = n36673 ^ n36671;
  assign n1620 = n1619 ^ n1592;
  assign n1630 = n1629 ^ n1620;
  assign n1637 = n1636 ^ n1630;
  assign n36698 = n36697 ^ n1637;
  assign n36702 = n36670 ^ n36669;
  assign n36699 = n34753 ^ n26149;
  assign n36700 = n36699 ^ n30613;
  assign n36701 = n36700 ^ n1614;
  assign n36703 = n36702 ^ n36701;
  assign n36707 = n36668 ^ n36666;
  assign n36708 = n36707 ^ n36706;
  assign n36729 = n36665 ^ n36664;
  assign n36712 = n36711 ^ n36664;
  assign n36723 = n36722 ^ n36720;
  assign n36724 = n36721 & ~n36723;
  assign n36725 = n36724 ^ n36717;
  assign n36726 = n36725 ^ n36664;
  assign n36727 = n36712 & ~n36726;
  assign n36728 = n36727 ^ n36711;
  assign n36730 = n36729 ^ n36728;
  assign n36731 = n34763 ^ n26164;
  assign n36732 = n36731 ^ n25005;
  assign n36733 = n36732 ^ n30634;
  assign n36734 = n36733 ^ n36729;
  assign n36735 = n36730 & ~n36734;
  assign n36736 = n36735 ^ n36733;
  assign n36737 = n36736 ^ n36707;
  assign n36738 = ~n36708 & n36737;
  assign n36739 = n36738 ^ n36706;
  assign n36740 = n36739 ^ n36702;
  assign n36741 = ~n36703 & n36740;
  assign n36742 = n36741 ^ n36701;
  assign n36743 = n36742 ^ n36697;
  assign n36744 = ~n36698 & n36743;
  assign n36745 = n36744 ^ n1637;
  assign n36746 = n36745 ^ n36695;
  assign n36747 = n36696 & ~n36746;
  assign n36748 = n36747 ^ n36694;
  assign n36750 = n36749 ^ n36748;
  assign n36751 = n34742 ^ n26137;
  assign n36752 = n36751 ^ n1709;
  assign n36753 = n36752 ^ n24994;
  assign n36754 = n36753 ^ n36749;
  assign n36755 = n36750 & ~n36754;
  assign n36756 = n36755 ^ n36753;
  assign n36757 = n36756 ^ n36687;
  assign n36758 = ~n36691 & n36757;
  assign n36759 = n36758 ^ n36690;
  assign n36760 = n36759 ^ n36682;
  assign n36761 = ~n36686 & n36760;
  assign n36762 = n36761 ^ n36685;
  assign n37160 = n36780 ^ n36762;
  assign n37161 = ~n36781 & n37160;
  assign n37162 = n37161 ^ n2237;
  assign n37164 = n37163 ^ n37162;
  assign n37165 = n37163 ^ n2252;
  assign n37166 = ~n37164 & n37165;
  assign n37167 = n37166 ^ n2252;
  assign n37168 = n37167 ^ n37158;
  assign n37169 = n37159 & ~n37168;
  assign n37170 = n37169 ^ n37157;
  assign n37172 = n37171 ^ n37170;
  assign n37176 = n37175 ^ n37171;
  assign n37177 = ~n37172 & n37176;
  assign n37178 = n37177 ^ n37175;
  assign n37179 = n37178 ^ n37150;
  assign n37180 = n37154 & ~n37179;
  assign n37181 = n37180 ^ n37153;
  assign n37183 = n37182 ^ n37181;
  assign n37184 = n34708 ^ n26217;
  assign n37185 = n37184 ^ n30568;
  assign n37186 = n37185 ^ n24970;
  assign n37187 = n37186 ^ n37182;
  assign n37188 = n37183 & ~n37187;
  assign n37189 = n37188 ^ n37186;
  assign n37190 = n37189 ^ n37145;
  assign n37191 = n37149 & ~n37190;
  assign n37192 = n37191 ^ n37148;
  assign n37193 = n37192 ^ n37142;
  assign n37194 = n37144 & ~n37193;
  assign n37195 = n37194 ^ n37143;
  assign n37196 = n37195 ^ n37138;
  assign n37197 = n37139 & ~n37196;
  assign n37198 = n37197 ^ n37137;
  assign n37199 = n37198 ^ n37133;
  assign n37200 = ~n37134 & n37199;
  assign n37201 = n37200 ^ n37132;
  assign n37202 = n37201 ^ n37128;
  assign n37203 = ~n37129 & n37202;
  assign n37204 = n37203 ^ n37127;
  assign n37205 = n37204 ^ n37120;
  assign n37206 = n37124 & ~n37205;
  assign n37207 = n37206 ^ n37123;
  assign n37208 = n37207 ^ n37115;
  assign n37209 = n37119 & ~n37208;
  assign n37210 = n37209 ^ n37118;
  assign n37211 = n37210 ^ n37113;
  assign n37212 = n37114 & ~n37211;
  assign n37213 = n37212 ^ n1090;
  assign n37214 = n37213 ^ n37111;
  assign n37215 = n37112 & ~n37214;
  assign n37216 = n37215 ^ n1108;
  assign n37217 = n37216 ^ n37109;
  assign n37218 = n37110 & ~n37217;
  assign n37219 = n37218 ^ n1245;
  assign n37220 = n37219 ^ n37104;
  assign n37221 = ~n37108 & n37220;
  assign n37222 = n37221 ^ n37107;
  assign n37224 = n37223 ^ n37222;
  assign n2283 = n2282 ^ n1337;
  assign n2296 = n2295 ^ n2283;
  assign n2303 = n2302 ^ n2296;
  assign n37225 = n37223 ^ n2303;
  assign n37226 = ~n37224 & n37225;
  assign n37227 = n37226 ^ n2303;
  assign n37228 = n37227 ^ n37099;
  assign n37229 = n37103 & ~n37228;
  assign n37230 = n37229 ^ n37102;
  assign n37287 = n37249 ^ n37230;
  assign n37288 = ~n37253 & n37287;
  assign n37289 = n37288 ^ n37252;
  assign n37293 = n37292 ^ n37289;
  assign n37312 = n37311 ^ n37293;
  assign n37283 = n35852 ^ n35267;
  assign n37284 = n36079 ^ n35852;
  assign n37285 = ~n37283 & ~n37284;
  assign n37286 = n37285 ^ n35267;
  assign n37313 = n37312 ^ n37286;
  assign n37254 = n37253 ^ n37230;
  assign n36786 = n35145 ^ n35111;
  assign n36787 = n36086 ^ n35111;
  assign n36788 = n36786 & ~n36787;
  assign n36789 = n36788 ^ n35145;
  assign n37255 = n37254 ^ n36789;
  assign n37260 = n37227 ^ n37103;
  assign n37256 = n35152 ^ n35119;
  assign n37257 = n36088 ^ n35119;
  assign n37258 = n37256 & ~n37257;
  assign n37259 = n37258 ^ n35152;
  assign n37261 = n37260 ^ n37259;
  assign n37266 = n37219 ^ n37108;
  assign n37267 = n35281 ^ n35134;
  assign n37268 = n36104 ^ n35134;
  assign n37269 = n37267 & ~n37268;
  assign n37270 = n37269 ^ n35281;
  assign n37271 = ~n37266 & ~n37270;
  assign n37262 = n35279 ^ n35132;
  assign n37263 = n36098 ^ n35132;
  assign n37264 = n37262 & ~n37263;
  assign n37265 = n37264 ^ n35279;
  assign n37272 = n37271 ^ n37265;
  assign n37273 = n37224 ^ n2303;
  assign n37274 = n37273 ^ n37265;
  assign n37275 = n37272 & ~n37274;
  assign n37276 = n37275 ^ n37271;
  assign n37277 = n37276 ^ n37260;
  assign n37278 = ~n37261 & ~n37277;
  assign n37279 = n37278 ^ n37259;
  assign n37280 = n37279 ^ n37254;
  assign n37281 = n37255 & ~n37280;
  assign n37282 = n37281 ^ n36789;
  assign n37337 = n37312 ^ n37282;
  assign n37338 = n37313 & ~n37337;
  assign n37339 = n37338 ^ n37286;
  assign n37406 = n37345 ^ n37339;
  assign n37407 = ~n37405 & n37406;
  assign n37408 = n37407 ^ n37343;
  assign n37413 = n37412 ^ n37408;
  assign n37415 = n37414 ^ n37413;
  assign n37344 = n37343 ^ n37339;
  assign n37346 = n37345 ^ n37344;
  assign n37347 = n37346 ^ n34359;
  assign n37314 = n37313 ^ n37282;
  assign n37315 = n37314 ^ n34343;
  assign n37316 = n37279 ^ n36789;
  assign n37317 = n37316 ^ n37254;
  assign n37318 = n37317 ^ n34324;
  assign n37319 = n37276 ^ n37261;
  assign n37320 = n37319 ^ n34330;
  assign n37321 = n37270 ^ n37266;
  assign n37322 = ~n33861 & n37321;
  assign n37323 = n37322 ^ n34336;
  assign n37324 = n37273 ^ n37272;
  assign n37325 = n37324 ^ n37322;
  assign n37326 = n37323 & ~n37325;
  assign n37327 = n37326 ^ n34336;
  assign n37328 = n37327 ^ n37319;
  assign n37329 = n37320 & n37328;
  assign n37330 = n37329 ^ n34330;
  assign n37331 = n37330 ^ n37317;
  assign n37332 = ~n37318 & ~n37331;
  assign n37333 = n37332 ^ n34324;
  assign n37334 = n37333 ^ n37314;
  assign n37335 = ~n37315 & n37334;
  assign n37336 = n37335 ^ n34343;
  assign n37401 = n37346 ^ n37336;
  assign n37402 = n37347 & ~n37401;
  assign n37403 = n37402 ^ n34359;
  assign n37404 = n37403 ^ n34365;
  assign n37416 = n37415 ^ n37404;
  assign n37348 = n37347 ^ n37336;
  assign n37349 = n37333 ^ n34343;
  assign n37350 = n37349 ^ n37314;
  assign n37351 = n37330 ^ n37318;
  assign n37352 = n37327 ^ n34330;
  assign n37353 = n37352 ^ n37319;
  assign n37354 = ~n37351 & ~n37353;
  assign n37355 = n37350 & n37354;
  assign n37400 = n37348 & ~n37355;
  assign n37417 = n37416 ^ n37400;
  assign n37418 = n37417 ^ n37399;
  assign n37356 = n37355 ^ n37348;
  assign n37360 = n37359 ^ n37356;
  assign n37361 = n37354 ^ n37350;
  assign n37365 = n37364 ^ n37361;
  assign n37367 = n35065 ^ n26963;
  assign n37368 = n37367 ^ n30865;
  assign n37369 = n37368 ^ n25181;
  assign n37366 = n37353 ^ n37351;
  assign n37370 = n37369 ^ n37366;
  assign n37371 = n35069 ^ n26971;
  assign n37372 = n37371 ^ n30874;
  assign n37373 = n37372 ^ n1556;
  assign n37374 = n37373 ^ n37353;
  assign n37377 = n35072 ^ n26967;
  assign n37378 = n37377 ^ n2654;
  assign n37379 = n37378 ^ n30869;
  assign n2571 = n2570 ^ n2501;
  assign n2572 = n2571 ^ n2555;
  assign n2579 = n2578 ^ n2572;
  assign n37375 = n37321 ^ n33861;
  assign n37376 = n2579 & ~n37375;
  assign n37380 = n37379 ^ n37376;
  assign n37381 = n37324 ^ n37323;
  assign n37382 = n37381 ^ n37379;
  assign n37383 = n37380 & ~n37382;
  assign n37384 = n37383 ^ n37376;
  assign n37385 = n37384 ^ n37353;
  assign n37386 = ~n37374 & n37385;
  assign n37387 = n37386 ^ n37373;
  assign n37388 = n37387 ^ n37369;
  assign n37389 = ~n37370 & ~n37388;
  assign n37390 = n37389 ^ n37366;
  assign n37391 = n37390 ^ n37361;
  assign n37392 = ~n37365 & ~n37391;
  assign n37393 = n37392 ^ n37364;
  assign n37394 = n37393 ^ n37356;
  assign n37395 = ~n37360 & n37394;
  assign n37396 = n37395 ^ n37359;
  assign n37952 = n37417 ^ n37396;
  assign n37953 = ~n37418 & n37952;
  assign n37954 = n37953 ^ n37399;
  assign n37827 = ~n37400 & ~n37416;
  assign n37724 = n37415 ^ n34365;
  assign n37725 = n37415 ^ n37403;
  assign n37726 = n37724 & n37725;
  assign n37727 = n37726 ^ n34365;
  assign n37825 = n37727 ^ n33859;
  assign n37592 = n37414 ^ n37412;
  assign n37593 = n37414 ^ n37408;
  assign n37594 = n37592 & n37593;
  assign n37595 = n37594 ^ n37412;
  assign n37587 = n36074 ^ n35122;
  assign n37588 = n36877 ^ n36074;
  assign n37589 = ~n37587 & ~n37588;
  assign n37590 = n37589 ^ n35122;
  assign n37721 = n37595 ^ n37590;
  assign n37586 = n36725 ^ n36712;
  assign n37722 = n37721 ^ n37586;
  assign n37826 = n37825 ^ n37722;
  assign n37950 = n37827 ^ n37826;
  assign n37947 = n35684 ^ n1684;
  assign n37948 = n37947 ^ n31229;
  assign n37949 = n37948 ^ n1790;
  assign n37951 = n37950 ^ n37949;
  assign n38131 = n37954 ^ n37951;
  assign n37444 = n36745 ^ n36696;
  assign n39429 = n38131 ^ n37444;
  assign n38087 = n36088 ^ n35134;
  assign n38088 = n37345 ^ n36088;
  assign n38089 = n38087 & n38088;
  assign n38090 = n38089 ^ n35134;
  assign n37504 = n36355 ^ n35514;
  assign n37505 = n37077 ^ n36355;
  assign n37506 = ~n37504 & n37505;
  assign n37507 = n37506 ^ n35514;
  assign n37503 = n37192 ^ n37144;
  assign n37508 = n37507 ^ n37503;
  assign n37511 = n36110 ^ n35158;
  assign n37512 = n36929 ^ n36110;
  assign n37513 = ~n37511 & n37512;
  assign n37514 = n37513 ^ n35158;
  assign n37510 = n37186 ^ n37183;
  assign n37515 = n37514 ^ n37510;
  assign n37517 = n36116 ^ n35165;
  assign n37518 = n36795 ^ n36116;
  assign n37519 = ~n37517 & n37518;
  assign n37520 = n37519 ^ n35165;
  assign n37516 = n37178 ^ n37154;
  assign n37521 = n37520 ^ n37516;
  assign n37526 = n37175 ^ n37172;
  assign n37522 = n36126 ^ n35175;
  assign n37523 = n36802 ^ n36126;
  assign n37524 = n37522 & ~n37523;
  assign n37525 = n37524 ^ n35175;
  assign n37527 = n37526 ^ n37525;
  assign n37532 = n37167 ^ n37159;
  assign n37528 = n36133 ^ n35178;
  assign n37529 = n36808 ^ n36133;
  assign n37530 = ~n37528 & ~n37529;
  assign n37531 = n37530 ^ n35178;
  assign n37533 = n37532 ^ n37531;
  assign n37538 = n37164 ^ n2252;
  assign n37534 = n36140 ^ n35185;
  assign n37535 = n36810 ^ n36140;
  assign n37536 = ~n37534 & ~n37535;
  assign n37537 = n37536 ^ n35185;
  assign n37539 = n37538 ^ n37537;
  assign n37540 = n36146 ^ n35191;
  assign n37541 = n36816 ^ n36146;
  assign n37542 = n37540 & ~n37541;
  assign n37543 = n37542 ^ n35191;
  assign n36782 = n36781 ^ n36762;
  assign n37544 = n37543 ^ n36782;
  assign n37545 = n36152 ^ n35197;
  assign n37546 = n36823 ^ n36152;
  assign n37547 = ~n37545 & ~n37546;
  assign n37548 = n37547 ^ n35197;
  assign n37422 = n36759 ^ n36686;
  assign n37549 = n37548 ^ n37422;
  assign n37550 = n36220 ^ n35203;
  assign n37551 = n36833 ^ n36220;
  assign n37552 = n37550 & ~n37551;
  assign n37553 = n37552 ^ n35203;
  assign n37430 = n36756 ^ n36691;
  assign n37554 = n37553 ^ n37430;
  assign n37555 = n36159 ^ n35210;
  assign n37556 = n36159 ^ n36060;
  assign n37557 = ~n37555 & n37556;
  assign n37558 = n37557 ^ n35210;
  assign n37437 = n36753 ^ n36750;
  assign n37559 = n37558 ^ n37437;
  assign n37560 = n36165 ^ n35220;
  assign n37561 = n36840 ^ n36165;
  assign n37562 = n37560 & n37561;
  assign n37563 = n37562 ^ n35220;
  assign n37564 = n37563 ^ n37444;
  assign n37565 = n36062 ^ n35227;
  assign n37566 = n36847 ^ n36062;
  assign n37567 = n37565 & n37566;
  assign n37568 = n37567 ^ n35227;
  assign n37451 = n36742 ^ n36698;
  assign n37569 = n37568 ^ n37451;
  assign n37570 = n36176 ^ n35234;
  assign n37571 = n36853 ^ n36176;
  assign n37572 = n37570 & n37571;
  assign n37573 = n37572 ^ n35234;
  assign n37458 = n36739 ^ n36703;
  assign n37574 = n37573 ^ n37458;
  assign n37575 = n36183 ^ n35241;
  assign n37576 = n36860 ^ n36183;
  assign n37577 = n37575 & ~n37576;
  assign n37578 = n37577 ^ n35241;
  assign n37464 = n36736 ^ n36708;
  assign n37579 = n37578 ^ n37464;
  assign n37581 = n36065 ^ n35113;
  assign n37582 = n36866 ^ n36065;
  assign n37583 = ~n37581 & ~n37582;
  assign n37584 = n37583 ^ n35113;
  assign n37580 = n36733 ^ n36730;
  assign n37585 = n37584 ^ n37580;
  assign n37591 = n37590 ^ n37586;
  assign n37596 = n37595 ^ n37586;
  assign n37597 = ~n37591 & ~n37596;
  assign n37598 = n37597 ^ n37590;
  assign n37599 = n37598 ^ n37580;
  assign n37600 = ~n37585 & ~n37599;
  assign n37601 = n37600 ^ n37584;
  assign n37602 = n37601 ^ n37464;
  assign n37603 = n37579 & n37602;
  assign n37604 = n37603 ^ n37578;
  assign n37605 = n37604 ^ n37458;
  assign n37606 = n37574 & ~n37605;
  assign n37607 = n37606 ^ n37573;
  assign n37608 = n37607 ^ n37451;
  assign n37609 = n37569 & ~n37608;
  assign n37610 = n37609 ^ n37568;
  assign n37611 = n37610 ^ n37444;
  assign n37612 = n37564 & n37611;
  assign n37613 = n37612 ^ n37563;
  assign n37614 = n37613 ^ n37437;
  assign n37615 = ~n37559 & n37614;
  assign n37616 = n37615 ^ n37558;
  assign n37617 = n37616 ^ n37430;
  assign n37618 = ~n37554 & n37617;
  assign n37619 = n37618 ^ n37553;
  assign n37620 = n37619 ^ n37422;
  assign n37621 = n37549 & n37620;
  assign n37622 = n37621 ^ n37548;
  assign n37623 = n37622 ^ n36782;
  assign n37624 = ~n37544 & ~n37623;
  assign n37625 = n37624 ^ n37543;
  assign n37626 = n37625 ^ n37538;
  assign n37627 = ~n37539 & ~n37626;
  assign n37628 = n37627 ^ n37537;
  assign n37629 = n37628 ^ n37532;
  assign n37630 = n37533 & n37629;
  assign n37631 = n37630 ^ n37531;
  assign n37632 = n37631 ^ n37526;
  assign n37633 = n37527 & ~n37632;
  assign n37634 = n37633 ^ n37525;
  assign n37635 = n37634 ^ n37516;
  assign n37636 = n37521 & ~n37635;
  assign n37637 = n37636 ^ n37520;
  assign n37638 = n37637 ^ n37510;
  assign n37639 = n37515 & n37638;
  assign n37640 = n37639 ^ n37514;
  assign n37509 = n37189 ^ n37149;
  assign n37641 = n37640 ^ n37509;
  assign n37642 = n36256 ^ n35157;
  assign n37643 = n37021 ^ n36256;
  assign n37644 = n37642 & n37643;
  assign n37645 = n37644 ^ n35157;
  assign n37646 = n37645 ^ n37509;
  assign n37647 = n37641 & n37646;
  assign n37648 = n37647 ^ n37645;
  assign n37649 = n37648 ^ n37503;
  assign n37650 = ~n37508 & ~n37649;
  assign n37651 = n37650 ^ n37507;
  assign n37498 = n36544 ^ n35779;
  assign n37499 = n37096 ^ n36544;
  assign n37500 = n37498 & ~n37499;
  assign n37501 = n37500 ^ n35779;
  assign n37682 = n37651 ^ n37501;
  assign n37497 = n37195 ^ n37139;
  assign n37683 = n37682 ^ n37497;
  assign n37684 = n37683 ^ n35039;
  assign n37685 = n37648 ^ n37507;
  assign n37686 = n37685 ^ n37503;
  assign n37687 = n37686 ^ n34997;
  assign n37688 = n37645 ^ n37641;
  assign n37689 = n37688 ^ n34955;
  assign n37690 = n37637 ^ n37514;
  assign n37691 = n37690 ^ n37510;
  assign n37692 = n37691 ^ n34905;
  assign n37693 = n37634 ^ n37521;
  assign n37694 = n37693 ^ n34872;
  assign n37695 = n37631 ^ n37527;
  assign n37696 = n37695 ^ n34659;
  assign n37697 = n37628 ^ n37533;
  assign n37698 = n37697 ^ n34585;
  assign n37699 = n37625 ^ n37539;
  assign n37700 = n37699 ^ n34430;
  assign n37701 = n37622 ^ n37544;
  assign n37702 = n37701 ^ n34414;
  assign n37703 = n37619 ^ n37549;
  assign n37704 = n37703 ^ n33777;
  assign n37749 = n37616 ^ n37554;
  assign n37705 = n37613 ^ n37559;
  assign n37706 = n37705 ^ n33804;
  assign n37707 = n37610 ^ n37563;
  assign n37708 = n37707 ^ n37444;
  assign n37709 = n37708 ^ n33817;
  assign n37710 = n37607 ^ n37569;
  assign n37711 = n37710 ^ n33828;
  assign n37712 = n37604 ^ n37573;
  assign n37713 = n37712 ^ n37458;
  assign n37714 = n37713 ^ n34388;
  assign n37715 = n37601 ^ n37578;
  assign n37716 = n37715 ^ n37464;
  assign n37717 = n37716 ^ n33841;
  assign n37718 = n37598 ^ n37584;
  assign n37719 = n37718 ^ n37580;
  assign n37720 = n37719 ^ n33848;
  assign n37723 = n37722 ^ n33859;
  assign n37728 = n37727 ^ n37722;
  assign n37729 = ~n37723 & ~n37728;
  assign n37730 = n37729 ^ n33859;
  assign n37731 = n37730 ^ n37719;
  assign n37732 = ~n37720 & ~n37731;
  assign n37733 = n37732 ^ n33848;
  assign n37734 = n37733 ^ n37716;
  assign n37735 = ~n37717 & n37734;
  assign n37736 = n37735 ^ n33841;
  assign n37737 = n37736 ^ n37713;
  assign n37738 = ~n37714 & ~n37737;
  assign n37739 = n37738 ^ n34388;
  assign n37740 = n37739 ^ n37710;
  assign n37741 = ~n37711 & n37740;
  assign n37742 = n37741 ^ n33828;
  assign n37743 = n37742 ^ n37708;
  assign n37744 = n37709 & n37743;
  assign n37745 = n37744 ^ n33817;
  assign n37746 = n37745 ^ n37705;
  assign n37747 = n37706 & ~n37746;
  assign n37748 = n37747 ^ n33804;
  assign n37750 = n37749 ^ n37748;
  assign n37751 = n37749 ^ n33797;
  assign n37752 = ~n37750 & ~n37751;
  assign n37753 = n37752 ^ n33797;
  assign n37754 = n37753 ^ n37703;
  assign n37755 = ~n37704 & ~n37754;
  assign n37756 = n37755 ^ n33777;
  assign n37757 = n37756 ^ n37701;
  assign n37758 = n37702 & n37757;
  assign n37759 = n37758 ^ n34414;
  assign n37760 = n37759 ^ n37699;
  assign n37761 = n37700 & n37760;
  assign n37762 = n37761 ^ n34430;
  assign n37763 = n37762 ^ n37697;
  assign n37764 = n37698 & ~n37763;
  assign n37765 = n37764 ^ n34585;
  assign n37766 = n37765 ^ n37695;
  assign n37767 = n37696 & n37766;
  assign n37768 = n37767 ^ n34659;
  assign n37769 = n37768 ^ n37693;
  assign n37770 = ~n37694 & ~n37769;
  assign n37771 = n37770 ^ n34872;
  assign n37772 = n37771 ^ n37691;
  assign n37773 = ~n37692 & n37772;
  assign n37774 = n37773 ^ n34905;
  assign n37775 = n37774 ^ n37688;
  assign n37776 = n37689 & ~n37775;
  assign n37777 = n37776 ^ n34955;
  assign n37778 = n37777 ^ n37686;
  assign n37779 = n37687 & ~n37778;
  assign n37780 = n37779 ^ n34997;
  assign n37781 = n37780 ^ n37683;
  assign n37782 = ~n37684 & ~n37781;
  assign n37783 = n37782 ^ n35039;
  assign n37815 = n37783 ^ n34292;
  assign n37502 = n37501 ^ n37497;
  assign n37652 = n37651 ^ n37497;
  assign n37653 = n37502 & n37652;
  assign n37654 = n37653 ^ n37501;
  assign n37492 = n35806 ^ n34879;
  assign n37493 = n37244 ^ n35806;
  assign n37494 = n37492 & ~n37493;
  assign n37495 = n37494 ^ n34879;
  assign n37679 = n37654 ^ n37495;
  assign n37491 = n37198 ^ n37134;
  assign n37680 = n37679 ^ n37491;
  assign n37816 = n37815 ^ n37680;
  assign n37817 = n37777 ^ n34997;
  assign n37818 = n37817 ^ n37686;
  assign n37819 = n37774 ^ n34955;
  assign n37820 = n37819 ^ n37688;
  assign n37821 = n37765 ^ n37696;
  assign n37822 = n37759 ^ n37700;
  assign n37823 = n37756 ^ n37702;
  assign n37824 = n37753 ^ n37704;
  assign n37828 = ~n37826 & n37827;
  assign n37829 = n37730 ^ n33848;
  assign n37830 = n37829 ^ n37719;
  assign n37831 = ~n37828 & ~n37830;
  assign n37832 = n37733 ^ n33841;
  assign n37833 = n37832 ^ n37716;
  assign n37834 = n37831 & n37833;
  assign n37835 = n37736 ^ n34388;
  assign n37836 = n37835 ^ n37713;
  assign n37837 = ~n37834 & ~n37836;
  assign n37838 = n37739 ^ n37711;
  assign n37839 = n37837 & n37838;
  assign n37840 = n37742 ^ n37709;
  assign n37841 = n37839 & ~n37840;
  assign n37842 = n37745 ^ n37706;
  assign n37843 = n37841 & n37842;
  assign n37844 = n37750 ^ n33797;
  assign n37845 = ~n37843 & n37844;
  assign n37846 = n37824 & ~n37845;
  assign n37847 = n37823 & n37846;
  assign n37848 = ~n37822 & n37847;
  assign n37849 = n37762 ^ n37698;
  assign n37850 = ~n37848 & ~n37849;
  assign n37851 = n37821 & ~n37850;
  assign n37852 = n37768 ^ n37694;
  assign n37853 = n37851 & n37852;
  assign n37854 = n37771 ^ n37692;
  assign n37855 = ~n37853 & n37854;
  assign n37856 = ~n37820 & n37855;
  assign n37857 = ~n37818 & n37856;
  assign n37858 = n37780 ^ n37684;
  assign n37859 = ~n37857 & ~n37858;
  assign n37860 = n37816 & n37859;
  assign n37681 = n37680 ^ n34292;
  assign n37784 = n37783 ^ n37680;
  assign n37785 = ~n37681 & ~n37784;
  assign n37786 = n37785 ^ n34292;
  assign n37813 = n37786 ^ n34290;
  assign n37496 = n37495 ^ n37491;
  assign n37655 = n37654 ^ n37491;
  assign n37656 = n37496 & n37655;
  assign n37657 = n37656 ^ n37495;
  assign n37485 = n35803 ^ n34915;
  assign n37486 = n37307 ^ n35803;
  assign n37487 = n37485 & ~n37486;
  assign n37488 = n37487 ^ n34915;
  assign n37676 = n37657 ^ n37488;
  assign n37489 = n37201 ^ n37129;
  assign n37677 = n37676 ^ n37489;
  assign n37814 = n37813 ^ n37677;
  assign n37883 = n37860 ^ n37814;
  assign n1365 = n1274 ^ n1197;
  assign n1375 = n1374 ^ n1365;
  assign n1382 = n1381 ^ n1375;
  assign n37884 = n37883 ^ n1382;
  assign n38023 = n37859 ^ n37816;
  assign n37885 = n37858 ^ n37857;
  assign n37889 = n37888 ^ n37885;
  assign n37893 = n37856 ^ n37818;
  assign n37894 = n37893 ^ n37892;
  assign n37896 = n35619 ^ n27068;
  assign n37897 = n37896 ^ n31617;
  assign n37898 = n37897 ^ n828;
  assign n37895 = n37855 ^ n37820;
  assign n37899 = n37898 ^ n37895;
  assign n37900 = n37854 ^ n37853;
  assign n726 = n725 ^ n707;
  assign n739 = n738 ^ n726;
  assign n752 = n751 ^ n739;
  assign n37901 = n37900 ^ n752;
  assign n37903 = n35625 ^ n27055;
  assign n37904 = n37903 ^ n31624;
  assign n37905 = n37904 ^ n749;
  assign n37902 = n37852 ^ n37851;
  assign n37906 = n37905 ^ n37902;
  assign n37908 = n35631 ^ n675;
  assign n37909 = n37908 ^ n31629;
  assign n37910 = n37909 ^ n25632;
  assign n37907 = n37850 ^ n37821;
  assign n37911 = n37910 ^ n37907;
  assign n37912 = n37849 ^ n37848;
  assign n37916 = n37915 ^ n37912;
  assign n37917 = n37847 ^ n37822;
  assign n37921 = n37920 ^ n37917;
  assign n37922 = n37846 ^ n37823;
  assign n37926 = n37925 ^ n37922;
  assign n37930 = n37845 ^ n37824;
  assign n37927 = n35650 ^ n26935;
  assign n37928 = n37927 ^ n31202;
  assign n37929 = n37928 ^ n25719;
  assign n37931 = n37930 ^ n37929;
  assign n37985 = n37844 ^ n37843;
  assign n37932 = n37842 ^ n37841;
  assign n37936 = n37935 ^ n37932;
  assign n37974 = n37840 ^ n37839;
  assign n37937 = n37838 ^ n37837;
  assign n37941 = n37940 ^ n37937;
  assign n37966 = n37836 ^ n37834;
  assign n37945 = n37833 ^ n37831;
  assign n37946 = n37945 ^ n37944;
  assign n37958 = n37830 ^ n37828;
  assign n37955 = n37954 ^ n37950;
  assign n37956 = n37951 & ~n37955;
  assign n37957 = n37956 ^ n37949;
  assign n37959 = n37958 ^ n37957;
  assign n1777 = n1770 ^ n1737;
  assign n1796 = n1795 ^ n1777;
  assign n1803 = n1802 ^ n1796;
  assign n37960 = n37958 ^ n1803;
  assign n37961 = ~n37959 & n37960;
  assign n37962 = n37961 ^ n1803;
  assign n37963 = n37962 ^ n37945;
  assign n37964 = n37946 & ~n37963;
  assign n37965 = n37964 ^ n37944;
  assign n37967 = n37966 ^ n37965;
  assign n1911 = n1910 ^ n1847;
  assign n1924 = n1923 ^ n1911;
  assign n1931 = n1930 ^ n1924;
  assign n37968 = n37966 ^ n1931;
  assign n37969 = n37967 & ~n37968;
  assign n37970 = n37969 ^ n1931;
  assign n37971 = n37970 ^ n37937;
  assign n37972 = ~n37941 & n37971;
  assign n37973 = n37972 ^ n37940;
  assign n37975 = n37974 ^ n37973;
  assign n37976 = n35666 ^ n26950;
  assign n37977 = n37976 ^ n2087;
  assign n37978 = n37977 ^ n25695;
  assign n37979 = n37978 ^ n37974;
  assign n37980 = ~n37975 & n37979;
  assign n37981 = n37980 ^ n37978;
  assign n37982 = n37981 ^ n37932;
  assign n37983 = ~n37936 & n37982;
  assign n37984 = n37983 ^ n37935;
  assign n37986 = n37985 ^ n37984;
  assign n37990 = n37989 ^ n37985;
  assign n37991 = n37986 & ~n37990;
  assign n37992 = n37991 ^ n37989;
  assign n37993 = n37992 ^ n37930;
  assign n37994 = n37931 & ~n37993;
  assign n37995 = n37994 ^ n37929;
  assign n37996 = n37995 ^ n37922;
  assign n37997 = ~n37926 & n37996;
  assign n37998 = n37997 ^ n37925;
  assign n37999 = n37998 ^ n37917;
  assign n38000 = n37921 & ~n37999;
  assign n38001 = n38000 ^ n37920;
  assign n38002 = n38001 ^ n37912;
  assign n38003 = n37916 & ~n38002;
  assign n38004 = n38003 ^ n37915;
  assign n38005 = n38004 ^ n37907;
  assign n38006 = n37911 & ~n38005;
  assign n38007 = n38006 ^ n37910;
  assign n38008 = n38007 ^ n37902;
  assign n38009 = ~n37906 & n38008;
  assign n38010 = n38009 ^ n37905;
  assign n38011 = n38010 ^ n37900;
  assign n38012 = ~n37901 & n38011;
  assign n38013 = n38012 ^ n752;
  assign n38014 = n38013 ^ n37895;
  assign n38015 = ~n37899 & n38014;
  assign n38016 = n38015 ^ n37898;
  assign n38017 = n38016 ^ n37893;
  assign n38018 = ~n37894 & n38017;
  assign n38019 = n38018 ^ n37892;
  assign n38020 = n38019 ^ n37885;
  assign n38021 = ~n37889 & n38020;
  assign n38022 = n38021 ^ n37888;
  assign n38024 = n38023 ^ n38022;
  assign n38028 = n38027 ^ n38023;
  assign n38029 = n38024 & ~n38028;
  assign n38030 = n38029 ^ n38027;
  assign n38031 = n38030 ^ n37883;
  assign n38032 = ~n37884 & n38031;
  assign n38033 = n38032 ^ n1382;
  assign n37678 = n37677 ^ n34290;
  assign n37787 = n37786 ^ n37677;
  assign n37788 = n37678 & n37787;
  assign n37789 = n37788 ^ n34290;
  assign n37862 = n37789 ^ n34284;
  assign n37490 = n37489 ^ n37488;
  assign n37658 = n37657 ^ n37489;
  assign n37659 = ~n37490 & ~n37658;
  assign n37660 = n37659 ^ n37488;
  assign n37480 = n35797 ^ n34960;
  assign n37481 = n36576 ^ n35797;
  assign n37482 = n37480 & n37481;
  assign n37483 = n37482 ^ n34960;
  assign n37673 = n37660 ^ n37483;
  assign n37479 = n37204 ^ n37124;
  assign n37674 = n37673 ^ n37479;
  assign n37863 = n37862 ^ n37674;
  assign n37861 = n37814 & n37860;
  assign n37881 = n37863 ^ n37861;
  assign n1392 = n1352 ^ n1289;
  assign n1393 = n1392 ^ n1389;
  assign n1397 = n1396 ^ n1393;
  assign n37882 = n37881 ^ n1397;
  assign n38086 = n38033 ^ n37882;
  assign n38159 = n38090 ^ n38086;
  assign n38160 = ~n35281 & ~n38159;
  assign n38161 = n38160 ^ n35279;
  assign n38034 = n38033 ^ n37881;
  assign n38035 = n37882 & ~n38034;
  assign n38036 = n38035 ^ n1397;
  assign n37864 = n37861 & ~n37863;
  assign n37675 = n37674 ^ n34284;
  assign n37790 = n37789 ^ n37674;
  assign n37791 = n37675 & n37790;
  assign n37792 = n37791 ^ n34284;
  assign n37811 = n37792 ^ n34278;
  assign n37484 = n37483 ^ n37479;
  assign n37661 = n37660 ^ n37479;
  assign n37662 = ~n37484 & ~n37661;
  assign n37663 = n37662 ^ n37483;
  assign n37474 = n35790 ^ n35006;
  assign n37475 = n36573 ^ n35790;
  assign n37476 = ~n37474 & n37475;
  assign n37477 = n37476 ^ n35006;
  assign n37670 = n37663 ^ n37477;
  assign n37473 = n37207 ^ n37119;
  assign n37671 = n37670 ^ n37473;
  assign n37812 = n37811 ^ n37671;
  assign n37879 = n37864 ^ n37812;
  assign n37876 = n35595 ^ n2332;
  assign n37877 = n37876 ^ n25775;
  assign n37878 = n37877 ^ n1407;
  assign n37880 = n37879 ^ n37878;
  assign n38093 = n38036 ^ n37880;
  assign n38091 = n38086 & ~n38090;
  assign n38082 = n36086 ^ n35132;
  assign n38083 = n37414 ^ n36086;
  assign n38084 = ~n38082 & n38083;
  assign n38085 = n38084 ^ n35132;
  assign n38092 = n38091 ^ n38085;
  assign n38162 = n38093 ^ n38092;
  assign n38163 = n38162 ^ n38160;
  assign n38164 = n38161 & ~n38163;
  assign n38165 = n38164 ^ n35279;
  assign n38094 = n38093 ^ n38085;
  assign n38095 = n38092 & ~n38094;
  assign n38096 = n38095 ^ n38091;
  assign n38076 = n36079 ^ n35119;
  assign n38077 = n37586 ^ n36079;
  assign n38078 = ~n38076 & ~n38077;
  assign n38079 = n38078 ^ n35119;
  assign n38156 = n38096 ^ n38079;
  assign n38037 = n38036 ^ n37878;
  assign n38038 = n37880 & ~n38037;
  assign n38039 = n38038 ^ n37879;
  assign n37872 = n35590 ^ n2344;
  assign n37873 = n37872 ^ n31594;
  assign n37874 = n37873 ^ n2457;
  assign n37672 = n37671 ^ n34278;
  assign n37793 = n37792 ^ n37671;
  assign n37794 = n37672 & ~n37793;
  assign n37795 = n37794 ^ n34278;
  assign n37866 = n37795 ^ n34265;
  assign n37478 = n37477 ^ n37473;
  assign n37664 = n37663 ^ n37473;
  assign n37665 = n37478 & n37664;
  assign n37666 = n37665 ^ n37477;
  assign n37472 = n37210 ^ n37114;
  assign n37667 = n37666 ^ n37472;
  assign n37468 = n35784 ^ n35049;
  assign n37469 = n36567 ^ n35784;
  assign n37470 = ~n37468 & ~n37469;
  assign n37471 = n37470 ^ n35049;
  assign n37668 = n37667 ^ n37471;
  assign n37867 = n37866 ^ n37668;
  assign n37865 = ~n37812 & ~n37864;
  assign n37871 = n37867 ^ n37865;
  assign n37875 = n37874 ^ n37871;
  assign n38080 = n38039 ^ n37875;
  assign n38157 = n38156 ^ n38080;
  assign n38158 = n38157 ^ n35152;
  assign n38216 = n38165 ^ n38158;
  assign n38166 = n38165 ^ n38157;
  assign n38167 = ~n38158 & ~n38166;
  assign n38168 = n38167 ^ n35152;
  assign n38081 = n38080 ^ n38079;
  assign n38097 = n38096 ^ n38080;
  assign n38098 = n38081 & n38097;
  assign n38099 = n38098 ^ n38079;
  assign n38071 = n36070 ^ n35111;
  assign n38072 = n37580 ^ n36070;
  assign n38073 = ~n38071 & n38072;
  assign n38074 = n38073 ^ n35111;
  assign n38153 = n38099 ^ n38074;
  assign n38040 = n38039 ^ n37871;
  assign n38041 = ~n37875 & n38040;
  assign n38042 = n38041 ^ n37874;
  assign n37868 = n37865 & ~n37867;
  assign n37805 = n37472 ^ n37471;
  assign n37806 = ~n37667 & n37805;
  assign n37807 = n37806 ^ n37471;
  assign n37804 = n37213 ^ n37112;
  assign n37808 = n37807 ^ n37804;
  assign n37800 = n35142 ^ n35104;
  assign n37801 = n36560 ^ n35142;
  assign n37802 = n37800 & n37801;
  assign n37803 = n37802 ^ n35104;
  assign n37809 = n37808 ^ n37803;
  assign n37669 = n37668 ^ n34265;
  assign n37796 = n37795 ^ n37668;
  assign n37797 = n37669 & n37796;
  assign n37798 = n37797 ^ n34265;
  assign n37799 = n37798 ^ n33873;
  assign n37810 = n37809 ^ n37799;
  assign n37869 = n37868 ^ n37810;
  assign n2434 = n2423 ^ n2397;
  assign n2447 = n2446 ^ n2434;
  assign n2460 = n2459 ^ n2447;
  assign n37870 = n37869 ^ n2460;
  assign n38070 = n38042 ^ n37870;
  assign n38154 = n38153 ^ n38070;
  assign n38155 = n38154 ^ n35145;
  assign n38217 = n38168 ^ n38155;
  assign n38218 = n38216 & ~n38217;
  assign n38169 = n38168 ^ n38154;
  assign n38170 = ~n38155 & n38169;
  assign n38171 = n38170 ^ n35145;
  assign n38075 = n38074 ^ n38070;
  assign n38100 = n38099 ^ n38070;
  assign n38101 = ~n38075 & n38100;
  assign n38102 = n38101 ^ n38074;
  assign n38066 = n37810 & n37868;
  assign n38062 = n37216 ^ n37110;
  assign n38059 = n37804 ^ n37803;
  assign n38060 = ~n37808 & ~n38059;
  assign n38061 = n38060 ^ n37803;
  assign n38063 = n38062 ^ n38061;
  assign n38055 = n35827 ^ n35287;
  assign n38056 = n36554 ^ n35827;
  assign n38057 = ~n38055 & ~n38056;
  assign n38058 = n38057 ^ n35287;
  assign n38064 = n38063 ^ n38058;
  assign n38050 = n37809 ^ n33873;
  assign n38051 = n37809 ^ n37798;
  assign n38052 = n38050 & n38051;
  assign n38053 = n38052 ^ n33873;
  assign n38054 = n38053 ^ n33867;
  assign n38065 = n38064 ^ n38054;
  assign n38067 = n38066 ^ n38065;
  assign n38046 = n35583 ^ n27232;
  assign n38047 = n38046 ^ n2576;
  assign n38048 = n38047 ^ n2467;
  assign n38043 = n38042 ^ n37869;
  assign n38044 = n37870 & ~n38043;
  assign n38045 = n38044 ^ n2460;
  assign n38049 = n38048 ^ n38045;
  assign n38068 = n38067 ^ n38049;
  assign n37463 = n36775 ^ n35852;
  assign n37465 = n37464 ^ n36775;
  assign n37466 = n37463 & n37465;
  assign n37467 = n37466 ^ n35852;
  assign n38069 = n38068 ^ n37467;
  assign n38151 = n38102 ^ n38069;
  assign n38152 = n38151 ^ n35267;
  assign n38215 = n38171 ^ n38152;
  assign n38264 = n38218 ^ n38215;
  assign n38261 = n35988 ^ n27197;
  assign n38262 = n38261 ^ n31905;
  assign n38263 = n38262 ^ n1532;
  assign n38265 = n38264 ^ n38263;
  assign n38286 = n38217 ^ n38216;
  assign n38266 = n35999 ^ n26154;
  assign n38267 = n38266 ^ n27119;
  assign n38268 = n38267 ^ n31919;
  assign n38269 = n38268 ^ n38216;
  assign n38270 = n28042 ^ n2602;
  assign n38271 = n38270 ^ n26590;
  assign n38272 = n38271 ^ n32538;
  assign n38273 = n38159 ^ n35281;
  assign n38274 = n38272 & n38273;
  assign n38278 = n38277 ^ n38274;
  assign n38279 = n38162 ^ n38161;
  assign n38280 = n38279 ^ n38277;
  assign n38281 = n38278 & ~n38280;
  assign n38282 = n38281 ^ n38274;
  assign n38283 = n38282 ^ n38216;
  assign n38284 = n38269 & ~n38283;
  assign n38285 = n38284 ^ n38268;
  assign n38287 = n38286 ^ n38285;
  assign n38288 = n35993 ^ n1559;
  assign n38289 = n38288 ^ n26164;
  assign n38290 = n38289 ^ n31910;
  assign n38291 = n38290 ^ n38286;
  assign n38292 = ~n38287 & n38291;
  assign n38293 = n38292 ^ n38290;
  assign n38294 = n38293 ^ n38264;
  assign n38295 = ~n38265 & n38294;
  assign n38296 = n38295 ^ n38263;
  assign n38257 = n35984 ^ n27284;
  assign n38258 = n38257 ^ n1565;
  assign n38259 = n38258 ^ n26149;
  assign n38172 = n38171 ^ n38151;
  assign n38173 = n38152 & ~n38172;
  assign n38174 = n38173 ^ n35267;
  assign n38103 = n38102 ^ n38068;
  assign n38104 = n38069 & n38103;
  assign n38105 = n38104 ^ n37467;
  assign n37457 = n36877 ^ n35922;
  assign n37459 = n37458 ^ n36877;
  assign n37460 = ~n37457 & n37459;
  assign n37461 = n37460 ^ n35922;
  assign n37456 = n37375 ^ n2579;
  assign n37462 = n37461 ^ n37456;
  assign n38149 = n38105 ^ n37462;
  assign n38150 = n38149 ^ n35137;
  assign n38220 = n38174 ^ n38150;
  assign n38219 = n38215 & n38218;
  assign n38256 = n38220 ^ n38219;
  assign n38260 = n38259 ^ n38256;
  assign n38904 = n38296 ^ n38260;
  assign n39430 = n38904 ^ n38131;
  assign n39431 = n39429 & n39430;
  assign n39432 = n39431 ^ n37444;
  assign n38510 = n37244 ^ n36355;
  assign n38511 = n37473 ^ n37244;
  assign n38512 = ~n38510 & n38511;
  assign n38513 = n38512 ^ n36355;
  assign n38392 = n38001 ^ n37916;
  assign n38514 = n38513 ^ n38392;
  assign n38515 = n37096 ^ n36256;
  assign n38516 = n37479 ^ n37096;
  assign n38517 = n38515 & ~n38516;
  assign n38518 = n38517 ^ n36256;
  assign n38399 = n37998 ^ n37921;
  assign n38519 = n38518 ^ n38399;
  assign n38520 = n37077 ^ n36110;
  assign n38521 = n37489 ^ n37077;
  assign n38522 = ~n38520 & ~n38521;
  assign n38523 = n38522 ^ n36110;
  assign n38406 = n37995 ^ n37926;
  assign n38524 = n38523 ^ n38406;
  assign n38525 = n37021 ^ n36116;
  assign n38526 = n37491 ^ n37021;
  assign n38527 = n38525 & ~n38526;
  assign n38528 = n38527 ^ n36116;
  assign n38413 = n37992 ^ n37931;
  assign n38529 = n38528 ^ n38413;
  assign n38530 = n36929 ^ n36126;
  assign n38531 = n37497 ^ n36929;
  assign n38532 = ~n38530 & n38531;
  assign n38533 = n38532 ^ n36126;
  assign n38420 = n37989 ^ n37986;
  assign n38534 = n38533 ^ n38420;
  assign n38535 = n36795 ^ n36133;
  assign n38536 = n37503 ^ n36795;
  assign n38537 = ~n38535 & ~n38536;
  assign n38538 = n38537 ^ n36133;
  assign n38427 = n37981 ^ n37936;
  assign n38539 = n38538 ^ n38427;
  assign n38540 = n36802 ^ n36140;
  assign n38541 = n37509 ^ n36802;
  assign n38542 = n38540 & ~n38541;
  assign n38543 = n38542 ^ n36140;
  assign n38434 = n37978 ^ n37975;
  assign n38544 = n38543 ^ n38434;
  assign n38545 = n36808 ^ n36146;
  assign n38546 = n37510 ^ n36808;
  assign n38547 = ~n38545 & ~n38546;
  assign n38548 = n38547 ^ n36146;
  assign n38440 = n37970 ^ n37941;
  assign n38549 = n38548 ^ n38440;
  assign n38362 = n36810 ^ n36152;
  assign n38363 = n37516 ^ n36810;
  assign n38364 = n38362 & ~n38363;
  assign n38365 = n38364 ^ n36152;
  assign n38361 = n37967 ^ n1931;
  assign n38366 = n38365 ^ n38361;
  assign n38341 = n37962 ^ n37946;
  assign n38337 = n36816 ^ n36220;
  assign n38338 = n37526 ^ n36816;
  assign n38339 = n38337 & ~n38338;
  assign n38340 = n38339 ^ n36220;
  assign n38342 = n38341 ^ n38340;
  assign n38206 = n37959 ^ n1803;
  assign n38202 = n36823 ^ n36159;
  assign n38203 = n37532 ^ n36823;
  assign n38204 = ~n38202 & ~n38203;
  assign n38205 = n38204 ^ n36159;
  assign n38207 = n38206 ^ n38205;
  assign n38127 = n36833 ^ n36165;
  assign n38128 = n37538 ^ n36833;
  assign n38129 = n38127 & ~n38128;
  assign n38130 = n38129 ^ n36165;
  assign n38132 = n38131 ^ n38130;
  assign n37419 = n37418 ^ n37396;
  assign n36063 = n36062 ^ n36060;
  assign n36783 = n36782 ^ n36060;
  assign n36784 = ~n36063 & n36783;
  assign n36785 = n36784 ^ n36062;
  assign n37420 = n37419 ^ n36785;
  assign n37426 = n37393 ^ n37360;
  assign n37421 = n36840 ^ n36176;
  assign n37423 = n37422 ^ n36840;
  assign n37424 = n37421 & ~n37423;
  assign n37425 = n37424 ^ n36176;
  assign n37427 = n37426 ^ n37425;
  assign n37429 = n36847 ^ n36183;
  assign n37431 = n37430 ^ n36847;
  assign n37432 = ~n37429 & n37431;
  assign n37433 = n37432 ^ n36183;
  assign n37428 = n37390 ^ n37365;
  assign n37434 = n37433 ^ n37428;
  assign n37436 = n36853 ^ n36065;
  assign n37438 = n37437 ^ n36853;
  assign n37439 = ~n37436 & n37438;
  assign n37440 = n37439 ^ n36065;
  assign n37435 = n37387 ^ n37370;
  assign n37441 = n37440 ^ n37435;
  assign n37443 = n36860 ^ n36074;
  assign n37445 = n37444 ^ n36860;
  assign n37446 = ~n37443 & n37445;
  assign n37447 = n37446 ^ n36074;
  assign n37442 = n37384 ^ n37374;
  assign n37448 = n37447 ^ n37442;
  assign n37450 = n36866 ^ n36054;
  assign n37452 = n37451 ^ n36866;
  assign n37453 = ~n37450 & ~n37452;
  assign n37454 = n37453 ^ n36054;
  assign n37449 = n37381 ^ n37380;
  assign n37455 = n37454 ^ n37449;
  assign n38106 = n38105 ^ n37456;
  assign n38107 = n37462 & n38106;
  assign n38108 = n38107 ^ n37461;
  assign n38109 = n38108 ^ n37449;
  assign n38110 = n37455 & n38109;
  assign n38111 = n38110 ^ n37454;
  assign n38112 = n38111 ^ n37442;
  assign n38113 = ~n37448 & n38112;
  assign n38114 = n38113 ^ n37447;
  assign n38115 = n38114 ^ n37435;
  assign n38116 = n37441 & n38115;
  assign n38117 = n38116 ^ n37440;
  assign n38118 = n38117 ^ n37428;
  assign n38119 = ~n37434 & n38118;
  assign n38120 = n38119 ^ n37433;
  assign n38121 = n38120 ^ n37426;
  assign n38122 = n37427 & ~n38121;
  assign n38123 = n38122 ^ n37425;
  assign n38124 = n38123 ^ n37419;
  assign n38125 = n37420 & ~n38124;
  assign n38126 = n38125 ^ n36785;
  assign n38199 = n38131 ^ n38126;
  assign n38200 = n38132 & n38199;
  assign n38201 = n38200 ^ n38130;
  assign n38334 = n38206 ^ n38201;
  assign n38335 = ~n38207 & ~n38334;
  assign n38336 = n38335 ^ n38205;
  assign n38358 = n38341 ^ n38336;
  assign n38359 = n38342 & n38358;
  assign n38360 = n38359 ^ n38340;
  assign n38550 = n38361 ^ n38360;
  assign n38551 = ~n38366 & n38550;
  assign n38552 = n38551 ^ n38365;
  assign n38553 = n38552 ^ n38440;
  assign n38554 = ~n38549 & n38553;
  assign n38555 = n38554 ^ n38548;
  assign n38556 = n38555 ^ n38434;
  assign n38557 = n38544 & ~n38556;
  assign n38558 = n38557 ^ n38543;
  assign n38559 = n38558 ^ n38427;
  assign n38560 = n38539 & n38559;
  assign n38561 = n38560 ^ n38538;
  assign n38562 = n38561 ^ n38420;
  assign n38563 = ~n38534 & ~n38562;
  assign n38564 = n38563 ^ n38533;
  assign n38565 = n38564 ^ n38413;
  assign n38566 = ~n38529 & ~n38565;
  assign n38567 = n38566 ^ n38528;
  assign n38568 = n38567 ^ n38406;
  assign n38569 = ~n38524 & ~n38568;
  assign n38570 = n38569 ^ n38523;
  assign n38571 = n38570 ^ n38399;
  assign n38572 = n38519 & ~n38571;
  assign n38573 = n38572 ^ n38518;
  assign n38574 = n38573 ^ n38392;
  assign n38575 = n38514 & ~n38574;
  assign n38576 = n38575 ^ n38513;
  assign n38505 = n37307 ^ n36544;
  assign n38506 = n37472 ^ n37307;
  assign n38507 = n38505 & ~n38506;
  assign n38508 = n38507 ^ n36544;
  assign n38604 = n38576 ^ n38508;
  assign n38385 = n38004 ^ n37911;
  assign n38605 = n38604 ^ n38385;
  assign n38606 = n38605 ^ n35779;
  assign n38607 = n38573 ^ n38514;
  assign n38608 = n38607 ^ n35514;
  assign n38609 = n38570 ^ n38519;
  assign n38610 = n38609 ^ n35157;
  assign n38611 = n38567 ^ n38524;
  assign n38612 = n38611 ^ n35158;
  assign n38613 = n38564 ^ n38529;
  assign n38614 = n38613 ^ n35165;
  assign n38615 = n38561 ^ n38534;
  assign n38616 = n38615 ^ n35175;
  assign n38617 = n38558 ^ n38539;
  assign n38618 = n38617 ^ n35178;
  assign n38619 = n38555 ^ n38544;
  assign n38620 = n38619 ^ n35185;
  assign n38621 = n38552 ^ n38548;
  assign n38622 = n38621 ^ n38440;
  assign n38623 = n38622 ^ n35191;
  assign n38367 = n38366 ^ n38360;
  assign n38368 = n38367 ^ n35197;
  assign n38343 = n38342 ^ n38336;
  assign n38344 = n38343 ^ n35203;
  assign n38208 = n38207 ^ n38201;
  assign n38209 = n38208 ^ n35210;
  assign n38133 = n38132 ^ n38126;
  assign n38134 = n38133 ^ n35220;
  assign n38135 = n38123 ^ n37420;
  assign n38136 = n38135 ^ n35227;
  assign n38137 = n38120 ^ n37427;
  assign n38138 = n38137 ^ n35234;
  assign n38139 = n38117 ^ n37434;
  assign n38140 = n38139 ^ n35241;
  assign n38141 = n38114 ^ n37440;
  assign n38142 = n38141 ^ n37435;
  assign n38143 = n38142 ^ n35113;
  assign n38144 = n38111 ^ n37448;
  assign n38145 = n38144 ^ n35122;
  assign n38146 = n38108 ^ n37454;
  assign n38147 = n38146 ^ n37449;
  assign n38148 = n38147 ^ n35128;
  assign n38175 = n38174 ^ n38149;
  assign n38176 = ~n38150 & n38175;
  assign n38177 = n38176 ^ n35137;
  assign n38178 = n38177 ^ n38147;
  assign n38179 = ~n38148 & ~n38178;
  assign n38180 = n38179 ^ n35128;
  assign n38181 = n38180 ^ n38144;
  assign n38182 = n38145 & n38181;
  assign n38183 = n38182 ^ n35122;
  assign n38184 = n38183 ^ n38142;
  assign n38185 = n38143 & n38184;
  assign n38186 = n38185 ^ n35113;
  assign n38187 = n38186 ^ n38139;
  assign n38188 = ~n38140 & ~n38187;
  assign n38189 = n38188 ^ n35241;
  assign n38190 = n38189 ^ n38137;
  assign n38191 = n38138 & ~n38190;
  assign n38192 = n38191 ^ n35234;
  assign n38193 = n38192 ^ n38135;
  assign n38194 = n38136 & ~n38193;
  assign n38195 = n38194 ^ n35227;
  assign n38196 = n38195 ^ n38133;
  assign n38197 = ~n38134 & ~n38196;
  assign n38198 = n38197 ^ n35220;
  assign n38331 = n38208 ^ n38198;
  assign n38332 = ~n38209 & n38331;
  assign n38333 = n38332 ^ n35210;
  assign n38355 = n38343 ^ n38333;
  assign n38356 = ~n38344 & n38355;
  assign n38357 = n38356 ^ n35203;
  assign n38624 = n38367 ^ n38357;
  assign n38625 = n38368 & n38624;
  assign n38626 = n38625 ^ n35197;
  assign n38627 = n38626 ^ n38622;
  assign n38628 = ~n38623 & ~n38627;
  assign n38629 = n38628 ^ n35191;
  assign n38630 = n38629 ^ n38619;
  assign n38631 = ~n38620 & ~n38630;
  assign n38632 = n38631 ^ n35185;
  assign n38633 = n38632 ^ n38617;
  assign n38634 = n38618 & n38633;
  assign n38635 = n38634 ^ n35178;
  assign n38636 = n38635 ^ n38615;
  assign n38637 = n38616 & ~n38636;
  assign n38638 = n38637 ^ n35175;
  assign n38639 = n38638 ^ n38613;
  assign n38640 = ~n38614 & n38639;
  assign n38641 = n38640 ^ n35165;
  assign n38642 = n38641 ^ n38611;
  assign n38643 = ~n38612 & ~n38642;
  assign n38644 = n38643 ^ n35158;
  assign n38645 = n38644 ^ n38609;
  assign n38646 = n38610 & n38645;
  assign n38647 = n38646 ^ n35157;
  assign n38648 = n38647 ^ n38607;
  assign n38649 = ~n38608 & ~n38648;
  assign n38650 = n38649 ^ n35514;
  assign n38651 = n38650 ^ n38605;
  assign n38652 = n38606 & n38651;
  assign n38653 = n38652 ^ n35779;
  assign n38509 = n38508 ^ n38385;
  assign n38577 = n38576 ^ n38385;
  assign n38578 = n38509 & ~n38577;
  assign n38579 = n38578 ^ n38508;
  assign n38500 = n36576 ^ n35806;
  assign n38501 = n37804 ^ n36576;
  assign n38502 = ~n38500 & ~n38501;
  assign n38503 = n38502 ^ n35806;
  assign n38378 = n38007 ^ n37906;
  assign n38504 = n38503 ^ n38378;
  assign n38602 = n38579 ^ n38504;
  assign n38603 = n38602 ^ n34879;
  assign n38683 = n38653 ^ n38603;
  assign n38684 = n38635 ^ n38616;
  assign n38685 = n38629 ^ n38620;
  assign n38369 = n38368 ^ n38357;
  assign n38345 = n38344 ^ n38333;
  assign n38210 = n38209 ^ n38198;
  assign n38211 = n38192 ^ n38136;
  assign n38212 = n38189 ^ n38138;
  assign n38213 = n38186 ^ n38140;
  assign n38214 = n38183 ^ n38143;
  assign n38221 = ~n38219 & n38220;
  assign n38222 = n38177 ^ n38148;
  assign n38223 = ~n38221 & ~n38222;
  assign n38224 = n38180 ^ n38145;
  assign n38225 = n38223 & ~n38224;
  assign n38226 = ~n38214 & ~n38225;
  assign n38227 = ~n38213 & n38226;
  assign n38228 = n38212 & ~n38227;
  assign n38229 = n38211 & n38228;
  assign n38230 = n38195 ^ n38134;
  assign n38231 = n38229 & ~n38230;
  assign n38346 = n38210 & n38231;
  assign n38370 = ~n38345 & ~n38346;
  assign n38686 = ~n38369 & ~n38370;
  assign n38687 = n38626 ^ n38623;
  assign n38688 = n38686 & ~n38687;
  assign n38689 = n38685 & n38688;
  assign n38690 = n38632 ^ n38618;
  assign n38691 = ~n38689 & ~n38690;
  assign n38692 = ~n38684 & ~n38691;
  assign n38693 = n38638 ^ n38614;
  assign n38694 = n38692 & n38693;
  assign n38695 = n38641 ^ n38612;
  assign n38696 = ~n38694 & ~n38695;
  assign n38697 = n38644 ^ n38610;
  assign n38698 = n38696 & ~n38697;
  assign n38699 = n38647 ^ n38608;
  assign n38700 = n38698 & ~n38699;
  assign n38701 = n38650 ^ n38606;
  assign n38702 = ~n38700 & n38701;
  assign n38703 = n38683 & n38702;
  assign n38654 = n38653 ^ n38602;
  assign n38655 = ~n38603 & ~n38654;
  assign n38656 = n38655 ^ n34879;
  assign n38580 = n38579 ^ n38378;
  assign n38581 = n38504 & n38580;
  assign n38582 = n38581 ^ n38503;
  assign n38498 = n38010 ^ n37901;
  assign n38494 = n36573 ^ n35803;
  assign n38495 = n38062 ^ n36573;
  assign n38496 = n38494 & ~n38495;
  assign n38497 = n38496 ^ n35803;
  assign n38499 = n38498 ^ n38497;
  assign n38600 = n38582 ^ n38499;
  assign n38601 = n38600 ^ n34915;
  assign n38682 = n38656 ^ n38601;
  assign n38726 = n38703 ^ n38682;
  assign n38723 = n36429 ^ n27983;
  assign n38724 = n38723 ^ n32466;
  assign n38725 = n38724 ^ n1224;
  assign n38727 = n38726 ^ n38725;
  assign n38800 = n38702 ^ n38683;
  assign n38729 = n36436 ^ n27990;
  assign n38730 = n38729 ^ n940;
  assign n38731 = n38730 ^ n1061;
  assign n38728 = n38701 ^ n38700;
  assign n38732 = n38731 ^ n38728;
  assign n38733 = n38699 ^ n38698;
  assign n907 = n887 ^ n861;
  assign n920 = n919 ^ n907;
  assign n933 = n932 ^ n920;
  assign n38734 = n38733 ^ n933;
  assign n38736 = n36443 ^ n808;
  assign n38737 = n38736 ^ n32415;
  assign n38738 = n38737 ^ n930;
  assign n38735 = n38697 ^ n38696;
  assign n38739 = n38738 ^ n38735;
  assign n38741 = n36448 ^ n793;
  assign n38742 = n38741 ^ n32420;
  assign n38743 = n38742 ^ n26498;
  assign n38740 = n38695 ^ n38694;
  assign n38744 = n38743 ^ n38740;
  assign n38748 = n38693 ^ n38692;
  assign n38749 = n38748 ^ n38747;
  assign n38753 = n38691 ^ n38684;
  assign n38750 = n36458 ^ n27584;
  assign n38751 = n38750 ^ n32387;
  assign n38752 = n38751 ^ n25808;
  assign n38754 = n38753 ^ n38752;
  assign n38774 = n38690 ^ n38689;
  assign n38756 = n36489 ^ n27594;
  assign n38757 = n38756 ^ n32391;
  assign n38758 = n38757 ^ n626;
  assign n38755 = n38688 ^ n38685;
  assign n38759 = n38758 ^ n38755;
  assign n38763 = n38687 ^ n38686;
  assign n38371 = n38370 ^ n38369;
  assign n38375 = n38374 ^ n38371;
  assign n38347 = n38346 ^ n38345;
  assign n38232 = n38231 ^ n38210;
  assign n38236 = n38235 ^ n38232;
  assign n38323 = n38230 ^ n38229;
  assign n38237 = n38228 ^ n38211;
  assign n38238 = n38237 ^ n2065;
  assign n38239 = n38227 ^ n38212;
  assign n2024 = n2005 ^ n1957;
  assign n2040 = n2039 ^ n2024;
  assign n2047 = n2046 ^ n2040;
  assign n38240 = n38239 ^ n2047;
  assign n38242 = n35963 ^ n1880;
  assign n38243 = n38242 ^ n31884;
  assign n38244 = n38243 ^ n2034;
  assign n38241 = n38226 ^ n38213;
  assign n38245 = n38244 ^ n38241;
  assign n38306 = n38225 ^ n38214;
  assign n38246 = n38224 ^ n38223;
  assign n38250 = n38249 ^ n38246;
  assign n38251 = n38222 ^ n38221;
  assign n38255 = n38254 ^ n38251;
  assign n38297 = n38296 ^ n38256;
  assign n38298 = ~n38260 & n38297;
  assign n38299 = n38298 ^ n38259;
  assign n38300 = n38299 ^ n38251;
  assign n38301 = ~n38255 & n38300;
  assign n38302 = n38301 ^ n38254;
  assign n38303 = n38302 ^ n38246;
  assign n38304 = n38250 & ~n38303;
  assign n38305 = n38304 ^ n38249;
  assign n38307 = n38306 ^ n38305;
  assign n38308 = n35969 ^ n1865;
  assign n38309 = n38308 ^ n31889;
  assign n38310 = n38309 ^ n26137;
  assign n38311 = n38310 ^ n38306;
  assign n38312 = ~n38307 & n38311;
  assign n38313 = n38312 ^ n38310;
  assign n38314 = n38313 ^ n38241;
  assign n38315 = ~n38245 & n38314;
  assign n38316 = n38315 ^ n38244;
  assign n38317 = n38316 ^ n38239;
  assign n38318 = n38240 & ~n38317;
  assign n38319 = n38318 ^ n2047;
  assign n38320 = n38319 ^ n38237;
  assign n38321 = ~n38238 & n38320;
  assign n38322 = n38321 ^ n2065;
  assign n38324 = n38323 ^ n38322;
  assign n2194 = n2190 ^ n2103;
  assign n2201 = n2200 ^ n2194;
  assign n2208 = n2207 ^ n2201;
  assign n38325 = n38323 ^ n2208;
  assign n38326 = ~n38324 & n38325;
  assign n38327 = n38326 ^ n2208;
  assign n38328 = n38327 ^ n38232;
  assign n38329 = ~n38236 & n38328;
  assign n38330 = n38329 ^ n38235;
  assign n38348 = n38347 ^ n38330;
  assign n38352 = n38351 ^ n38347;
  assign n38353 = ~n38348 & n38352;
  assign n38354 = n38353 ^ n38351;
  assign n38760 = n38371 ^ n38354;
  assign n38761 = ~n38375 & n38760;
  assign n38762 = n38761 ^ n38374;
  assign n38764 = n38763 ^ n38762;
  assign n38765 = n36468 ^ n27599;
  assign n38766 = n38765 ^ n32374;
  assign n38767 = n38766 ^ n26217;
  assign n38768 = n38767 ^ n38763;
  assign n38769 = ~n38764 & n38768;
  assign n38770 = n38769 ^ n38767;
  assign n38771 = n38770 ^ n38755;
  assign n38772 = ~n38759 & n38771;
  assign n38773 = n38772 ^ n38758;
  assign n38775 = n38774 ^ n38773;
  assign n38776 = n36463 ^ n27589;
  assign n38777 = n38776 ^ n32397;
  assign n38778 = n38777 ^ n26243;
  assign n38779 = n38778 ^ n38774;
  assign n38780 = ~n38775 & n38779;
  assign n38781 = n38780 ^ n38778;
  assign n38782 = n38781 ^ n38753;
  assign n38783 = ~n38754 & n38782;
  assign n38784 = n38783 ^ n38752;
  assign n38785 = n38784 ^ n38748;
  assign n38786 = ~n38749 & n38785;
  assign n38787 = n38786 ^ n38747;
  assign n38788 = n38787 ^ n38740;
  assign n38789 = n38744 & ~n38788;
  assign n38790 = n38789 ^ n38743;
  assign n38791 = n38790 ^ n38735;
  assign n38792 = ~n38739 & n38791;
  assign n38793 = n38792 ^ n38738;
  assign n38794 = n38793 ^ n38733;
  assign n38795 = ~n38734 & n38794;
  assign n38796 = n38795 ^ n933;
  assign n38797 = n38796 ^ n38728;
  assign n38798 = n38732 & ~n38797;
  assign n38799 = n38798 ^ n38731;
  assign n38801 = n38800 ^ n38799;
  assign n1044 = n1043 ^ n977;
  assign n1057 = n1056 ^ n1044;
  assign n1064 = n1063 ^ n1057;
  assign n38802 = n38800 ^ n1064;
  assign n38803 = n38801 & ~n38802;
  assign n38804 = n38803 ^ n1064;
  assign n38805 = n38804 ^ n38726;
  assign n38806 = ~n38727 & n38805;
  assign n38807 = n38806 ^ n38725;
  assign n38719 = n36424 ^ n27978;
  assign n38720 = n38719 ^ n26487;
  assign n38721 = n38720 ^ n1229;
  assign n38704 = n38682 & n38703;
  assign n38657 = n38656 ^ n38600;
  assign n38658 = n38601 & n38657;
  assign n38659 = n38658 ^ n34915;
  assign n38583 = n38582 ^ n38498;
  assign n38584 = ~n38499 & ~n38583;
  assign n38585 = n38584 ^ n38497;
  assign n38492 = n38013 ^ n37899;
  assign n38488 = n36567 ^ n35797;
  assign n38489 = n37266 ^ n36567;
  assign n38490 = n38488 & ~n38489;
  assign n38491 = n38490 ^ n35797;
  assign n38493 = n38492 ^ n38491;
  assign n38598 = n38585 ^ n38493;
  assign n38599 = n38598 ^ n34960;
  assign n38681 = n38659 ^ n38599;
  assign n38718 = n38704 ^ n38681;
  assign n38722 = n38721 ^ n38718;
  assign n38870 = n38807 ^ n38722;
  assign n38866 = n37586 ^ n36088;
  assign n38867 = n37586 ^ n37456;
  assign n38868 = ~n38866 & n38867;
  assign n38869 = n38868 ^ n36088;
  assign n38992 = n38870 ^ n38869;
  assign n39222 = n38992 ^ n35134;
  assign n39219 = n37292 ^ n28640;
  assign n39220 = n39219 ^ n33369;
  assign n39221 = n39220 ^ n2570;
  assign n39428 = n39222 ^ n39221;
  assign n39433 = n39432 ^ n39428;
  assign n39495 = n38793 ^ n38734;
  assign n39490 = n37254 ^ n36560;
  assign n39491 = n38093 ^ n37254;
  assign n39492 = ~n39490 & n39491;
  assign n39493 = n39492 ^ n36560;
  assign n39467 = n38790 ^ n38739;
  assign n39463 = n37260 ^ n36567;
  assign n39464 = n38086 ^ n37260;
  assign n39465 = ~n39463 & ~n39464;
  assign n39466 = n39465 ^ n36567;
  assign n39468 = n39467 ^ n39466;
  assign n39445 = n38787 ^ n38744;
  assign n39441 = n37273 ^ n36573;
  assign n38833 = n38030 ^ n37884;
  assign n39442 = n38833 ^ n37273;
  assign n39443 = n39441 & n39442;
  assign n39444 = n39443 ^ n36573;
  assign n39446 = n39445 ^ n39444;
  assign n39331 = n38781 ^ n38754;
  assign n39326 = n38062 ^ n37307;
  assign n38592 = n38019 ^ n37889;
  assign n39327 = n38592 ^ n38062;
  assign n39328 = n39326 & n39327;
  assign n39329 = n39328 ^ n37307;
  assign n39448 = n39331 ^ n39329;
  assign n39127 = n37804 ^ n37244;
  assign n38486 = n38016 ^ n37894;
  assign n39128 = n38486 ^ n37804;
  assign n39129 = ~n39127 & n39128;
  assign n39130 = n39129 ^ n37244;
  assign n39126 = n38778 ^ n38775;
  assign n39131 = n39130 ^ n39126;
  assign n39069 = n37472 ^ n37096;
  assign n39070 = n38492 ^ n37472;
  assign n39071 = n39069 & n39070;
  assign n39072 = n39071 ^ n37096;
  assign n39068 = n38770 ^ n38759;
  assign n39073 = n39072 ^ n39068;
  assign n38947 = n38767 ^ n38764;
  assign n38943 = n37473 ^ n37077;
  assign n38944 = n38498 ^ n37473;
  assign n38945 = ~n38943 & n38944;
  assign n38946 = n38945 ^ n37077;
  assign n38948 = n38947 ^ n38946;
  assign n38377 = n37479 ^ n37021;
  assign n38379 = n38378 ^ n37479;
  assign n38380 = ~n38377 & n38379;
  assign n38381 = n38380 ^ n37021;
  assign n38376 = n38375 ^ n38354;
  assign n38382 = n38381 ^ n38376;
  assign n38384 = n37489 ^ n36929;
  assign n38386 = n38385 ^ n37489;
  assign n38387 = n38384 & n38386;
  assign n38388 = n38387 ^ n36929;
  assign n38383 = n38351 ^ n38348;
  assign n38389 = n38388 ^ n38383;
  assign n38391 = n37491 ^ n36795;
  assign n38393 = n38392 ^ n37491;
  assign n38394 = ~n38391 & n38393;
  assign n38395 = n38394 ^ n36795;
  assign n38390 = n38327 ^ n38236;
  assign n38396 = n38395 ^ n38390;
  assign n38398 = n37497 ^ n36802;
  assign n38400 = n38399 ^ n37497;
  assign n38401 = n38398 & ~n38400;
  assign n38402 = n38401 ^ n36802;
  assign n38397 = n38324 ^ n2208;
  assign n38403 = n38402 ^ n38397;
  assign n38405 = n37503 ^ n36808;
  assign n38407 = n38406 ^ n37503;
  assign n38408 = ~n38405 & n38407;
  assign n38409 = n38408 ^ n36808;
  assign n38404 = n38319 ^ n38238;
  assign n38410 = n38409 ^ n38404;
  assign n38412 = n37509 ^ n36810;
  assign n38414 = n38413 ^ n37509;
  assign n38415 = n38412 & ~n38414;
  assign n38416 = n38415 ^ n36810;
  assign n38411 = n38316 ^ n38240;
  assign n38417 = n38416 ^ n38411;
  assign n38419 = n37510 ^ n36816;
  assign n38421 = n38420 ^ n37510;
  assign n38422 = ~n38419 & ~n38421;
  assign n38423 = n38422 ^ n36816;
  assign n38418 = n38313 ^ n38245;
  assign n38424 = n38423 ^ n38418;
  assign n38426 = n37516 ^ n36823;
  assign n38428 = n38427 ^ n37516;
  assign n38429 = n38426 & n38428;
  assign n38430 = n38429 ^ n36823;
  assign n38425 = n38310 ^ n38307;
  assign n38431 = n38430 ^ n38425;
  assign n38433 = n37526 ^ n36833;
  assign n38435 = n38434 ^ n37526;
  assign n38436 = n38433 & ~n38435;
  assign n38437 = n38436 ^ n36833;
  assign n38432 = n38302 ^ n38250;
  assign n38438 = n38437 ^ n38432;
  assign n38444 = n38299 ^ n38255;
  assign n38439 = n37532 ^ n36060;
  assign n38441 = n38440 ^ n37532;
  assign n38442 = n38439 & n38441;
  assign n38443 = n38442 ^ n36060;
  assign n38445 = n38444 ^ n38443;
  assign n38450 = n38293 ^ n38265;
  assign n38446 = n36847 ^ n36782;
  assign n38447 = n38341 ^ n36782;
  assign n38448 = ~n38446 & n38447;
  assign n38449 = n38448 ^ n36847;
  assign n38451 = n38450 ^ n38449;
  assign n38456 = n38290 ^ n38287;
  assign n38452 = n37422 ^ n36853;
  assign n38453 = n38206 ^ n37422;
  assign n38454 = ~n38452 & n38453;
  assign n38455 = n38454 ^ n36853;
  assign n38457 = n38456 ^ n38455;
  assign n38463 = n38279 ^ n38278;
  assign n38459 = n37437 ^ n36866;
  assign n38460 = n37437 ^ n37419;
  assign n38461 = n38459 & ~n38460;
  assign n38462 = n38461 ^ n36866;
  assign n38464 = n38463 ^ n38462;
  assign n38469 = n38273 ^ n38272;
  assign n38465 = n37444 ^ n36877;
  assign n38466 = n37444 ^ n37426;
  assign n38467 = n38465 & n38466;
  assign n38468 = n38467 ^ n36877;
  assign n38470 = n38469 ^ n38468;
  assign n38676 = n38027 ^ n38024;
  assign n38482 = n36560 ^ n35790;
  assign n38483 = n37273 ^ n36560;
  assign n38484 = ~n38482 & ~n38483;
  assign n38485 = n38484 ^ n35790;
  assign n38487 = n38486 ^ n38485;
  assign n38586 = n38585 ^ n38492;
  assign n38587 = n38493 & n38586;
  assign n38588 = n38587 ^ n38491;
  assign n38589 = n38588 ^ n38486;
  assign n38590 = n38487 & ~n38589;
  assign n38591 = n38590 ^ n38485;
  assign n38593 = n38592 ^ n38591;
  assign n38478 = n36554 ^ n35784;
  assign n38479 = n37260 ^ n36554;
  assign n38480 = n38478 & n38479;
  assign n38481 = n38480 ^ n35784;
  assign n38673 = n38592 ^ n38481;
  assign n38674 = ~n38593 & n38673;
  assign n38675 = n38674 ^ n38481;
  assign n38677 = n38676 ^ n38675;
  assign n38669 = n36104 ^ n35142;
  assign n38670 = n37254 ^ n36104;
  assign n38671 = n38669 & ~n38670;
  assign n38672 = n38671 ^ n35142;
  assign n38678 = n38677 ^ n38672;
  assign n38679 = n38678 ^ n35104;
  assign n38594 = n38593 ^ n38481;
  assign n38595 = n38594 ^ n35049;
  assign n38596 = n38588 ^ n38487;
  assign n38597 = n38596 ^ n35006;
  assign n38660 = n38659 ^ n38598;
  assign n38661 = ~n38599 & ~n38660;
  assign n38662 = n38661 ^ n34960;
  assign n38663 = n38662 ^ n38596;
  assign n38664 = ~n38597 & ~n38663;
  assign n38665 = n38664 ^ n35006;
  assign n38666 = n38665 ^ n38594;
  assign n38667 = ~n38595 & n38666;
  assign n38668 = n38667 ^ n35049;
  assign n38680 = n38679 ^ n38668;
  assign n38705 = n38681 & n38704;
  assign n38706 = n38662 ^ n38597;
  assign n38707 = ~n38705 & n38706;
  assign n38708 = n38665 ^ n35049;
  assign n38709 = n38708 ^ n38594;
  assign n38710 = n38707 & ~n38709;
  assign n38844 = n38680 & n38710;
  assign n38837 = n36098 ^ n35827;
  assign n38838 = n37312 ^ n36098;
  assign n38839 = ~n38837 & n38838;
  assign n38840 = n38839 ^ n35827;
  assign n38834 = n38676 ^ n38672;
  assign n38835 = ~n38677 & n38834;
  assign n38836 = n38835 ^ n38672;
  assign n38841 = n38840 ^ n38836;
  assign n38842 = n38841 ^ n38833;
  assign n38829 = n38678 ^ n38668;
  assign n38830 = n38679 & n38829;
  assign n38831 = n38830 ^ n35104;
  assign n38832 = n38831 ^ n35287;
  assign n38843 = n38842 ^ n38832;
  assign n38845 = n38844 ^ n38843;
  assign n38825 = n36404 ^ n2531;
  assign n38826 = n38825 ^ n32369;
  assign n38827 = n38826 ^ n26569;
  assign n38711 = n38710 ^ n38680;
  assign n38475 = n36408 ^ n2516;
  assign n38476 = n38475 ^ n26480;
  assign n38477 = n38476 ^ n32499;
  assign n38712 = n38711 ^ n38477;
  assign n38714 = n36414 ^ n27973;
  assign n38715 = n38714 ^ n32494;
  assign n38716 = n38715 ^ n26543;
  assign n38713 = n38709 ^ n38707;
  assign n38717 = n38716 ^ n38713;
  assign n38811 = n38706 ^ n38705;
  assign n38808 = n38807 ^ n38718;
  assign n38809 = ~n38722 & n38808;
  assign n38810 = n38809 ^ n38721;
  assign n38812 = n38811 ^ n38810;
  assign n38813 = n36419 ^ n2282;
  assign n38814 = n38813 ^ n28011;
  assign n38815 = n38814 ^ n32472;
  assign n38816 = n38815 ^ n38811;
  assign n38817 = n38812 & ~n38816;
  assign n38818 = n38817 ^ n38815;
  assign n38819 = n38818 ^ n38713;
  assign n38820 = ~n38717 & n38819;
  assign n38821 = n38820 ^ n38716;
  assign n38822 = n38821 ^ n38711;
  assign n38823 = n38712 & ~n38822;
  assign n38824 = n38823 ^ n38477;
  assign n38828 = n38827 ^ n38824;
  assign n38846 = n38845 ^ n38828;
  assign n38471 = n37451 ^ n36775;
  assign n38472 = n37451 ^ n37428;
  assign n38473 = ~n38471 & n38472;
  assign n38474 = n38473 ^ n36775;
  assign n38847 = n38846 ^ n38474;
  assign n38852 = n38821 ^ n38712;
  assign n38848 = n37458 ^ n36070;
  assign n38849 = n37458 ^ n37435;
  assign n38850 = ~n38848 & ~n38849;
  assign n38851 = n38850 ^ n36070;
  assign n38853 = n38852 ^ n38851;
  assign n38858 = n38818 ^ n38717;
  assign n38854 = n37464 ^ n36079;
  assign n38855 = n37464 ^ n37442;
  assign n38856 = ~n38854 & ~n38855;
  assign n38857 = n38856 ^ n36079;
  assign n38859 = n38858 ^ n38857;
  assign n38864 = n38815 ^ n38812;
  assign n38860 = n37580 ^ n36086;
  assign n38861 = n37580 ^ n37449;
  assign n38862 = n38860 & n38861;
  assign n38863 = n38862 ^ n36086;
  assign n38865 = n38864 ^ n38863;
  assign n38871 = ~n38869 & ~n38870;
  assign n38872 = n38871 ^ n38864;
  assign n38873 = ~n38865 & ~n38872;
  assign n38874 = n38873 ^ n38871;
  assign n38875 = n38874 ^ n38858;
  assign n38876 = ~n38859 & n38875;
  assign n38877 = n38876 ^ n38857;
  assign n38878 = n38877 ^ n38852;
  assign n38879 = n38853 & ~n38878;
  assign n38880 = n38879 ^ n38851;
  assign n38881 = n38880 ^ n38846;
  assign n38882 = ~n38847 & n38881;
  assign n38883 = n38882 ^ n38474;
  assign n38884 = n38883 ^ n38469;
  assign n38885 = n38470 & ~n38884;
  assign n38886 = n38885 ^ n38468;
  assign n38887 = n38886 ^ n38463;
  assign n38888 = ~n38464 & ~n38887;
  assign n38889 = n38888 ^ n38462;
  assign n38458 = n38282 ^ n38269;
  assign n38890 = n38889 ^ n38458;
  assign n38891 = n37430 ^ n36860;
  assign n38892 = n38131 ^ n37430;
  assign n38893 = n38891 & n38892;
  assign n38894 = n38893 ^ n36860;
  assign n38895 = n38894 ^ n38458;
  assign n38896 = n38890 & ~n38895;
  assign n38897 = n38896 ^ n38894;
  assign n38898 = n38897 ^ n38456;
  assign n38899 = n38457 & n38898;
  assign n38900 = n38899 ^ n38455;
  assign n38901 = n38900 ^ n38449;
  assign n38902 = ~n38451 & ~n38901;
  assign n38903 = n38902 ^ n38450;
  assign n38905 = n38904 ^ n38903;
  assign n38906 = n37538 ^ n36840;
  assign n38907 = n38361 ^ n37538;
  assign n38908 = ~n38906 & n38907;
  assign n38909 = n38908 ^ n36840;
  assign n38910 = n38909 ^ n38903;
  assign n38911 = n38905 & ~n38910;
  assign n38912 = n38911 ^ n38904;
  assign n38913 = n38912 ^ n38444;
  assign n38914 = ~n38445 & ~n38913;
  assign n38915 = n38914 ^ n38443;
  assign n38916 = n38915 ^ n38432;
  assign n38917 = n38438 & ~n38916;
  assign n38918 = n38917 ^ n38437;
  assign n38919 = n38918 ^ n38425;
  assign n38920 = n38431 & ~n38919;
  assign n38921 = n38920 ^ n38430;
  assign n38922 = n38921 ^ n38418;
  assign n38923 = ~n38424 & n38922;
  assign n38924 = n38923 ^ n38423;
  assign n38925 = n38924 ^ n38411;
  assign n38926 = n38417 & ~n38925;
  assign n38927 = n38926 ^ n38416;
  assign n38928 = n38927 ^ n38404;
  assign n38929 = n38410 & n38928;
  assign n38930 = n38929 ^ n38409;
  assign n38931 = n38930 ^ n38397;
  assign n38932 = n38403 & n38931;
  assign n38933 = n38932 ^ n38402;
  assign n38934 = n38933 ^ n38390;
  assign n38935 = ~n38396 & n38934;
  assign n38936 = n38935 ^ n38395;
  assign n38937 = n38936 ^ n38383;
  assign n38938 = ~n38389 & ~n38937;
  assign n38939 = n38938 ^ n38388;
  assign n38940 = n38939 ^ n38376;
  assign n38941 = n38382 & ~n38940;
  assign n38942 = n38941 ^ n38381;
  assign n39065 = n38947 ^ n38942;
  assign n39066 = ~n38948 & n39065;
  assign n39067 = n39066 ^ n38946;
  assign n39123 = n39068 ^ n39067;
  assign n39124 = ~n39073 & ~n39123;
  assign n39125 = n39124 ^ n39072;
  assign n39323 = n39126 ^ n39125;
  assign n39324 = ~n39131 & ~n39323;
  assign n39325 = n39324 ^ n39130;
  assign n39449 = n39331 ^ n39325;
  assign n39450 = ~n39448 & ~n39449;
  assign n39451 = n39450 ^ n39329;
  assign n39447 = n38784 ^ n38749;
  assign n39452 = n39451 ^ n39447;
  assign n39453 = n37266 ^ n36576;
  assign n39454 = n38676 ^ n37266;
  assign n39455 = ~n39453 & ~n39454;
  assign n39456 = n39455 ^ n36576;
  assign n39457 = n39456 ^ n39447;
  assign n39458 = n39452 & ~n39457;
  assign n39459 = n39458 ^ n39456;
  assign n39460 = n39459 ^ n39445;
  assign n39461 = n39446 & ~n39460;
  assign n39462 = n39461 ^ n39444;
  assign n39487 = n39467 ^ n39462;
  assign n39488 = n39468 & n39487;
  assign n39489 = n39488 ^ n39466;
  assign n39494 = n39493 ^ n39489;
  assign n39496 = n39495 ^ n39494;
  assign n39497 = n39496 ^ n35790;
  assign n39469 = n39468 ^ n39462;
  assign n39470 = n39469 ^ n35797;
  assign n39471 = n39459 ^ n39446;
  assign n39472 = n39471 ^ n35803;
  assign n39476 = n39456 ^ n39452;
  assign n39330 = n39329 ^ n39325;
  assign n39332 = n39331 ^ n39330;
  assign n39333 = n39332 ^ n36544;
  assign n39132 = n39131 ^ n39125;
  assign n39133 = n39132 ^ n36355;
  assign n39074 = n39073 ^ n39067;
  assign n39075 = n39074 ^ n36256;
  assign n38949 = n38948 ^ n38942;
  assign n38950 = n38949 ^ n36110;
  assign n38951 = n38939 ^ n38382;
  assign n38952 = n38951 ^ n36116;
  assign n38953 = n38936 ^ n38389;
  assign n38954 = n38953 ^ n36126;
  assign n38955 = n38933 ^ n38396;
  assign n38956 = n38955 ^ n36133;
  assign n38957 = n38930 ^ n38403;
  assign n38958 = n38957 ^ n36140;
  assign n38959 = n38927 ^ n38410;
  assign n38960 = n38959 ^ n36146;
  assign n38961 = n38924 ^ n38417;
  assign n38962 = n38961 ^ n36152;
  assign n38963 = n38921 ^ n38423;
  assign n38964 = n38963 ^ n38418;
  assign n38965 = n38964 ^ n36220;
  assign n38966 = n38918 ^ n38430;
  assign n38967 = n38966 ^ n38425;
  assign n38968 = n38967 ^ n36159;
  assign n38969 = n38915 ^ n38437;
  assign n38970 = n38969 ^ n38432;
  assign n38971 = n38970 ^ n36165;
  assign n38972 = n38912 ^ n38443;
  assign n38973 = n38972 ^ n38444;
  assign n38974 = n38973 ^ n36062;
  assign n38975 = n38897 ^ n38455;
  assign n38976 = n38975 ^ n38456;
  assign n38977 = n38976 ^ n36065;
  assign n38978 = n38894 ^ n38890;
  assign n38979 = n38978 ^ n36074;
  assign n38980 = n38886 ^ n38462;
  assign n38981 = n38980 ^ n38463;
  assign n38982 = n38981 ^ n36054;
  assign n38983 = n38883 ^ n38470;
  assign n38984 = n38983 ^ n35922;
  assign n38985 = n38880 ^ n38847;
  assign n38986 = n38985 ^ n35852;
  assign n38987 = n38877 ^ n38851;
  assign n38988 = n38987 ^ n38852;
  assign n38989 = n38988 ^ n35111;
  assign n38990 = n38874 ^ n38859;
  assign n38991 = n38990 ^ n35119;
  assign n38993 = ~n35134 & n38992;
  assign n38994 = n38993 ^ n35132;
  assign n38995 = n38871 ^ n38863;
  assign n38996 = n38995 ^ n38864;
  assign n38997 = n38996 ^ n38993;
  assign n38998 = n38994 & ~n38997;
  assign n38999 = n38998 ^ n35132;
  assign n39000 = n38999 ^ n38990;
  assign n39001 = n38991 & n39000;
  assign n39002 = n39001 ^ n35119;
  assign n39003 = n39002 ^ n38988;
  assign n39004 = ~n38989 & n39003;
  assign n39005 = n39004 ^ n35111;
  assign n39006 = n39005 ^ n38985;
  assign n39007 = ~n38986 & ~n39006;
  assign n39008 = n39007 ^ n35852;
  assign n39009 = n39008 ^ n38983;
  assign n39010 = ~n38984 & ~n39009;
  assign n39011 = n39010 ^ n35922;
  assign n39012 = n39011 ^ n38981;
  assign n39013 = ~n38982 & ~n39012;
  assign n39014 = n39013 ^ n36054;
  assign n39015 = n39014 ^ n38978;
  assign n39016 = n38979 & ~n39015;
  assign n39017 = n39016 ^ n36074;
  assign n39018 = n39017 ^ n38976;
  assign n39019 = n38977 & n39018;
  assign n39020 = n39019 ^ n36065;
  assign n39021 = n39020 ^ n36183;
  assign n39022 = n38900 ^ n38451;
  assign n39023 = n39022 ^ n39020;
  assign n39024 = n39021 & ~n39023;
  assign n39025 = n39024 ^ n36183;
  assign n39026 = n39025 ^ n36176;
  assign n39027 = n38909 ^ n38904;
  assign n39028 = n39027 ^ n38903;
  assign n39029 = n39028 ^ n39025;
  assign n39030 = n39026 & ~n39029;
  assign n39031 = n39030 ^ n36176;
  assign n39032 = n39031 ^ n38973;
  assign n39033 = ~n38974 & n39032;
  assign n39034 = n39033 ^ n36062;
  assign n39035 = n39034 ^ n38970;
  assign n39036 = n38971 & n39035;
  assign n39037 = n39036 ^ n36165;
  assign n39038 = n39037 ^ n38967;
  assign n39039 = ~n38968 & ~n39038;
  assign n39040 = n39039 ^ n36159;
  assign n39041 = n39040 ^ n38964;
  assign n39042 = ~n38965 & ~n39041;
  assign n39043 = n39042 ^ n36220;
  assign n39044 = n39043 ^ n38961;
  assign n39045 = n38962 & ~n39044;
  assign n39046 = n39045 ^ n36152;
  assign n39047 = n39046 ^ n38959;
  assign n39048 = n38960 & ~n39047;
  assign n39049 = n39048 ^ n36146;
  assign n39050 = n39049 ^ n38957;
  assign n39051 = ~n38958 & n39050;
  assign n39052 = n39051 ^ n36140;
  assign n39053 = n39052 ^ n38955;
  assign n39054 = n38956 & n39053;
  assign n39055 = n39054 ^ n36133;
  assign n39056 = n39055 ^ n38953;
  assign n39057 = ~n38954 & ~n39056;
  assign n39058 = n39057 ^ n36126;
  assign n39059 = n39058 ^ n38951;
  assign n39060 = n38952 & n39059;
  assign n39061 = n39060 ^ n36116;
  assign n39062 = n39061 ^ n38949;
  assign n39063 = n38950 & n39062;
  assign n39064 = n39063 ^ n36110;
  assign n39120 = n39074 ^ n39064;
  assign n39121 = n39075 & ~n39120;
  assign n39122 = n39121 ^ n36256;
  assign n39320 = n39132 ^ n39122;
  assign n39321 = ~n39133 & n39320;
  assign n39322 = n39321 ^ n36355;
  assign n39473 = n39332 ^ n39322;
  assign n39474 = n39333 & ~n39473;
  assign n39475 = n39474 ^ n36544;
  assign n39477 = n39476 ^ n39475;
  assign n39478 = n39476 ^ n35806;
  assign n39479 = n39477 & n39478;
  assign n39480 = n39479 ^ n35806;
  assign n39481 = n39480 ^ n39471;
  assign n39482 = n39472 & n39481;
  assign n39483 = n39482 ^ n35803;
  assign n39484 = n39483 ^ n39469;
  assign n39485 = ~n39470 & ~n39484;
  assign n39486 = n39485 ^ n35797;
  assign n39498 = n39497 ^ n39486;
  assign n39499 = n39483 ^ n39470;
  assign n39500 = n39477 ^ n35806;
  assign n39334 = n39333 ^ n39322;
  assign n39076 = n39075 ^ n39064;
  assign n39077 = n39055 ^ n38954;
  assign n39078 = n39037 ^ n38968;
  assign n39079 = n39022 ^ n36183;
  assign n39080 = n39079 ^ n39020;
  assign n39081 = n38999 ^ n38991;
  assign n39082 = n39002 ^ n38989;
  assign n39083 = ~n39081 & ~n39082;
  assign n39084 = n39005 ^ n38986;
  assign n39085 = n39083 & ~n39084;
  assign n39086 = n39008 ^ n38984;
  assign n39087 = ~n39085 & ~n39086;
  assign n39088 = n39011 ^ n38982;
  assign n39089 = ~n39087 & ~n39088;
  assign n39090 = n39014 ^ n38979;
  assign n39091 = n39089 & ~n39090;
  assign n39092 = n39017 ^ n38977;
  assign n39093 = ~n39091 & n39092;
  assign n39094 = ~n39080 & n39093;
  assign n39095 = n39028 ^ n36176;
  assign n39096 = n39095 ^ n39025;
  assign n39097 = ~n39094 & n39096;
  assign n39098 = n39031 ^ n38974;
  assign n39099 = n39097 & ~n39098;
  assign n39100 = n39034 ^ n38971;
  assign n39101 = n39099 & n39100;
  assign n39102 = n39078 & n39101;
  assign n39103 = n39040 ^ n36220;
  assign n39104 = n39103 ^ n38964;
  assign n39105 = ~n39102 & n39104;
  assign n39106 = n39043 ^ n38962;
  assign n39107 = ~n39105 & ~n39106;
  assign n39108 = n39046 ^ n38960;
  assign n39109 = n39107 & ~n39108;
  assign n39110 = n39049 ^ n38958;
  assign n39111 = n39109 & n39110;
  assign n39112 = n39052 ^ n38956;
  assign n39113 = ~n39111 & n39112;
  assign n39114 = ~n39077 & ~n39113;
  assign n39115 = n39058 ^ n38952;
  assign n39116 = n39114 & ~n39115;
  assign n39117 = n39061 ^ n38950;
  assign n39118 = ~n39116 & ~n39117;
  assign n39119 = n39076 & n39118;
  assign n39134 = n39133 ^ n39122;
  assign n39335 = n39119 & ~n39134;
  assign n39501 = ~n39334 & ~n39335;
  assign n39502 = ~n39500 & n39501;
  assign n39503 = n39480 ^ n39472;
  assign n39504 = n39502 & n39503;
  assign n39505 = n39499 & n39504;
  assign n39506 = n39498 & ~n39505;
  assign n39514 = n37312 ^ n36554;
  assign n39515 = n38080 ^ n37312;
  assign n39516 = n39514 & ~n39515;
  assign n39517 = n39516 ^ n36554;
  assign n39510 = n39495 ^ n39493;
  assign n39511 = n39495 ^ n39489;
  assign n39512 = ~n39510 & ~n39511;
  assign n39513 = n39512 ^ n39493;
  assign n39518 = n39517 ^ n39513;
  assign n39342 = n38796 ^ n38732;
  assign n39519 = n39518 ^ n39342;
  assign n39520 = n39519 ^ n35784;
  assign n39507 = n39496 ^ n39486;
  assign n39508 = ~n39497 & n39507;
  assign n39509 = n39508 ^ n35790;
  assign n39521 = n39520 ^ n39509;
  assign n39522 = n39506 & ~n39521;
  assign n39534 = n38801 ^ n1064;
  assign n39530 = n39517 ^ n39342;
  assign n39531 = n39513 ^ n39342;
  assign n39532 = ~n39530 & ~n39531;
  assign n39533 = n39532 ^ n39517;
  assign n39535 = n39534 ^ n39533;
  assign n39526 = n37345 ^ n36104;
  assign n39527 = n38070 ^ n37345;
  assign n39528 = ~n39526 & ~n39527;
  assign n39529 = n39528 ^ n36104;
  assign n39536 = n39535 ^ n39529;
  assign n39537 = n39536 ^ n35142;
  assign n39523 = n39519 ^ n39509;
  assign n39524 = n39520 & ~n39523;
  assign n39525 = n39524 ^ n35784;
  assign n39538 = n39537 ^ n39525;
  assign n39594 = n39522 & ~n39538;
  assign n39588 = n39534 ^ n39529;
  assign n39589 = ~n39535 & n39588;
  assign n39590 = n39589 ^ n39529;
  assign n39587 = n38804 ^ n38727;
  assign n39591 = n39590 ^ n39587;
  assign n39583 = n37414 ^ n36098;
  assign n39584 = n38068 ^ n37414;
  assign n39585 = n39583 & ~n39584;
  assign n39586 = n39585 ^ n36098;
  assign n39592 = n39591 ^ n39586;
  assign n39579 = n39536 ^ n39525;
  assign n39580 = n39537 & ~n39579;
  assign n39581 = n39580 ^ n35142;
  assign n39582 = n39581 ^ n35827;
  assign n39593 = n39592 ^ n39582;
  assign n39595 = n39594 ^ n39593;
  assign n39540 = n37102 ^ n28438;
  assign n39541 = n39540 ^ n33189;
  assign n39542 = n39541 ^ n2423;
  assign n39539 = n39538 ^ n39522;
  assign n39543 = n39542 ^ n39539;
  assign n39544 = n39521 ^ n39506;
  assign n2325 = n2324 ^ n2303;
  assign n2338 = n2337 ^ n2325;
  assign n2345 = n2344 ^ n2338;
  assign n39545 = n39544 ^ n2345;
  assign n39547 = n37107 ^ n28625;
  assign n39548 = n39547 ^ n1360;
  assign n39549 = n39548 ^ n2332;
  assign n39546 = n39505 ^ n39498;
  assign n39550 = n39549 ^ n39546;
  assign n39551 = n39504 ^ n39499;
  assign n1339 = n1329 ^ n1245;
  assign n1346 = n1345 ^ n1339;
  assign n1353 = n1352 ^ n1346;
  assign n39552 = n39551 ^ n1353;
  assign n39553 = n39503 ^ n39502;
  assign n1190 = n1153 ^ n1108;
  assign n1191 = n1190 ^ n1187;
  assign n1198 = n1197 ^ n1191;
  assign n39554 = n39553 ^ n1198;
  assign n39558 = n39501 ^ n39500;
  assign n39336 = n39335 ^ n39334;
  assign n39340 = n39339 ^ n39336;
  assign n39136 = n37123 ^ n995;
  assign n39137 = n39136 ^ n33270;
  assign n39138 = n39137 ^ n27076;
  assign n39135 = n39134 ^ n39119;
  assign n39139 = n39138 ^ n39135;
  assign n39143 = n39118 ^ n39076;
  assign n39144 = n39143 ^ n39142;
  assign n39146 = n37132 ^ n28460;
  assign n39147 = n39146 ^ n33280;
  assign n39148 = n39147 ^ n725;
  assign n39145 = n39117 ^ n39116;
  assign n39149 = n39148 ^ n39145;
  assign n39303 = n39115 ^ n39114;
  assign n39151 = n37142 ^ n28470;
  assign n39152 = n39151 ^ n33250;
  assign n39153 = n39152 ^ n675;
  assign n39150 = n39113 ^ n39077;
  assign n39154 = n39153 ^ n39150;
  assign n39292 = n39112 ^ n39111;
  assign n39158 = n39110 ^ n39109;
  assign n39155 = n37186 ^ n28477;
  assign n39156 = n39155 ^ n33260;
  assign n39157 = n39156 ^ n26930;
  assign n39159 = n39158 ^ n39157;
  assign n39160 = n39108 ^ n39107;
  assign n39164 = n39163 ^ n39160;
  assign n39165 = n39106 ^ n39105;
  assign n39169 = n39168 ^ n39165;
  assign n39275 = n39104 ^ n39102;
  assign n39170 = n39101 ^ n39078;
  assign n39174 = n39173 ^ n39170;
  assign n39176 = n2237 ^ n2157;
  assign n39177 = n39176 ^ n33220;
  assign n39178 = n39177 ^ n26950;
  assign n39175 = n39100 ^ n39099;
  assign n39179 = n39178 ^ n39175;
  assign n39181 = n36685 ^ n2139;
  assign n39182 = n39181 ^ n33225;
  assign n39183 = n39182 ^ n26955;
  assign n39180 = n39098 ^ n39097;
  assign n39184 = n39183 ^ n39180;
  assign n39185 = n39096 ^ n39094;
  assign n39189 = n39188 ^ n39185;
  assign n39191 = n36753 ^ n28504;
  assign n39192 = n39191 ^ n1775;
  assign n39193 = n39192 ^ n27012;
  assign n39190 = n39093 ^ n39080;
  assign n39194 = n39193 ^ n39190;
  assign n39252 = n39092 ^ n39091;
  assign n39195 = n39090 ^ n39089;
  assign n1659 = n1658 ^ n1637;
  assign n1678 = n1677 ^ n1659;
  assign n1685 = n1684 ^ n1678;
  assign n39196 = n39195 ^ n1685;
  assign n39200 = n39088 ^ n39087;
  assign n39197 = n36701 ^ n28510;
  assign n39198 = n39197 ^ n32680;
  assign n39199 = n39198 ^ n1672;
  assign n39201 = n39200 ^ n39199;
  assign n39205 = n39086 ^ n39085;
  assign n39206 = n39205 ^ n39204;
  assign n39208 = n36733 ^ n28515;
  assign n39209 = n39208 ^ n32687;
  assign n39210 = n39209 ^ n26959;
  assign n39207 = n39084 ^ n39083;
  assign n39211 = n39210 ^ n39207;
  assign n39232 = n39082 ^ n39081;
  assign n39212 = n36720 ^ n28525;
  assign n39213 = n39212 ^ n32700;
  assign n39214 = n39213 ^ n26971;
  assign n39215 = n39214 ^ n39081;
  assign n39223 = n39221 & ~n39222;
  assign n39216 = n36715 ^ n26967;
  assign n39217 = n39216 ^ n32696;
  assign n39218 = n39217 ^ n28520;
  assign n39224 = n39223 ^ n39218;
  assign n39225 = n38996 ^ n38994;
  assign n39226 = n39225 ^ n39218;
  assign n39227 = n39224 & ~n39226;
  assign n39228 = n39227 ^ n39223;
  assign n39229 = n39228 ^ n39214;
  assign n39230 = ~n39215 & ~n39229;
  assign n39231 = n39230 ^ n39081;
  assign n39233 = n39232 ^ n39231;
  assign n39237 = n39236 ^ n39232;
  assign n39238 = ~n39233 & ~n39237;
  assign n39239 = n39238 ^ n39236;
  assign n39240 = n39239 ^ n39207;
  assign n39241 = n39211 & ~n39240;
  assign n39242 = n39241 ^ n39210;
  assign n39243 = n39242 ^ n39205;
  assign n39244 = n39206 & ~n39243;
  assign n39245 = n39244 ^ n39204;
  assign n39246 = n39245 ^ n39200;
  assign n39247 = ~n39201 & n39246;
  assign n39248 = n39247 ^ n39199;
  assign n39249 = n39248 ^ n39195;
  assign n39250 = n39196 & ~n39249;
  assign n39251 = n39250 ^ n1685;
  assign n39253 = n39252 ^ n39251;
  assign n39254 = n36694 ^ n28556;
  assign n39255 = n39254 ^ n32668;
  assign n39256 = n39255 ^ n1770;
  assign n39257 = n39256 ^ n39252;
  assign n39258 = n39253 & ~n39257;
  assign n39259 = n39258 ^ n39256;
  assign n39260 = n39259 ^ n39190;
  assign n39261 = ~n39194 & n39260;
  assign n39262 = n39261 ^ n39193;
  assign n39263 = n39262 ^ n39185;
  assign n39264 = n39189 & ~n39263;
  assign n39265 = n39264 ^ n39188;
  assign n39266 = n39265 ^ n39183;
  assign n39267 = n39184 & ~n39266;
  assign n39268 = n39267 ^ n39180;
  assign n39269 = n39268 ^ n39175;
  assign n39270 = ~n39179 & n39269;
  assign n39271 = n39270 ^ n39178;
  assign n39272 = n39271 ^ n39170;
  assign n39273 = ~n39174 & n39272;
  assign n39274 = n39273 ^ n39173;
  assign n39276 = n39275 ^ n39274;
  assign n39277 = n37157 ^ n28492;
  assign n39278 = n39277 ^ n33209;
  assign n39279 = n39278 ^ n26940;
  assign n39280 = n39279 ^ n39275;
  assign n39281 = n39276 & ~n39280;
  assign n39282 = n39281 ^ n39279;
  assign n39283 = n39282 ^ n39165;
  assign n39284 = ~n39169 & n39283;
  assign n39285 = n39284 ^ n39168;
  assign n39286 = n39285 ^ n39160;
  assign n39287 = n39164 & ~n39286;
  assign n39288 = n39287 ^ n39163;
  assign n39289 = n39288 ^ n39158;
  assign n39290 = ~n39159 & n39289;
  assign n39291 = n39290 ^ n39157;
  assign n39293 = n39292 ^ n39291;
  assign n39297 = n39296 ^ n39292;
  assign n39298 = n39293 & ~n39297;
  assign n39299 = n39298 ^ n39296;
  assign n39300 = n39299 ^ n39150;
  assign n39301 = ~n39154 & n39300;
  assign n39302 = n39301 ^ n39153;
  assign n39304 = n39303 ^ n39302;
  assign n39305 = n37137 ^ n28464;
  assign n39306 = n39305 ^ n680;
  assign n39307 = n39306 ^ n27055;
  assign n39308 = n39307 ^ n39303;
  assign n39309 = ~n39304 & n39308;
  assign n39310 = n39309 ^ n39307;
  assign n39311 = n39310 ^ n39145;
  assign n39312 = n39149 & ~n39311;
  assign n39313 = n39312 ^ n39148;
  assign n39314 = n39313 ^ n39143;
  assign n39315 = n39144 & ~n39314;
  assign n39316 = n39315 ^ n39142;
  assign n39317 = n39316 ^ n39135;
  assign n39318 = ~n39139 & n39317;
  assign n39319 = n39318 ^ n39138;
  assign n39555 = n39336 ^ n39319;
  assign n39556 = ~n39340 & n39555;
  assign n39557 = n39556 ^ n39339;
  assign n39559 = n39558 ^ n39557;
  assign n1157 = n1138 ^ n1090;
  assign n1173 = n1172 ^ n1157;
  assign n1180 = n1179 ^ n1173;
  assign n39560 = n39558 ^ n1180;
  assign n39561 = ~n39559 & n39560;
  assign n39562 = n39561 ^ n1180;
  assign n39563 = n39562 ^ n39553;
  assign n39564 = ~n39554 & n39563;
  assign n39565 = n39564 ^ n1198;
  assign n39566 = n39565 ^ n39551;
  assign n39567 = ~n39552 & n39566;
  assign n39568 = n39567 ^ n1353;
  assign n39569 = n39568 ^ n39546;
  assign n39570 = ~n39550 & n39569;
  assign n39571 = n39570 ^ n39549;
  assign n39572 = n39571 ^ n39544;
  assign n39573 = ~n39545 & n39572;
  assign n39574 = n39573 ^ n2345;
  assign n39575 = n39574 ^ n39539;
  assign n39576 = ~n39543 & n39575;
  assign n39577 = n39576 ^ n39542;
  assign n39438 = n37252 ^ n28433;
  assign n39439 = n39438 ^ n2432;
  assign n39440 = n39439 ^ n27232;
  assign n39578 = n39577 ^ n39440;
  assign n39596 = n39595 ^ n39578;
  assign n39434 = n37451 ^ n37419;
  assign n39435 = n38450 ^ n37419;
  assign n39436 = n39434 & ~n39435;
  assign n39437 = n39436 ^ n37451;
  assign n39597 = n39596 ^ n39437;
  assign n39599 = n37458 ^ n37426;
  assign n39600 = n38456 ^ n37426;
  assign n39601 = n39599 & n39600;
  assign n39602 = n39601 ^ n37458;
  assign n39598 = n39574 ^ n39543;
  assign n39603 = n39602 ^ n39598;
  assign n39608 = n39571 ^ n39545;
  assign n39604 = n37464 ^ n37428;
  assign n39605 = n38458 ^ n37428;
  assign n39606 = ~n39604 & ~n39605;
  assign n39607 = n39606 ^ n37464;
  assign n39609 = n39608 ^ n39607;
  assign n39614 = n37586 ^ n37442;
  assign n39615 = n38469 ^ n37442;
  assign n39616 = ~n39614 & n39615;
  assign n39617 = n39616 ^ n37586;
  assign n39618 = n39565 ^ n39552;
  assign n39619 = n39617 & ~n39618;
  assign n39610 = n37580 ^ n37435;
  assign n39611 = n38463 ^ n37435;
  assign n39612 = n39610 & n39611;
  assign n39613 = n39612 ^ n37580;
  assign n39620 = n39619 ^ n39613;
  assign n39621 = n39568 ^ n39550;
  assign n39622 = n39621 ^ n39613;
  assign n39623 = ~n39620 & ~n39622;
  assign n39624 = n39623 ^ n39619;
  assign n39625 = n39624 ^ n39608;
  assign n39626 = n39609 & n39625;
  assign n39627 = n39626 ^ n39607;
  assign n39628 = n39627 ^ n39598;
  assign n39629 = n39603 & ~n39628;
  assign n39630 = n39629 ^ n39602;
  assign n39631 = n39630 ^ n39596;
  assign n39632 = n39597 & ~n39631;
  assign n39633 = n39632 ^ n39437;
  assign n39634 = n39633 ^ n39428;
  assign n39635 = ~n39433 & ~n39634;
  assign n39636 = n39635 ^ n39432;
  assign n39422 = n38206 ^ n37437;
  assign n39423 = n38444 ^ n38206;
  assign n39424 = ~n39422 & n39423;
  assign n39425 = n39424 ^ n37437;
  assign n39715 = n39636 ^ n39425;
  assign n39426 = n39225 ^ n39224;
  assign n39716 = n39715 ^ n39426;
  assign n39717 = n39716 ^ n36866;
  assign n39718 = n39633 ^ n39433;
  assign n39719 = n39718 ^ n36877;
  assign n39720 = n39630 ^ n39597;
  assign n39721 = n39720 ^ n36775;
  assign n39722 = n39627 ^ n39602;
  assign n39723 = n39722 ^ n39598;
  assign n39724 = n39723 ^ n36070;
  assign n39725 = n39624 ^ n39609;
  assign n39726 = n39725 ^ n36079;
  assign n39727 = n39618 ^ n39617;
  assign n39728 = ~n36088 & ~n39727;
  assign n39729 = n39728 ^ n36086;
  assign n39730 = n39621 ^ n39620;
  assign n39731 = n39730 ^ n39728;
  assign n39732 = ~n39729 & ~n39731;
  assign n39733 = n39732 ^ n36086;
  assign n39734 = n39733 ^ n39725;
  assign n39735 = n39726 & n39734;
  assign n39736 = n39735 ^ n36079;
  assign n39737 = n39736 ^ n39723;
  assign n39738 = ~n39724 & n39737;
  assign n39739 = n39738 ^ n36070;
  assign n39740 = n39739 ^ n39720;
  assign n39741 = ~n39721 & n39740;
  assign n39742 = n39741 ^ n36775;
  assign n39743 = n39742 ^ n39718;
  assign n39744 = n39719 & ~n39743;
  assign n39745 = n39744 ^ n36877;
  assign n39746 = n39745 ^ n39716;
  assign n39747 = n39717 & n39746;
  assign n39748 = n39747 ^ n36866;
  assign n39427 = n39426 ^ n39425;
  assign n39637 = n39636 ^ n39426;
  assign n39638 = ~n39427 & ~n39637;
  assign n39639 = n39638 ^ n39425;
  assign n39420 = n39228 ^ n39215;
  assign n39416 = n38341 ^ n37430;
  assign n39417 = n38432 ^ n38341;
  assign n39418 = ~n39416 & ~n39417;
  assign n39419 = n39418 ^ n37430;
  assign n39421 = n39420 ^ n39419;
  assign n39713 = n39639 ^ n39421;
  assign n39714 = n39713 ^ n36860;
  assign n39819 = n39748 ^ n39714;
  assign n39810 = n39745 ^ n39717;
  assign n39811 = n39742 ^ n39719;
  assign n39812 = n39739 ^ n39721;
  assign n39813 = n39733 ^ n39726;
  assign n39814 = n39736 ^ n39724;
  assign n39815 = n39813 & n39814;
  assign n39816 = n39812 & n39815;
  assign n39817 = n39811 & ~n39816;
  assign n39818 = ~n39810 & ~n39817;
  assign n39892 = n39819 ^ n39818;
  assign n39893 = n39892 ^ n39891;
  assign n39894 = n39817 ^ n39810;
  assign n39898 = n39897 ^ n39894;
  assign n39899 = n39816 ^ n39811;
  assign n39903 = n39902 ^ n39899;
  assign n39905 = n37369 ^ n28803;
  assign n39906 = n39905 ^ n33683;
  assign n39907 = n39906 ^ n27197;
  assign n39904 = n39815 ^ n39812;
  assign n39908 = n39907 ^ n39904;
  assign n39929 = n39814 ^ n39813;
  assign n39909 = n37379 ^ n28816;
  assign n39910 = n39909 ^ n33696;
  assign n39911 = n39910 ^ n27119;
  assign n39912 = n39911 ^ n39813;
  assign n39918 = n33691 ^ n28811;
  assign n39919 = n39918 ^ n2579;
  assign n39920 = n39919 ^ n2636;
  assign n39913 = n38048 ^ n29449;
  assign n39914 = n39913 ^ n2542;
  assign n39915 = n39914 ^ n28042;
  assign n39916 = n39727 ^ n36088;
  assign n39917 = n39915 & n39916;
  assign n39921 = n39920 ^ n39917;
  assign n39922 = n39730 ^ n39729;
  assign n39923 = n39922 ^ n39920;
  assign n39924 = n39921 & n39923;
  assign n39925 = n39924 ^ n39917;
  assign n39926 = n39925 ^ n39813;
  assign n39927 = n39912 & ~n39926;
  assign n39928 = n39927 ^ n39911;
  assign n39930 = n39929 ^ n39928;
  assign n39931 = n37373 ^ n28807;
  assign n39932 = n39931 ^ n33687;
  assign n39933 = n39932 ^ n1559;
  assign n39934 = n39933 ^ n39929;
  assign n39935 = n39930 & ~n39934;
  assign n39936 = n39935 ^ n39933;
  assign n39937 = n39936 ^ n39904;
  assign n39938 = ~n39908 & n39937;
  assign n39939 = n39938 ^ n39907;
  assign n39940 = n39939 ^ n39899;
  assign n39941 = ~n39903 & n39940;
  assign n39942 = n39941 ^ n39902;
  assign n39943 = n39942 ^ n39894;
  assign n39944 = ~n39898 & n39943;
  assign n39945 = n39944 ^ n39897;
  assign n39946 = n39945 ^ n39892;
  assign n39947 = ~n39893 & n39946;
  assign n39948 = n39947 ^ n39891;
  assign n39820 = n39818 & n39819;
  assign n39749 = n39748 ^ n39713;
  assign n39750 = n39714 & ~n39749;
  assign n39751 = n39750 ^ n36860;
  assign n39640 = n39639 ^ n39420;
  assign n39641 = n39421 & ~n39640;
  assign n39642 = n39641 ^ n39419;
  assign n39411 = n38361 ^ n37422;
  assign n39412 = n38425 ^ n38361;
  assign n39413 = n39411 & n39412;
  assign n39414 = n39413 ^ n37422;
  assign n39710 = n39642 ^ n39414;
  assign n39410 = n39236 ^ n39233;
  assign n39711 = n39710 ^ n39410;
  assign n39712 = n39711 ^ n36853;
  assign n39809 = n39751 ^ n39712;
  assign n39887 = n39820 ^ n39809;
  assign n39884 = n37949 ^ n1744;
  assign n39885 = n39884 ^ n33662;
  assign n39886 = n39885 ^ n1865;
  assign n39888 = n39887 ^ n39886;
  assign n40038 = n39948 ^ n39888;
  assign n39380 = n39256 ^ n39253;
  assign n41679 = n40038 ^ n39380;
  assign n40239 = n29264 ^ n1397;
  assign n40240 = n40239 ^ n34142;
  assign n40241 = n40240 ^ n28011;
  assign n40114 = n39307 ^ n39304;
  assign n40110 = n38086 ^ n37266;
  assign n40111 = n39534 ^ n38086;
  assign n40112 = ~n40110 & n40111;
  assign n40113 = n40112 ^ n37266;
  assign n40115 = n40114 ^ n40113;
  assign n40120 = n39299 ^ n39154;
  assign n40116 = n38833 ^ n38062;
  assign n40117 = n39342 ^ n38833;
  assign n40118 = ~n40116 & n40117;
  assign n40119 = n40118 ^ n38062;
  assign n40121 = n40120 ^ n40119;
  assign n40123 = n38676 ^ n37804;
  assign n40124 = n39495 ^ n38676;
  assign n40125 = ~n40123 & ~n40124;
  assign n40126 = n40125 ^ n37804;
  assign n40122 = n39296 ^ n39293;
  assign n40127 = n40126 ^ n40122;
  assign n40018 = n39288 ^ n39159;
  assign n39798 = n39285 ^ n39164;
  assign n39683 = n39282 ^ n39169;
  assign n39679 = n38492 ^ n37479;
  assign n39680 = n39447 ^ n38492;
  assign n39681 = ~n39679 & ~n39680;
  assign n39682 = n39681 ^ n37479;
  assign n39684 = n39683 ^ n39682;
  assign n39348 = n39279 ^ n39276;
  assign n39344 = n38498 ^ n37489;
  assign n39345 = n39331 ^ n38498;
  assign n39346 = n39344 & ~n39345;
  assign n39347 = n39346 ^ n37489;
  assign n39349 = n39348 ^ n39347;
  assign n39354 = n39271 ^ n39174;
  assign n39350 = n38378 ^ n37491;
  assign n39351 = n39126 ^ n38378;
  assign n39352 = n39350 & n39351;
  assign n39353 = n39352 ^ n37491;
  assign n39355 = n39354 ^ n39353;
  assign n39360 = n39268 ^ n39179;
  assign n39356 = n38385 ^ n37497;
  assign n39357 = n39068 ^ n38385;
  assign n39358 = n39356 & n39357;
  assign n39359 = n39358 ^ n37497;
  assign n39361 = n39360 ^ n39359;
  assign n39363 = n38392 ^ n37503;
  assign n39364 = n38947 ^ n38392;
  assign n39365 = n39363 & ~n39364;
  assign n39366 = n39365 ^ n37503;
  assign n39362 = n39265 ^ n39184;
  assign n39367 = n39366 ^ n39362;
  assign n39372 = n39262 ^ n39189;
  assign n39368 = n38399 ^ n37509;
  assign n39369 = n38399 ^ n38376;
  assign n39370 = n39368 & n39369;
  assign n39371 = n39370 ^ n37509;
  assign n39373 = n39372 ^ n39371;
  assign n39375 = n38406 ^ n37510;
  assign n39376 = n38406 ^ n38383;
  assign n39377 = n39375 & n39376;
  assign n39378 = n39377 ^ n37510;
  assign n39374 = n39259 ^ n39194;
  assign n39379 = n39378 ^ n39374;
  assign n39381 = n38413 ^ n37516;
  assign n39382 = n38413 ^ n38390;
  assign n39383 = n39381 & n39382;
  assign n39384 = n39383 ^ n37516;
  assign n39385 = n39384 ^ n39380;
  assign n39387 = n38420 ^ n37526;
  assign n39388 = n38420 ^ n38397;
  assign n39389 = ~n39387 & n39388;
  assign n39390 = n39389 ^ n37526;
  assign n39386 = n39248 ^ n39196;
  assign n39391 = n39390 ^ n39386;
  assign n39393 = n38427 ^ n37532;
  assign n39394 = n38427 ^ n38404;
  assign n39395 = ~n39393 & ~n39394;
  assign n39396 = n39395 ^ n37532;
  assign n39392 = n39245 ^ n39201;
  assign n39397 = n39396 ^ n39392;
  assign n39399 = n38434 ^ n37538;
  assign n39400 = n38434 ^ n38411;
  assign n39401 = n39399 & ~n39400;
  assign n39402 = n39401 ^ n37538;
  assign n39398 = n39242 ^ n39206;
  assign n39403 = n39402 ^ n39398;
  assign n39405 = n38440 ^ n36782;
  assign n39406 = n38440 ^ n38418;
  assign n39407 = n39405 & ~n39406;
  assign n39408 = n39407 ^ n36782;
  assign n39404 = n39239 ^ n39211;
  assign n39409 = n39408 ^ n39404;
  assign n39415 = n39414 ^ n39410;
  assign n39643 = n39642 ^ n39410;
  assign n39644 = ~n39415 & n39643;
  assign n39645 = n39644 ^ n39414;
  assign n39646 = n39645 ^ n39404;
  assign n39647 = ~n39409 & n39646;
  assign n39648 = n39647 ^ n39408;
  assign n39649 = n39648 ^ n39398;
  assign n39650 = n39403 & n39649;
  assign n39651 = n39650 ^ n39402;
  assign n39652 = n39651 ^ n39392;
  assign n39653 = ~n39397 & n39652;
  assign n39654 = n39653 ^ n39396;
  assign n39655 = n39654 ^ n39386;
  assign n39656 = n39391 & ~n39655;
  assign n39657 = n39656 ^ n39390;
  assign n39658 = n39657 ^ n39380;
  assign n39659 = ~n39385 & n39658;
  assign n39660 = n39659 ^ n39384;
  assign n39661 = n39660 ^ n39374;
  assign n39662 = n39379 & n39661;
  assign n39663 = n39662 ^ n39378;
  assign n39664 = n39663 ^ n39372;
  assign n39665 = n39373 & n39664;
  assign n39666 = n39665 ^ n39371;
  assign n39667 = n39666 ^ n39362;
  assign n39668 = n39367 & ~n39667;
  assign n39669 = n39668 ^ n39366;
  assign n39670 = n39669 ^ n39360;
  assign n39671 = ~n39361 & n39670;
  assign n39672 = n39671 ^ n39359;
  assign n39673 = n39672 ^ n39354;
  assign n39674 = n39355 & n39673;
  assign n39675 = n39674 ^ n39353;
  assign n39676 = n39675 ^ n39348;
  assign n39677 = n39349 & ~n39676;
  assign n39678 = n39677 ^ n39347;
  assign n39795 = n39683 ^ n39678;
  assign n39796 = ~n39684 & ~n39795;
  assign n39797 = n39796 ^ n39682;
  assign n39799 = n39798 ^ n39797;
  assign n39791 = n38486 ^ n37473;
  assign n39792 = n39445 ^ n38486;
  assign n39793 = ~n39791 & n39792;
  assign n39794 = n39793 ^ n37473;
  assign n40015 = n39798 ^ n39794;
  assign n40016 = ~n39799 & n40015;
  assign n40017 = n40016 ^ n39794;
  assign n40019 = n40018 ^ n40017;
  assign n40011 = n38592 ^ n37472;
  assign n40012 = n39467 ^ n38592;
  assign n40013 = ~n40011 & ~n40012;
  assign n40014 = n40013 ^ n37472;
  assign n40128 = n40018 ^ n40014;
  assign n40129 = n40019 & ~n40128;
  assign n40130 = n40129 ^ n40014;
  assign n40131 = n40130 ^ n40122;
  assign n40132 = ~n40127 & n40131;
  assign n40133 = n40132 ^ n40126;
  assign n40134 = n40133 ^ n40120;
  assign n40135 = ~n40121 & n40134;
  assign n40136 = n40135 ^ n40119;
  assign n40137 = n40136 ^ n40114;
  assign n40138 = ~n40115 & ~n40137;
  assign n40139 = n40138 ^ n40113;
  assign n40104 = n38093 ^ n37273;
  assign n40105 = n39587 ^ n38093;
  assign n40106 = n40104 & n40105;
  assign n40107 = n40106 ^ n37273;
  assign n40162 = n40139 ^ n40107;
  assign n40108 = n39310 ^ n39149;
  assign n40163 = n40162 ^ n40108;
  assign n40164 = n40163 ^ n36573;
  assign n40165 = n40136 ^ n40113;
  assign n40166 = n40165 ^ n40114;
  assign n40167 = n40166 ^ n36576;
  assign n40168 = n40133 ^ n40119;
  assign n40169 = n40168 ^ n40120;
  assign n40170 = n40169 ^ n37307;
  assign n40171 = n40130 ^ n40126;
  assign n40172 = n40171 ^ n40122;
  assign n40173 = n40172 ^ n37244;
  assign n40020 = n40019 ^ n40014;
  assign n40174 = n40020 ^ n37096;
  assign n39800 = n39799 ^ n39794;
  assign n39801 = n39800 ^ n37077;
  assign n39685 = n39684 ^ n39678;
  assign n39686 = n39685 ^ n37021;
  assign n39687 = n39675 ^ n39349;
  assign n39688 = n39687 ^ n36929;
  assign n39689 = n39672 ^ n39355;
  assign n39690 = n39689 ^ n36795;
  assign n39691 = n39669 ^ n39361;
  assign n39692 = n39691 ^ n36802;
  assign n39693 = n39666 ^ n39367;
  assign n39694 = n39693 ^ n36808;
  assign n39695 = n39663 ^ n39373;
  assign n39696 = n39695 ^ n36810;
  assign n39697 = n39660 ^ n39379;
  assign n39698 = n39697 ^ n36816;
  assign n39699 = n39657 ^ n39385;
  assign n39700 = n39699 ^ n36823;
  assign n39701 = n39654 ^ n39390;
  assign n39702 = n39701 ^ n39386;
  assign n39703 = n39702 ^ n36833;
  assign n39704 = n39651 ^ n39397;
  assign n39705 = n39704 ^ n36060;
  assign n39706 = n39648 ^ n39403;
  assign n39707 = n39706 ^ n36840;
  assign n39708 = n39645 ^ n39409;
  assign n39709 = n39708 ^ n36847;
  assign n39752 = n39751 ^ n39711;
  assign n39753 = n39712 & n39752;
  assign n39754 = n39753 ^ n36853;
  assign n39755 = n39754 ^ n39708;
  assign n39756 = n39709 & ~n39755;
  assign n39757 = n39756 ^ n36847;
  assign n39758 = n39757 ^ n39706;
  assign n39759 = n39707 & n39758;
  assign n39760 = n39759 ^ n36840;
  assign n39761 = n39760 ^ n39704;
  assign n39762 = ~n39705 & ~n39761;
  assign n39763 = n39762 ^ n36060;
  assign n39764 = n39763 ^ n39702;
  assign n39765 = n39703 & ~n39764;
  assign n39766 = n39765 ^ n36833;
  assign n39767 = n39766 ^ n39699;
  assign n39768 = ~n39700 & n39767;
  assign n39769 = n39768 ^ n36823;
  assign n39770 = n39769 ^ n39697;
  assign n39771 = n39698 & ~n39770;
  assign n39772 = n39771 ^ n36816;
  assign n39773 = n39772 ^ n39695;
  assign n39774 = ~n39696 & n39773;
  assign n39775 = n39774 ^ n36810;
  assign n39776 = n39775 ^ n39693;
  assign n39777 = ~n39694 & ~n39776;
  assign n39778 = n39777 ^ n36808;
  assign n39779 = n39778 ^ n39691;
  assign n39780 = ~n39692 & ~n39779;
  assign n39781 = n39780 ^ n36802;
  assign n39782 = n39781 ^ n39689;
  assign n39783 = n39690 & ~n39782;
  assign n39784 = n39783 ^ n36795;
  assign n39785 = n39784 ^ n39687;
  assign n39786 = n39688 & n39785;
  assign n39787 = n39786 ^ n36929;
  assign n39788 = n39787 ^ n39685;
  assign n39789 = ~n39686 & n39788;
  assign n39790 = n39789 ^ n37021;
  assign n40007 = n39800 ^ n39790;
  assign n40008 = ~n39801 & n40007;
  assign n40009 = n40008 ^ n37077;
  assign n40175 = n40020 ^ n40009;
  assign n40176 = ~n40174 & ~n40175;
  assign n40177 = n40176 ^ n37096;
  assign n40178 = n40177 ^ n40172;
  assign n40179 = n40173 & n40178;
  assign n40180 = n40179 ^ n37244;
  assign n40181 = n40180 ^ n40169;
  assign n40182 = ~n40170 & ~n40181;
  assign n40183 = n40182 ^ n37307;
  assign n40184 = n40183 ^ n40166;
  assign n40185 = ~n40167 & n40184;
  assign n40186 = n40185 ^ n36576;
  assign n40187 = n40186 ^ n40163;
  assign n40188 = ~n40164 & n40187;
  assign n40189 = n40188 ^ n36573;
  assign n40109 = n40108 ^ n40107;
  assign n40140 = n40139 ^ n40108;
  assign n40141 = n40109 & n40140;
  assign n40142 = n40141 ^ n40107;
  assign n40098 = n38080 ^ n37260;
  assign n40099 = n38870 ^ n38080;
  assign n40100 = ~n40098 & ~n40099;
  assign n40101 = n40100 ^ n37260;
  assign n40159 = n40142 ^ n40101;
  assign n40102 = n39313 ^ n39144;
  assign n40160 = n40159 ^ n40102;
  assign n40161 = n40160 ^ n36567;
  assign n40213 = n40189 ^ n40161;
  assign n40214 = n40180 ^ n40170;
  assign n39802 = n39801 ^ n39790;
  assign n39803 = n39781 ^ n39690;
  assign n39804 = n39778 ^ n39692;
  assign n39805 = n39775 ^ n39694;
  assign n39806 = n39769 ^ n39698;
  assign n39807 = n39766 ^ n39700;
  assign n39808 = n39763 ^ n39703;
  assign n39821 = ~n39809 & ~n39820;
  assign n39822 = n39754 ^ n39709;
  assign n39823 = n39821 & n39822;
  assign n39824 = n39757 ^ n39707;
  assign n39825 = ~n39823 & ~n39824;
  assign n39826 = n39760 ^ n39705;
  assign n39827 = n39825 & ~n39826;
  assign n39828 = ~n39808 & n39827;
  assign n39829 = n39807 & n39828;
  assign n39830 = n39806 & ~n39829;
  assign n39831 = n39772 ^ n39696;
  assign n39832 = ~n39830 & n39831;
  assign n39833 = n39805 & n39832;
  assign n39834 = ~n39804 & n39833;
  assign n39835 = n39803 & ~n39834;
  assign n39836 = n39784 ^ n39688;
  assign n39837 = ~n39835 & ~n39836;
  assign n39838 = n39787 ^ n39686;
  assign n39839 = n39837 & ~n39838;
  assign n40006 = n39802 & ~n39839;
  assign n40010 = n40009 ^ n37096;
  assign n40021 = n40020 ^ n40010;
  assign n40215 = n40006 & n40021;
  assign n40216 = n40177 ^ n37244;
  assign n40217 = n40216 ^ n40172;
  assign n40218 = n40215 & n40217;
  assign n40219 = ~n40214 & ~n40218;
  assign n40220 = n40183 ^ n40167;
  assign n40221 = n40219 & n40220;
  assign n40222 = n40186 ^ n40164;
  assign n40223 = n40221 & n40222;
  assign n40224 = n40213 & n40223;
  assign n40190 = n40189 ^ n40160;
  assign n40191 = ~n40161 & ~n40190;
  assign n40192 = n40191 ^ n36567;
  assign n40103 = n40102 ^ n40101;
  assign n40143 = n40142 ^ n40102;
  assign n40144 = n40103 & ~n40143;
  assign n40145 = n40144 ^ n40101;
  assign n40092 = n38070 ^ n37254;
  assign n40093 = n38864 ^ n38070;
  assign n40094 = ~n40092 & n40093;
  assign n40095 = n40094 ^ n37254;
  assign n40156 = n40145 ^ n40095;
  assign n40096 = n39316 ^ n39139;
  assign n40157 = n40156 ^ n40096;
  assign n40158 = n40157 ^ n36560;
  assign n40212 = n40192 ^ n40158;
  assign n40238 = n40224 ^ n40212;
  assign n40242 = n40241 ^ n40238;
  assign n40278 = n40223 ^ n40213;
  assign n40246 = n40222 ^ n40221;
  assign n40243 = n38027 ^ n1281;
  assign n40244 = n40243 ^ n34221;
  assign n40245 = n40244 ^ n27983;
  assign n40247 = n40246 ^ n40245;
  assign n40267 = n40220 ^ n40219;
  assign n40251 = n40218 ^ n40214;
  assign n40252 = n40251 ^ n40250;
  assign n40256 = n40217 ^ n40215;
  assign n40022 = n40021 ^ n40006;
  assign n774 = n773 ^ n752;
  assign n802 = n801 ^ n774;
  assign n809 = n808 ^ n802;
  assign n40023 = n40022 ^ n809;
  assign n39841 = n37905 ^ n29282;
  assign n39842 = n39841 ^ n34154;
  assign n39843 = n39842 ^ n793;
  assign n39840 = n39839 ^ n39802;
  assign n39844 = n39843 ^ n39840;
  assign n39995 = n39838 ^ n39837;
  assign n39846 = n37915 ^ n29289;
  assign n39847 = n39846 ^ n34159;
  assign n39848 = n39847 ^ n27584;
  assign n39845 = n39836 ^ n39835;
  assign n39849 = n39848 ^ n39845;
  assign n39984 = n39834 ^ n39803;
  assign n39851 = n37925 ^ n29299;
  assign n39852 = n39851 ^ n33634;
  assign n39853 = n39852 ^ n27594;
  assign n39850 = n39833 ^ n39804;
  assign n39854 = n39853 ^ n39850;
  assign n39858 = n39832 ^ n39805;
  assign n39855 = n37929 ^ n29304;
  assign n39856 = n39855 ^ n33639;
  assign n39857 = n39856 ^ n27599;
  assign n39859 = n39858 ^ n39857;
  assign n39860 = n39831 ^ n39830;
  assign n39864 = n39863 ^ n39860;
  assign n39865 = n39829 ^ n39806;
  assign n39869 = n39868 ^ n39865;
  assign n39871 = n37978 ^ n29319;
  assign n39872 = n39871 ^ n2192;
  assign n39873 = n39872 ^ n27609;
  assign n39870 = n39828 ^ n39807;
  assign n39874 = n39873 ^ n39870;
  assign n39961 = n39827 ^ n39808;
  assign n39875 = n39826 ^ n39825;
  assign n1998 = n1997 ^ n1931;
  assign n2014 = n2013 ^ n1998;
  assign n2021 = n2020 ^ n2014;
  assign n39876 = n39875 ^ n2021;
  assign n39880 = n39824 ^ n39823;
  assign n39881 = n39880 ^ n39879;
  assign n39882 = n39822 ^ n39821;
  assign n1849 = n1839 ^ n1803;
  assign n1874 = n1873 ^ n1849;
  assign n1881 = n1880 ^ n1874;
  assign n39883 = n39882 ^ n1881;
  assign n39949 = n39948 ^ n39887;
  assign n39950 = n39888 & ~n39949;
  assign n39951 = n39950 ^ n39886;
  assign n39952 = n39951 ^ n39882;
  assign n39953 = n39883 & ~n39952;
  assign n39954 = n39953 ^ n1881;
  assign n39955 = n39954 ^ n39880;
  assign n39956 = ~n39881 & n39955;
  assign n39957 = n39956 ^ n39879;
  assign n39958 = n39957 ^ n39875;
  assign n39959 = n39876 & ~n39958;
  assign n39960 = n39959 ^ n2021;
  assign n39962 = n39961 ^ n39960;
  assign n39966 = n39965 ^ n39961;
  assign n39967 = ~n39962 & n39966;
  assign n39968 = n39967 ^ n39965;
  assign n39969 = n39968 ^ n39870;
  assign n39970 = ~n39874 & n39969;
  assign n39971 = n39970 ^ n39873;
  assign n39972 = n39971 ^ n39865;
  assign n39973 = ~n39869 & n39972;
  assign n39974 = n39973 ^ n39868;
  assign n39975 = n39974 ^ n39860;
  assign n39976 = n39864 & ~n39975;
  assign n39977 = n39976 ^ n39863;
  assign n39978 = n39977 ^ n39858;
  assign n39979 = ~n39859 & n39978;
  assign n39980 = n39979 ^ n39857;
  assign n39981 = n39980 ^ n39850;
  assign n39982 = n39854 & ~n39981;
  assign n39983 = n39982 ^ n39853;
  assign n39985 = n39984 ^ n39983;
  assign n39986 = n37920 ^ n29294;
  assign n39987 = n39986 ^ n33775;
  assign n39988 = n39987 ^ n27589;
  assign n39989 = n39988 ^ n39984;
  assign n39990 = n39985 & ~n39989;
  assign n39991 = n39990 ^ n39988;
  assign n39992 = n39991 ^ n39845;
  assign n39993 = ~n39849 & n39992;
  assign n39994 = n39993 ^ n39848;
  assign n39996 = n39995 ^ n39994;
  assign n39997 = n37910 ^ n699;
  assign n39998 = n39997 ^ n34167;
  assign n39999 = n39998 ^ n27579;
  assign n40000 = n39999 ^ n39995;
  assign n40001 = ~n39996 & n40000;
  assign n40002 = n40001 ^ n39999;
  assign n40003 = n40002 ^ n39840;
  assign n40004 = ~n39844 & n40003;
  assign n40005 = n40004 ^ n39843;
  assign n40253 = n40022 ^ n40005;
  assign n40254 = n40023 & ~n40253;
  assign n40255 = n40254 ^ n809;
  assign n40257 = n40256 ^ n40255;
  assign n40258 = n37898 ^ n29371;
  assign n40259 = n40258 ^ n34174;
  assign n40260 = n40259 ^ n887;
  assign n40261 = n40260 ^ n40256;
  assign n40262 = ~n40257 & n40261;
  assign n40263 = n40262 ^ n40260;
  assign n40264 = n40263 ^ n40251;
  assign n40265 = ~n40252 & n40264;
  assign n40266 = n40265 ^ n40250;
  assign n40268 = n40267 ^ n40266;
  assign n40272 = n40271 ^ n40267;
  assign n40273 = n40268 & ~n40272;
  assign n40274 = n40273 ^ n40271;
  assign n40275 = n40274 ^ n40246;
  assign n40276 = ~n40247 & n40275;
  assign n40277 = n40276 ^ n40245;
  assign n40279 = n40278 ^ n40277;
  assign n40280 = n1382 ^ n1299;
  assign n40281 = n40280 ^ n34147;
  assign n40282 = n40281 ^ n27978;
  assign n40283 = n40282 ^ n40278;
  assign n40284 = n40279 & ~n40283;
  assign n40285 = n40284 ^ n40282;
  assign n40286 = n40285 ^ n40238;
  assign n40287 = n40242 & ~n40286;
  assign n40288 = n40287 ^ n40241;
  assign n40193 = n40192 ^ n40157;
  assign n40194 = n40158 & n40193;
  assign n40195 = n40194 ^ n36560;
  assign n40149 = n38068 ^ n37312;
  assign n40150 = n38858 ^ n38068;
  assign n40151 = ~n40149 & n40150;
  assign n40152 = n40151 ^ n37312;
  assign n40097 = n40096 ^ n40095;
  assign n40146 = n40145 ^ n40096;
  assign n40147 = n40097 & n40146;
  assign n40148 = n40147 ^ n40095;
  assign n40153 = n40152 ^ n40148;
  assign n39341 = n39340 ^ n39319;
  assign n40154 = n40153 ^ n39341;
  assign n40155 = n40154 ^ n36554;
  assign n40226 = n40195 ^ n40155;
  assign n40225 = ~n40212 & ~n40224;
  assign n40236 = n40226 ^ n40225;
  assign n40233 = n37878 ^ n2389;
  assign n40234 = n40233 ^ n34136;
  assign n40235 = n40234 ^ n27973;
  assign n40237 = n40236 ^ n40235;
  assign n40326 = n40288 ^ n40237;
  assign n40322 = n38450 ^ n37428;
  assign n40323 = n39420 ^ n38450;
  assign n40324 = ~n40322 & ~n40323;
  assign n40325 = n40324 ^ n37428;
  assign n40327 = n40326 ^ n40325;
  assign n40332 = n40285 ^ n40242;
  assign n40328 = n38456 ^ n37435;
  assign n40329 = n39426 ^ n38456;
  assign n40330 = ~n40328 & ~n40329;
  assign n40331 = n40330 ^ n37435;
  assign n40333 = n40332 ^ n40331;
  assign n40334 = n38458 ^ n37442;
  assign n40335 = n39428 ^ n38458;
  assign n40336 = ~n40334 & n40335;
  assign n40337 = n40336 ^ n37442;
  assign n40338 = n40282 ^ n40279;
  assign n40339 = ~n40337 & ~n40338;
  assign n40340 = n40339 ^ n40332;
  assign n40341 = n40333 & n40340;
  assign n40342 = n40341 ^ n40339;
  assign n40343 = n40342 ^ n40326;
  assign n40344 = n40327 & ~n40343;
  assign n40345 = n40344 ^ n40325;
  assign n40316 = n38904 ^ n37426;
  assign n40317 = n39410 ^ n38904;
  assign n40318 = n40316 & n40317;
  assign n40319 = n40318 ^ n37426;
  assign n40412 = n40345 ^ n40319;
  assign n40289 = n40288 ^ n40236;
  assign n40290 = n40237 & ~n40289;
  assign n40291 = n40290 ^ n40235;
  assign n40229 = n37874 ^ n2404;
  assign n40230 = n40229 ^ n34132;
  assign n40231 = n40230 ^ n2516;
  assign n40227 = n40225 & n40226;
  assign n40208 = n39559 ^ n1180;
  assign n40203 = n37456 ^ n37345;
  assign n40204 = n38852 ^ n37456;
  assign n40205 = ~n40203 & n40204;
  assign n40206 = n40205 ^ n37345;
  assign n40199 = n40152 ^ n39341;
  assign n40200 = n40148 ^ n39341;
  assign n40201 = n40199 & ~n40200;
  assign n40202 = n40201 ^ n40152;
  assign n40207 = n40206 ^ n40202;
  assign n40209 = n40208 ^ n40207;
  assign n40210 = n40209 ^ n36104;
  assign n40196 = n40195 ^ n40154;
  assign n40197 = n40155 & n40196;
  assign n40198 = n40197 ^ n36554;
  assign n40211 = n40210 ^ n40198;
  assign n40228 = n40227 ^ n40211;
  assign n40232 = n40231 ^ n40228;
  assign n40320 = n40291 ^ n40232;
  assign n40413 = n40412 ^ n40320;
  assign n40414 = n40413 ^ n37458;
  assign n40415 = n40342 ^ n40327;
  assign n40416 = n40415 ^ n37464;
  assign n40417 = n40338 ^ n40337;
  assign n40418 = n37586 & n40417;
  assign n40419 = n40418 ^ n37580;
  assign n40420 = n40339 ^ n40331;
  assign n40421 = n40420 ^ n40332;
  assign n40422 = n40421 ^ n40418;
  assign n40423 = ~n40419 & n40422;
  assign n40424 = n40423 ^ n37580;
  assign n40425 = n40424 ^ n40415;
  assign n40426 = ~n40416 & n40425;
  assign n40427 = n40426 ^ n37464;
  assign n40428 = n40427 ^ n40413;
  assign n40429 = ~n40414 & n40428;
  assign n40430 = n40429 ^ n37458;
  assign n40321 = n40320 ^ n40319;
  assign n40346 = n40345 ^ n40320;
  assign n40347 = n40321 & n40346;
  assign n40348 = n40347 ^ n40319;
  assign n40312 = ~n40211 & n40227;
  assign n40304 = n37449 ^ n37414;
  assign n40305 = n38846 ^ n37449;
  assign n40306 = n40304 & n40305;
  assign n40307 = n40306 ^ n37414;
  assign n40303 = n39562 ^ n39554;
  assign n40308 = n40307 ^ n40303;
  assign n40299 = n40208 ^ n40206;
  assign n40300 = n40208 ^ n40202;
  assign n40301 = n40299 & n40300;
  assign n40302 = n40301 ^ n40206;
  assign n40309 = n40308 ^ n40302;
  assign n40310 = n40309 ^ n36098;
  assign n40296 = n40209 ^ n40198;
  assign n40297 = n40210 & ~n40296;
  assign n40298 = n40297 ^ n36104;
  assign n40311 = n40310 ^ n40298;
  assign n40313 = n40312 ^ n40311;
  assign n40292 = n40291 ^ n40228;
  assign n40293 = ~n40232 & n40292;
  assign n40294 = n40293 ^ n40231;
  assign n2503 = n2499 ^ n2460;
  assign n2525 = n2524 ^ n2503;
  assign n2532 = n2531 ^ n2525;
  assign n40295 = n40294 ^ n2532;
  assign n40314 = n40313 ^ n40295;
  assign n40088 = n38444 ^ n37419;
  assign n40089 = n39404 ^ n38444;
  assign n40090 = n40088 & n40089;
  assign n40091 = n40090 ^ n37419;
  assign n40315 = n40314 ^ n40091;
  assign n40410 = n40348 ^ n40315;
  assign n40411 = n40410 ^ n37451;
  assign n40488 = n40430 ^ n40411;
  assign n40489 = n40424 ^ n40416;
  assign n40490 = n40427 ^ n40414;
  assign n40491 = ~n40489 & ~n40490;
  assign n40492 = n40488 & n40491;
  assign n40431 = n40430 ^ n40410;
  assign n40432 = n40411 & ~n40431;
  assign n40433 = n40432 ^ n37451;
  assign n40349 = n40348 ^ n40314;
  assign n40350 = n40315 & ~n40349;
  assign n40351 = n40350 ^ n40091;
  assign n40083 = n38432 ^ n38131;
  assign n40084 = n39398 ^ n38432;
  assign n40085 = n40083 & ~n40084;
  assign n40086 = n40085 ^ n38131;
  assign n40082 = n39916 ^ n39915;
  assign n40087 = n40086 ^ n40082;
  assign n40408 = n40351 ^ n40087;
  assign n40409 = n40408 ^ n37444;
  assign n40487 = n40433 ^ n40409;
  assign n40549 = n40492 ^ n40487;
  assign n40546 = n38263 ^ n29666;
  assign n40547 = n40546 ^ n34753;
  assign n40548 = n40547 ^ n1584;
  assign n40550 = n40549 ^ n40548;
  assign n40554 = n40491 ^ n40488;
  assign n40551 = n38290 ^ n1562;
  assign n40552 = n40551 ^ n34758;
  assign n40553 = n40552 ^ n28515;
  assign n40555 = n40554 ^ n40553;
  assign n40576 = n40490 ^ n40489;
  assign n40559 = n40558 ^ n40489;
  assign n40563 = n38827 ^ n2609;
  assign n40564 = n40563 ^ n35028;
  assign n40565 = n40564 ^ n28640;
  assign n40566 = n40417 ^ n37586;
  assign n40567 = n40565 & n40566;
  assign n40560 = n38272 ^ n29674;
  assign n40561 = n40560 ^ n34767;
  assign n40562 = n40561 ^ n28520;
  assign n40568 = n40567 ^ n40562;
  assign n40569 = n40421 ^ n40419;
  assign n40570 = n40569 ^ n40562;
  assign n40571 = n40568 & ~n40570;
  assign n40572 = n40571 ^ n40567;
  assign n40573 = n40572 ^ n40489;
  assign n40574 = ~n40559 & n40573;
  assign n40575 = n40574 ^ n40558;
  assign n40577 = n40576 ^ n40575;
  assign n40578 = n38268 ^ n29671;
  assign n40579 = n40578 ^ n34763;
  assign n40580 = n40579 ^ n28534;
  assign n40581 = n40580 ^ n40576;
  assign n40582 = n40577 & ~n40581;
  assign n40583 = n40582 ^ n40580;
  assign n40584 = n40583 ^ n40554;
  assign n40585 = ~n40555 & n40584;
  assign n40586 = n40585 ^ n40553;
  assign n40587 = n40586 ^ n40549;
  assign n40588 = ~n40550 & n40587;
  assign n40589 = n40588 ^ n40548;
  assign n40542 = n38259 ^ n29662;
  assign n40543 = n40542 ^ n1592;
  assign n40544 = n40543 ^ n28510;
  assign n40434 = n40433 ^ n40408;
  assign n40435 = ~n40409 & ~n40434;
  assign n40436 = n40435 ^ n37444;
  assign n40352 = n40351 ^ n40082;
  assign n40353 = n40087 & n40352;
  assign n40354 = n40353 ^ n40086;
  assign n40077 = n38425 ^ n38206;
  assign n40078 = n39392 ^ n38425;
  assign n40079 = n40077 & n40078;
  assign n40080 = n40079 ^ n38206;
  assign n40405 = n40354 ^ n40080;
  assign n40076 = n39922 ^ n39921;
  assign n40406 = n40405 ^ n40076;
  assign n40407 = n40406 ^ n37437;
  assign n40494 = n40436 ^ n40407;
  assign n40493 = n40487 & ~n40492;
  assign n40541 = n40494 ^ n40493;
  assign n40545 = n40544 ^ n40541;
  assign n40732 = n40589 ^ n40545;
  assign n41680 = n40732 ^ n40038;
  assign n41681 = ~n41679 & n41680;
  assign n41682 = n41681 ^ n39380;
  assign n40787 = n39534 ^ n38676;
  assign n40788 = n40096 ^ n39534;
  assign n40789 = n40787 & ~n40788;
  assign n40790 = n40789 ^ n38676;
  assign n40682 = n39988 ^ n39985;
  assign n40791 = n40790 ^ n40682;
  assign n40792 = n39342 ^ n38592;
  assign n40793 = n40102 ^ n39342;
  assign n40794 = ~n40792 & ~n40793;
  assign n40795 = n40794 ^ n38592;
  assign n40689 = n39980 ^ n39854;
  assign n40796 = n40795 ^ n40689;
  assign n40797 = n39495 ^ n38486;
  assign n40798 = n40108 ^ n39495;
  assign n40799 = n40797 & n40798;
  assign n40800 = n40799 ^ n38486;
  assign n40695 = n39977 ^ n39859;
  assign n40801 = n40800 ^ n40695;
  assign n40802 = n39467 ^ n38492;
  assign n40803 = n40114 ^ n39467;
  assign n40804 = n40802 & n40803;
  assign n40805 = n40804 ^ n38492;
  assign n40702 = n39974 ^ n39864;
  assign n40806 = n40805 ^ n40702;
  assign n40807 = n39445 ^ n38498;
  assign n40808 = n40120 ^ n39445;
  assign n40809 = ~n40807 & n40808;
  assign n40810 = n40809 ^ n38498;
  assign n40710 = n39971 ^ n39869;
  assign n40811 = n40810 ^ n40710;
  assign n40812 = n39447 ^ n38378;
  assign n40813 = n40122 ^ n39447;
  assign n40814 = n40812 & ~n40813;
  assign n40815 = n40814 ^ n38378;
  assign n40716 = n39968 ^ n39874;
  assign n40816 = n40815 ^ n40716;
  assign n40646 = n39965 ^ n39962;
  assign n40642 = n39331 ^ n38385;
  assign n40643 = n40018 ^ n39331;
  assign n40644 = ~n40642 & ~n40643;
  assign n40645 = n40644 ^ n38385;
  assign n40647 = n40646 ^ n40645;
  assign n40476 = n39957 ^ n39876;
  assign n40472 = n39126 ^ n38392;
  assign n40473 = n39798 ^ n39126;
  assign n40474 = n40472 & ~n40473;
  assign n40475 = n40474 ^ n38392;
  assign n40477 = n40476 ^ n40475;
  assign n40386 = n39954 ^ n39881;
  assign n40382 = n39068 ^ n38399;
  assign n40383 = n39683 ^ n39068;
  assign n40384 = ~n40382 & ~n40383;
  assign n40385 = n40384 ^ n38399;
  assign n40387 = n40386 ^ n40385;
  assign n40032 = n39951 ^ n39883;
  assign n40028 = n38947 ^ n38406;
  assign n40029 = n39348 ^ n38947;
  assign n40030 = ~n40028 & n40029;
  assign n40031 = n40030 ^ n38406;
  assign n40033 = n40032 ^ n40031;
  assign n40034 = n38413 ^ n38376;
  assign n40035 = n39354 ^ n38376;
  assign n40036 = ~n40034 & ~n40035;
  assign n40037 = n40036 ^ n38413;
  assign n40039 = n40038 ^ n40037;
  assign n40041 = n38420 ^ n38383;
  assign n40042 = n39360 ^ n38383;
  assign n40043 = ~n40041 & n40042;
  assign n40044 = n40043 ^ n38420;
  assign n40040 = n39945 ^ n39893;
  assign n40045 = n40044 ^ n40040;
  assign n40050 = n39942 ^ n39898;
  assign n40046 = n38427 ^ n38390;
  assign n40047 = n39362 ^ n38390;
  assign n40048 = n40046 & n40047;
  assign n40049 = n40048 ^ n38427;
  assign n40051 = n40050 ^ n40049;
  assign n40056 = n39939 ^ n39903;
  assign n40052 = n38434 ^ n38397;
  assign n40053 = n39372 ^ n38397;
  assign n40054 = n40052 & ~n40053;
  assign n40055 = n40054 ^ n38434;
  assign n40057 = n40056 ^ n40055;
  assign n40059 = n38440 ^ n38404;
  assign n40060 = n39374 ^ n38404;
  assign n40061 = n40059 & ~n40060;
  assign n40062 = n40061 ^ n38440;
  assign n40058 = n39936 ^ n39908;
  assign n40063 = n40062 ^ n40058;
  assign n40065 = n38411 ^ n38361;
  assign n40066 = n39380 ^ n38411;
  assign n40067 = ~n40065 & n40066;
  assign n40068 = n40067 ^ n38361;
  assign n40064 = n39933 ^ n39930;
  assign n40069 = n40068 ^ n40064;
  assign n40071 = n38418 ^ n38341;
  assign n40072 = n39386 ^ n38418;
  assign n40073 = ~n40071 & n40072;
  assign n40074 = n40073 ^ n38341;
  assign n40070 = n39925 ^ n39912;
  assign n40075 = n40074 ^ n40070;
  assign n40081 = n40080 ^ n40076;
  assign n40355 = n40354 ^ n40076;
  assign n40356 = ~n40081 & n40355;
  assign n40357 = n40356 ^ n40080;
  assign n40358 = n40357 ^ n40070;
  assign n40359 = n40075 & ~n40358;
  assign n40360 = n40359 ^ n40074;
  assign n40361 = n40360 ^ n40064;
  assign n40362 = n40069 & n40361;
  assign n40363 = n40362 ^ n40068;
  assign n40364 = n40363 ^ n40058;
  assign n40365 = n40063 & ~n40364;
  assign n40366 = n40365 ^ n40062;
  assign n40367 = n40366 ^ n40056;
  assign n40368 = ~n40057 & ~n40367;
  assign n40369 = n40368 ^ n40055;
  assign n40370 = n40369 ^ n40050;
  assign n40371 = n40051 & n40370;
  assign n40372 = n40371 ^ n40049;
  assign n40373 = n40372 ^ n40040;
  assign n40374 = n40045 & ~n40373;
  assign n40375 = n40374 ^ n40044;
  assign n40376 = n40375 ^ n40038;
  assign n40377 = n40039 & n40376;
  assign n40378 = n40377 ^ n40037;
  assign n40379 = n40378 ^ n40032;
  assign n40380 = ~n40033 & ~n40379;
  assign n40381 = n40380 ^ n40031;
  assign n40469 = n40386 ^ n40381;
  assign n40470 = ~n40387 & ~n40469;
  assign n40471 = n40470 ^ n40385;
  assign n40639 = n40476 ^ n40471;
  assign n40640 = n40477 & ~n40639;
  assign n40641 = n40640 ^ n40475;
  assign n40817 = n40646 ^ n40641;
  assign n40818 = n40647 & ~n40817;
  assign n40819 = n40818 ^ n40645;
  assign n40820 = n40819 ^ n40716;
  assign n40821 = n40816 & n40820;
  assign n40822 = n40821 ^ n40815;
  assign n40823 = n40822 ^ n40710;
  assign n40824 = n40811 & ~n40823;
  assign n40825 = n40824 ^ n40810;
  assign n40826 = n40825 ^ n40702;
  assign n40827 = ~n40806 & n40826;
  assign n40828 = n40827 ^ n40805;
  assign n40829 = n40828 ^ n40695;
  assign n40830 = n40801 & ~n40829;
  assign n40831 = n40830 ^ n40800;
  assign n40832 = n40831 ^ n40689;
  assign n40833 = ~n40796 & n40832;
  assign n40834 = n40833 ^ n40795;
  assign n40835 = n40834 ^ n40682;
  assign n40836 = n40791 & ~n40835;
  assign n40837 = n40836 ^ n40790;
  assign n40782 = n39587 ^ n38833;
  assign n40783 = n39587 ^ n39341;
  assign n40784 = n40782 & ~n40783;
  assign n40785 = n40784 ^ n38833;
  assign n40858 = n40837 ^ n40785;
  assign n40675 = n39991 ^ n39849;
  assign n40859 = n40858 ^ n40675;
  assign n40860 = n40859 ^ n38062;
  assign n40861 = n40834 ^ n40791;
  assign n40862 = n40861 ^ n37804;
  assign n40863 = n40831 ^ n40796;
  assign n40864 = n40863 ^ n37472;
  assign n40865 = n40828 ^ n40801;
  assign n40866 = n40865 ^ n37473;
  assign n40867 = n40825 ^ n40806;
  assign n40868 = n40867 ^ n37479;
  assign n40869 = n40822 ^ n40811;
  assign n40870 = n40869 ^ n37489;
  assign n40871 = n40819 ^ n40816;
  assign n40872 = n40871 ^ n37491;
  assign n40648 = n40647 ^ n40641;
  assign n40649 = n40648 ^ n37497;
  assign n40478 = n40477 ^ n40471;
  assign n40479 = n40478 ^ n37503;
  assign n40388 = n40387 ^ n40381;
  assign n40389 = n40388 ^ n37509;
  assign n40390 = n40378 ^ n40033;
  assign n40391 = n40390 ^ n37510;
  assign n40392 = n40375 ^ n40039;
  assign n40393 = n40392 ^ n37516;
  assign n40394 = n40369 ^ n40051;
  assign n40395 = n40394 ^ n37532;
  assign n40396 = n40366 ^ n40057;
  assign n40397 = n40396 ^ n37538;
  assign n40398 = n40363 ^ n40063;
  assign n40399 = n40398 ^ n36782;
  assign n40400 = n40360 ^ n40068;
  assign n40401 = n40400 ^ n40064;
  assign n40402 = n40401 ^ n37422;
  assign n40403 = n40357 ^ n40075;
  assign n40404 = n40403 ^ n37430;
  assign n40437 = n40436 ^ n40406;
  assign n40438 = n40407 & n40437;
  assign n40439 = n40438 ^ n37437;
  assign n40440 = n40439 ^ n40403;
  assign n40441 = ~n40404 & n40440;
  assign n40442 = n40441 ^ n37430;
  assign n40443 = n40442 ^ n40401;
  assign n40444 = ~n40402 & n40443;
  assign n40445 = n40444 ^ n37422;
  assign n40446 = n40445 ^ n40398;
  assign n40447 = n40399 & ~n40446;
  assign n40448 = n40447 ^ n36782;
  assign n40449 = n40448 ^ n40396;
  assign n40450 = n40397 & n40449;
  assign n40451 = n40450 ^ n37538;
  assign n40452 = n40451 ^ n40394;
  assign n40453 = n40395 & ~n40452;
  assign n40454 = n40453 ^ n37532;
  assign n40455 = n40454 ^ n37526;
  assign n40456 = n40372 ^ n40045;
  assign n40457 = n40456 ^ n40454;
  assign n40458 = n40455 & n40457;
  assign n40459 = n40458 ^ n37526;
  assign n40460 = n40459 ^ n40392;
  assign n40461 = ~n40393 & n40460;
  assign n40462 = n40461 ^ n37516;
  assign n40463 = n40462 ^ n40390;
  assign n40464 = n40391 & n40463;
  assign n40465 = n40464 ^ n37510;
  assign n40466 = n40465 ^ n40388;
  assign n40467 = n40389 & n40466;
  assign n40468 = n40467 ^ n37509;
  assign n40636 = n40478 ^ n40468;
  assign n40637 = n40479 & ~n40636;
  assign n40638 = n40637 ^ n37503;
  assign n40873 = n40648 ^ n40638;
  assign n40874 = n40649 & ~n40873;
  assign n40875 = n40874 ^ n37497;
  assign n40876 = n40875 ^ n40871;
  assign n40877 = ~n40872 & ~n40876;
  assign n40878 = n40877 ^ n37491;
  assign n40879 = n40878 ^ n40869;
  assign n40880 = n40870 & ~n40879;
  assign n40881 = n40880 ^ n37489;
  assign n40882 = n40881 ^ n40867;
  assign n40883 = n40868 & n40882;
  assign n40884 = n40883 ^ n37479;
  assign n40885 = n40884 ^ n40865;
  assign n40886 = ~n40866 & n40885;
  assign n40887 = n40886 ^ n37473;
  assign n40888 = n40887 ^ n40863;
  assign n40889 = n40864 & ~n40888;
  assign n40890 = n40889 ^ n37472;
  assign n40891 = n40890 ^ n40861;
  assign n40892 = ~n40862 & n40891;
  assign n40893 = n40892 ^ n37804;
  assign n40894 = n40893 ^ n40859;
  assign n40895 = ~n40860 & n40894;
  assign n40896 = n40895 ^ n38062;
  assign n40786 = n40785 ^ n40675;
  assign n40838 = n40837 ^ n40675;
  assign n40839 = n40786 & ~n40838;
  assign n40840 = n40839 ^ n40785;
  assign n40777 = n38870 ^ n38086;
  assign n40778 = n40208 ^ n38870;
  assign n40779 = ~n40777 & n40778;
  assign n40780 = n40779 ^ n38086;
  assign n40668 = n39999 ^ n39996;
  assign n40781 = n40780 ^ n40668;
  assign n40856 = n40840 ^ n40781;
  assign n40857 = n40856 ^ n37266;
  assign n40920 = n40896 ^ n40857;
  assign n40921 = n40881 ^ n40868;
  assign n40480 = n40479 ^ n40468;
  assign n40481 = n40465 ^ n40389;
  assign n40482 = n40451 ^ n40395;
  assign n40483 = n40448 ^ n40397;
  assign n40484 = n40445 ^ n40399;
  assign n40485 = n40442 ^ n40402;
  assign n40486 = n40439 ^ n40404;
  assign n40495 = ~n40493 & ~n40494;
  assign n40496 = ~n40486 & n40495;
  assign n40497 = n40485 & ~n40496;
  assign n40498 = ~n40484 & n40497;
  assign n40499 = n40483 & ~n40498;
  assign n40500 = ~n40482 & n40499;
  assign n40501 = n40456 ^ n37526;
  assign n40502 = n40501 ^ n40454;
  assign n40503 = n40500 & n40502;
  assign n40504 = n40459 ^ n40393;
  assign n40505 = n40503 & n40504;
  assign n40506 = n40462 ^ n40391;
  assign n40507 = ~n40505 & n40506;
  assign n40508 = n40481 & ~n40507;
  assign n40635 = ~n40480 & n40508;
  assign n40650 = n40649 ^ n40638;
  assign n40922 = n40635 & ~n40650;
  assign n40923 = n40875 ^ n40872;
  assign n40924 = ~n40922 & ~n40923;
  assign n40925 = n40878 ^ n40870;
  assign n40926 = ~n40924 & n40925;
  assign n40927 = n40921 & n40926;
  assign n40928 = n40884 ^ n40866;
  assign n40929 = ~n40927 & ~n40928;
  assign n40930 = n40887 ^ n40864;
  assign n40931 = n40929 & n40930;
  assign n40932 = n40890 ^ n40862;
  assign n40933 = n40931 & ~n40932;
  assign n40934 = n40893 ^ n40860;
  assign n40935 = ~n40933 & n40934;
  assign n40936 = ~n40920 & n40935;
  assign n40897 = n40896 ^ n40856;
  assign n40898 = n40857 & n40897;
  assign n40899 = n40898 ^ n37266;
  assign n40841 = n40840 ^ n40668;
  assign n40842 = n40781 & n40841;
  assign n40843 = n40842 ^ n40780;
  assign n40772 = n38864 ^ n38093;
  assign n40773 = n40303 ^ n38864;
  assign n40774 = ~n40772 & ~n40773;
  assign n40775 = n40774 ^ n38093;
  assign n40661 = n40002 ^ n39844;
  assign n40776 = n40775 ^ n40661;
  assign n40854 = n40843 ^ n40776;
  assign n40855 = n40854 ^ n37273;
  assign n40919 = n40899 ^ n40855;
  assign n40988 = n40936 ^ n40919;
  assign n1131 = n1130 ^ n1064;
  assign n1147 = n1146 ^ n1131;
  assign n1154 = n1153 ^ n1147;
  assign n40989 = n40988 ^ n1154;
  assign n41046 = n40935 ^ n40920;
  assign n40990 = n40934 ^ n40933;
  assign n979 = n969 ^ n933;
  assign n1004 = n1003 ^ n979;
  assign n1011 = n1010 ^ n1004;
  assign n40991 = n40990 ^ n1011;
  assign n40993 = n38738 ^ n868;
  assign n40994 = n40993 ^ n34678;
  assign n40995 = n40994 ^ n995;
  assign n40992 = n40932 ^ n40931;
  assign n40996 = n40995 ^ n40992;
  assign n40998 = n38743 ^ n853;
  assign n40999 = n40998 ^ n34683;
  assign n41000 = n40999 ^ n28455;
  assign n40997 = n40930 ^ n40929;
  assign n41001 = n41000 ^ n40997;
  assign n41002 = n40928 ^ n40927;
  assign n41006 = n41005 ^ n41002;
  assign n41026 = n40926 ^ n40921;
  assign n41010 = n40925 ^ n40924;
  assign n41007 = n38778 ^ n30124;
  assign n41008 = n41007 ^ n34697;
  assign n41009 = n41008 ^ n28470;
  assign n41011 = n41010 ^ n41009;
  assign n41013 = n38758 ^ n29768;
  assign n41014 = n41013 ^ n34703;
  assign n41015 = n41014 ^ n644;
  assign n41012 = n40923 ^ n40922;
  assign n41016 = n41015 ^ n41012;
  assign n40652 = n38767 ^ n29762;
  assign n40653 = n40652 ^ n34824;
  assign n40654 = n40653 ^ n28477;
  assign n40651 = n40650 ^ n40635;
  assign n40655 = n40654 ^ n40651;
  assign n40509 = n40508 ^ n40480;
  assign n40513 = n40512 ^ n40509;
  assign n40514 = n40507 ^ n40481;
  assign n40518 = n40517 ^ n40514;
  assign n40621 = n40506 ^ n40505;
  assign n40520 = n29646 ^ n2208;
  assign n40521 = n40520 ^ n34722;
  assign n40522 = n40521 ^ n28497;
  assign n40519 = n40504 ^ n40503;
  assign n40523 = n40522 ^ n40519;
  assign n40613 = n40502 ^ n40500;
  assign n40524 = n40499 ^ n40482;
  assign n2114 = n2095 ^ n2047;
  assign n2133 = n2132 ^ n2114;
  assign n2140 = n2139 ^ n2133;
  assign n40525 = n40524 ^ n2140;
  assign n40527 = n38244 ^ n1964;
  assign n40528 = n40527 ^ n34732;
  assign n40529 = n40528 ^ n2124;
  assign n40526 = n40498 ^ n40483;
  assign n40530 = n40529 ^ n40526;
  assign n40532 = n38310 ^ n1949;
  assign n40533 = n40532 ^ n34737;
  assign n40534 = n40533 ^ n28504;
  assign n40531 = n40497 ^ n40484;
  assign n40535 = n40534 ^ n40531;
  assign n40596 = n40496 ^ n40485;
  assign n40539 = n40495 ^ n40486;
  assign n40536 = n38254 ^ n29704;
  assign n40537 = n40536 ^ n34746;
  assign n40538 = n40537 ^ n1658;
  assign n40540 = n40539 ^ n40538;
  assign n40590 = n40589 ^ n40541;
  assign n40591 = ~n40545 & n40590;
  assign n40592 = n40591 ^ n40544;
  assign n40593 = n40592 ^ n40539;
  assign n40594 = n40540 & ~n40593;
  assign n40595 = n40594 ^ n40538;
  assign n40597 = n40596 ^ n40595;
  assign n40598 = n38249 ^ n29656;
  assign n40599 = n40598 ^ n34742;
  assign n40600 = n40599 ^ n28556;
  assign n40601 = n40600 ^ n40596;
  assign n40602 = n40597 & ~n40601;
  assign n40603 = n40602 ^ n40600;
  assign n40604 = n40603 ^ n40531;
  assign n40605 = ~n40535 & n40604;
  assign n40606 = n40605 ^ n40534;
  assign n40607 = n40606 ^ n40526;
  assign n40608 = n40530 & ~n40607;
  assign n40609 = n40608 ^ n40529;
  assign n40610 = n40609 ^ n40524;
  assign n40611 = n40525 & ~n40610;
  assign n40612 = n40611 ^ n2140;
  assign n40614 = n40613 ^ n40612;
  assign n40615 = n40613 ^ n2158;
  assign n40616 = n40614 & ~n40615;
  assign n40617 = n40616 ^ n2158;
  assign n40618 = n40617 ^ n40519;
  assign n40619 = ~n40523 & n40618;
  assign n40620 = n40619 ^ n40522;
  assign n40622 = n40621 ^ n40620;
  assign n40626 = n40625 ^ n40621;
  assign n40627 = n40622 & ~n40626;
  assign n40628 = n40627 ^ n40625;
  assign n40629 = n40628 ^ n40514;
  assign n40630 = n40518 & ~n40629;
  assign n40631 = n40630 ^ n40517;
  assign n40632 = n40631 ^ n40509;
  assign n40633 = n40513 & ~n40632;
  assign n40634 = n40633 ^ n40512;
  assign n41017 = n40651 ^ n40634;
  assign n41018 = n40655 & ~n41017;
  assign n41019 = n41018 ^ n40654;
  assign n41020 = n41019 ^ n41012;
  assign n41021 = n41016 & ~n41020;
  assign n41022 = n41021 ^ n41015;
  assign n41023 = n41022 ^ n41010;
  assign n41024 = n41011 & ~n41023;
  assign n41025 = n41024 ^ n41009;
  assign n41027 = n41026 ^ n41025;
  assign n41028 = n38752 ^ n30137;
  assign n41029 = n41028 ^ n34692;
  assign n41030 = n41029 ^ n28464;
  assign n41031 = n41030 ^ n41026;
  assign n41032 = n41027 & ~n41031;
  assign n41033 = n41032 ^ n41030;
  assign n41034 = n41033 ^ n41002;
  assign n41035 = n41006 & ~n41034;
  assign n41036 = n41035 ^ n41005;
  assign n41037 = n41036 ^ n40997;
  assign n41038 = n41001 & ~n41037;
  assign n41039 = n41038 ^ n41000;
  assign n41040 = n41039 ^ n40992;
  assign n41041 = ~n40996 & n41040;
  assign n41042 = n41041 ^ n40995;
  assign n41043 = n41042 ^ n40990;
  assign n41044 = n40991 & ~n41043;
  assign n41045 = n41044 ^ n1011;
  assign n41047 = n41046 ^ n41045;
  assign n41048 = n38731 ^ n30108;
  assign n41049 = n41048 ^ n1021;
  assign n41050 = n41049 ^ n1138;
  assign n41051 = n41050 ^ n41046;
  assign n41052 = ~n41047 & n41051;
  assign n41053 = n41052 ^ n41050;
  assign n41054 = n41053 ^ n40988;
  assign n41055 = n40989 & ~n41054;
  assign n41056 = n41055 ^ n1154;
  assign n40937 = ~n40919 & n40936;
  assign n40900 = n40899 ^ n40854;
  assign n40901 = ~n40855 & ~n40900;
  assign n40902 = n40901 ^ n37273;
  assign n40847 = n38858 ^ n38080;
  assign n40848 = n39618 ^ n38858;
  assign n40849 = n40847 & ~n40848;
  assign n40850 = n40849 ^ n38080;
  assign n40024 = n40023 ^ n40005;
  assign n40851 = n40850 ^ n40024;
  assign n40844 = n40843 ^ n40661;
  assign n40845 = ~n40776 & n40844;
  assign n40846 = n40845 ^ n40775;
  assign n40852 = n40851 ^ n40846;
  assign n40853 = n40852 ^ n37260;
  assign n40918 = n40902 ^ n40853;
  assign n40986 = n40937 ^ n40918;
  assign n40983 = n38725 ^ n30163;
  assign n40984 = n40983 ^ n34667;
  assign n40985 = n40984 ^ n1329;
  assign n40987 = n40986 ^ n40985;
  assign n41112 = n41056 ^ n40987;
  assign n41113 = n39420 ^ n38458;
  assign n41114 = n40082 ^ n39420;
  assign n41115 = ~n41113 & n41114;
  assign n41116 = n41115 ^ n38458;
  assign n41117 = ~n41112 & n41116;
  assign n41106 = n39410 ^ n38456;
  assign n41107 = n40076 ^ n39410;
  assign n41108 = n41106 & n41107;
  assign n41109 = n41108 ^ n38456;
  assign n41248 = n41117 ^ n41109;
  assign n41062 = n38721 ^ n30101;
  assign n41063 = n41062 ^ n1337;
  assign n41064 = n41063 ^ n28625;
  assign n40938 = n40918 & n40937;
  assign n40914 = n40260 ^ n40257;
  assign n40909 = n38852 ^ n38070;
  assign n40910 = n39621 ^ n38852;
  assign n40911 = n40909 & n40910;
  assign n40912 = n40911 ^ n38070;
  assign n40906 = n40846 ^ n40024;
  assign n40907 = ~n40851 & ~n40906;
  assign n40908 = n40907 ^ n40850;
  assign n40913 = n40912 ^ n40908;
  assign n40915 = n40914 ^ n40913;
  assign n40916 = n40915 ^ n37254;
  assign n40903 = n40902 ^ n40852;
  assign n40904 = ~n40853 & n40903;
  assign n40905 = n40904 ^ n37260;
  assign n40917 = n40916 ^ n40905;
  assign n41060 = n40938 ^ n40917;
  assign n41057 = n41056 ^ n40986;
  assign n41058 = ~n40987 & n41057;
  assign n41059 = n41058 ^ n40985;
  assign n41061 = n41060 ^ n41059;
  assign n41110 = n41064 ^ n41061;
  assign n41249 = n41248 ^ n41110;
  assign n41245 = n41116 ^ n41112;
  assign n41246 = ~n37442 & ~n41245;
  assign n41247 = n41246 ^ n37435;
  assign n41474 = n41249 ^ n41247;
  assign n41470 = n39221 ^ n30621;
  assign n41471 = n41470 ^ n35072;
  assign n41472 = n41471 ^ n28811;
  assign n41465 = n41245 ^ n37442;
  assign n41466 = n39440 ^ n30976;
  assign n41467 = n41466 ^ n2501;
  assign n41468 = n41467 ^ n29449;
  assign n41469 = n41465 & n41468;
  assign n41473 = n41472 ^ n41469;
  assign n41678 = n41474 ^ n41473;
  assign n41683 = n41682 ^ n41678;
  assign n41685 = n40040 ^ n39386;
  assign n40738 = n40586 ^ n40550;
  assign n41686 = n40738 ^ n40040;
  assign n41687 = ~n41685 & ~n41686;
  assign n41688 = n41687 ^ n39386;
  assign n41684 = n41468 ^ n41465;
  assign n41689 = n41688 ^ n41684;
  assign n41728 = n41042 ^ n40991;
  assign n41699 = n39598 ^ n38852;
  assign n41700 = n40332 ^ n39598;
  assign n41701 = ~n41699 & n41700;
  assign n41702 = n41701 ^ n38852;
  assign n41698 = n41039 ^ n40996;
  assign n41703 = n41702 ^ n41698;
  assign n41705 = n39608 ^ n38858;
  assign n41706 = n40338 ^ n39608;
  assign n41707 = n41705 & ~n41706;
  assign n41708 = n41707 ^ n38858;
  assign n41704 = n41036 ^ n41001;
  assign n41709 = n41708 ^ n41704;
  assign n41711 = n39621 ^ n38864;
  assign n41087 = n40274 ^ n40247;
  assign n41712 = n41087 ^ n39621;
  assign n41713 = n41711 & ~n41712;
  assign n41714 = n41713 ^ n38864;
  assign n41710 = n41033 ^ n41006;
  assign n41715 = n41714 ^ n41710;
  assign n41583 = n39618 ^ n38870;
  assign n40968 = n40271 ^ n40268;
  assign n41584 = n40968 ^ n39618;
  assign n41585 = n41583 & ~n41584;
  assign n41586 = n41585 ^ n38870;
  assign n41582 = n41030 ^ n41027;
  assign n41587 = n41586 ^ n41582;
  assign n41332 = n41022 ^ n41011;
  assign n41327 = n40303 ^ n39587;
  assign n40952 = n40263 ^ n40252;
  assign n41328 = n40952 ^ n40303;
  assign n41329 = n41327 & ~n41328;
  assign n41330 = n41329 ^ n39587;
  assign n41578 = n41332 ^ n41330;
  assign n41190 = n40208 ^ n39534;
  assign n41191 = n40914 ^ n40208;
  assign n41192 = ~n41190 & ~n41191;
  assign n41193 = n41192 ^ n39534;
  assign n41189 = n41019 ^ n41016;
  assign n41194 = n41193 ^ n41189;
  assign n40656 = n40655 ^ n40634;
  assign n39343 = n39342 ^ n39341;
  assign n40025 = n40024 ^ n39341;
  assign n40026 = ~n39343 & n40025;
  assign n40027 = n40026 ^ n39342;
  assign n40657 = n40656 ^ n40027;
  assign n40660 = n40096 ^ n39495;
  assign n40662 = n40661 ^ n40096;
  assign n40663 = n40660 & ~n40662;
  assign n40664 = n40663 ^ n39495;
  assign n40658 = n40631 ^ n40512;
  assign n40659 = n40658 ^ n40509;
  assign n40665 = n40664 ^ n40659;
  assign n40667 = n40102 ^ n39467;
  assign n40669 = n40668 ^ n40102;
  assign n40670 = ~n40667 & ~n40669;
  assign n40671 = n40670 ^ n39467;
  assign n40666 = n40628 ^ n40518;
  assign n40672 = n40671 ^ n40666;
  assign n40674 = n40108 ^ n39445;
  assign n40676 = n40675 ^ n40108;
  assign n40677 = n40674 & n40676;
  assign n40678 = n40677 ^ n39445;
  assign n40673 = n40625 ^ n40622;
  assign n40679 = n40678 ^ n40673;
  assign n40681 = n40114 ^ n39447;
  assign n40683 = n40682 ^ n40114;
  assign n40684 = ~n40681 & n40683;
  assign n40685 = n40684 ^ n39447;
  assign n40680 = n40617 ^ n40523;
  assign n40686 = n40685 ^ n40680;
  assign n40688 = n40120 ^ n39331;
  assign n40690 = n40689 ^ n40120;
  assign n40691 = n40688 & n40690;
  assign n40692 = n40691 ^ n39331;
  assign n40687 = n40614 ^ n2158;
  assign n40693 = n40692 ^ n40687;
  assign n40699 = n40609 ^ n40525;
  assign n40694 = n40122 ^ n39126;
  assign n40696 = n40695 ^ n40122;
  assign n40697 = ~n40694 & ~n40696;
  assign n40698 = n40697 ^ n39126;
  assign n40700 = n40699 ^ n40698;
  assign n40706 = n40606 ^ n40530;
  assign n40701 = n40018 ^ n39068;
  assign n40703 = n40702 ^ n40018;
  assign n40704 = n40701 & n40703;
  assign n40705 = n40704 ^ n39068;
  assign n40707 = n40706 ^ n40705;
  assign n40709 = n39798 ^ n38947;
  assign n40711 = n40710 ^ n39798;
  assign n40712 = n40709 & n40711;
  assign n40713 = n40712 ^ n38947;
  assign n40708 = n40603 ^ n40535;
  assign n40714 = n40713 ^ n40708;
  assign n40720 = n40600 ^ n40597;
  assign n40715 = n39683 ^ n38376;
  assign n40717 = n40716 ^ n39683;
  assign n40718 = n40715 & ~n40717;
  assign n40719 = n40718 ^ n38376;
  assign n40721 = n40720 ^ n40719;
  assign n40726 = n40592 ^ n40540;
  assign n40722 = n39348 ^ n38383;
  assign n40723 = n40646 ^ n39348;
  assign n40724 = ~n40722 & n40723;
  assign n40725 = n40724 ^ n38383;
  assign n40727 = n40726 ^ n40725;
  assign n40728 = n39354 ^ n38390;
  assign n40729 = n40476 ^ n39354;
  assign n40730 = n40728 & n40729;
  assign n40731 = n40730 ^ n38390;
  assign n40733 = n40732 ^ n40731;
  assign n40734 = n39360 ^ n38397;
  assign n40735 = n40386 ^ n39360;
  assign n40736 = ~n40734 & ~n40735;
  assign n40737 = n40736 ^ n38397;
  assign n40739 = n40738 ^ n40737;
  assign n40741 = n39362 ^ n38404;
  assign n40742 = n40032 ^ n39362;
  assign n40743 = ~n40741 & ~n40742;
  assign n40744 = n40743 ^ n38404;
  assign n40740 = n40583 ^ n40555;
  assign n40745 = n40744 ^ n40740;
  assign n40747 = n39372 ^ n38411;
  assign n40748 = n40038 ^ n39372;
  assign n40749 = n40747 & ~n40748;
  assign n40750 = n40749 ^ n38411;
  assign n40746 = n40580 ^ n40577;
  assign n40751 = n40750 ^ n40746;
  assign n40754 = n39380 ^ n38425;
  assign n40755 = n40050 ^ n39380;
  assign n40756 = ~n40754 & ~n40755;
  assign n40757 = n40756 ^ n38425;
  assign n40753 = n40569 ^ n40568;
  assign n40758 = n40757 ^ n40753;
  assign n40763 = n40566 ^ n40565;
  assign n40759 = n39386 ^ n38432;
  assign n40760 = n40056 ^ n39386;
  assign n40761 = n40759 & n40760;
  assign n40762 = n40761 ^ n38432;
  assign n40764 = n40763 ^ n40762;
  assign n40939 = n40917 & ~n40938;
  assign n40947 = n38846 ^ n38068;
  assign n40948 = n39608 ^ n38846;
  assign n40949 = ~n40947 & ~n40948;
  assign n40950 = n40949 ^ n38068;
  assign n40943 = n40914 ^ n40912;
  assign n40944 = n40914 ^ n40908;
  assign n40945 = n40943 & n40944;
  assign n40946 = n40945 ^ n40912;
  assign n40951 = n40950 ^ n40946;
  assign n40953 = n40952 ^ n40951;
  assign n40954 = n40953 ^ n37312;
  assign n40940 = n40915 ^ n40905;
  assign n40941 = n40916 & n40940;
  assign n40942 = n40941 ^ n37254;
  assign n40955 = n40954 ^ n40942;
  assign n40956 = n40939 & ~n40955;
  assign n40964 = n40952 ^ n40950;
  assign n40965 = n40952 ^ n40946;
  assign n40966 = ~n40964 & n40965;
  assign n40967 = n40966 ^ n40950;
  assign n40969 = n40968 ^ n40967;
  assign n40960 = n38469 ^ n37456;
  assign n40961 = n39598 ^ n38469;
  assign n40962 = ~n40960 & n40961;
  assign n40963 = n40962 ^ n37456;
  assign n40970 = n40969 ^ n40963;
  assign n40971 = n40970 ^ n37345;
  assign n40957 = n40953 ^ n40942;
  assign n40958 = n40954 & ~n40957;
  assign n40959 = n40958 ^ n37312;
  assign n40972 = n40971 ^ n40959;
  assign n41090 = n40956 & ~n40972;
  assign n41082 = n38463 ^ n37449;
  assign n41083 = n39596 ^ n38463;
  assign n41084 = n41082 & n41083;
  assign n41085 = n41084 ^ n37449;
  assign n41079 = n40968 ^ n40963;
  assign n41080 = n40969 & n41079;
  assign n41081 = n41080 ^ n40963;
  assign n41086 = n41085 ^ n41081;
  assign n41088 = n41087 ^ n41086;
  assign n41075 = n40970 ^ n40959;
  assign n41076 = n40971 & n41075;
  assign n41077 = n41076 ^ n37345;
  assign n41078 = n41077 ^ n37414;
  assign n41089 = n41088 ^ n41078;
  assign n41091 = n41090 ^ n41089;
  assign n40974 = n38716 ^ n30091;
  assign n40975 = n40974 ^ n34939;
  assign n40976 = n40975 ^ n28438;
  assign n40973 = n40972 ^ n40956;
  assign n40977 = n40976 ^ n40973;
  assign n40979 = n38815 ^ n30096;
  assign n40980 = n40979 ^ n34913;
  assign n40981 = n40980 ^ n2324;
  assign n40978 = n40955 ^ n40939;
  assign n40982 = n40981 ^ n40978;
  assign n41065 = n41064 ^ n41060;
  assign n41066 = n41061 & ~n41065;
  assign n41067 = n41066 ^ n41064;
  assign n41068 = n41067 ^ n40978;
  assign n41069 = ~n40982 & n41068;
  assign n41070 = n41069 ^ n40981;
  assign n41071 = n41070 ^ n40973;
  assign n41072 = ~n40977 & n41071;
  assign n41073 = n41072 ^ n40976;
  assign n40769 = n38477 ^ n2600;
  assign n40770 = n40769 ^ n35004;
  assign n40771 = n40770 ^ n28433;
  assign n41074 = n41073 ^ n40771;
  assign n41092 = n41091 ^ n41074;
  assign n40765 = n39392 ^ n38444;
  assign n40766 = n40058 ^ n39392;
  assign n40767 = n40765 & ~n40766;
  assign n40768 = n40767 ^ n38444;
  assign n41093 = n41092 ^ n40768;
  assign n41095 = n39398 ^ n38904;
  assign n41096 = n40064 ^ n39398;
  assign n41097 = ~n41095 & n41096;
  assign n41098 = n41097 ^ n38904;
  assign n41094 = n41070 ^ n40977;
  assign n41099 = n41098 ^ n41094;
  assign n41104 = n41067 ^ n40982;
  assign n41100 = n39404 ^ n38450;
  assign n41101 = n40070 ^ n39404;
  assign n41102 = ~n41100 & ~n41101;
  assign n41103 = n41102 ^ n38450;
  assign n41105 = n41104 ^ n41103;
  assign n41111 = n41110 ^ n41109;
  assign n41118 = n41117 ^ n41110;
  assign n41119 = n41111 & ~n41118;
  assign n41120 = n41119 ^ n41117;
  assign n41121 = n41120 ^ n41104;
  assign n41122 = n41105 & n41121;
  assign n41123 = n41122 ^ n41103;
  assign n41124 = n41123 ^ n41094;
  assign n41125 = n41099 & ~n41124;
  assign n41126 = n41125 ^ n41098;
  assign n41127 = n41126 ^ n41092;
  assign n41128 = n41093 & ~n41127;
  assign n41129 = n41128 ^ n40768;
  assign n41130 = n41129 ^ n40763;
  assign n41131 = n40764 & n41130;
  assign n41132 = n41131 ^ n40762;
  assign n41133 = n41132 ^ n40753;
  assign n41134 = n40758 & ~n41133;
  assign n41135 = n41134 ^ n40757;
  assign n40752 = n40572 ^ n40559;
  assign n41136 = n41135 ^ n40752;
  assign n41137 = n39374 ^ n38418;
  assign n41138 = n40040 ^ n39374;
  assign n41139 = n41137 & ~n41138;
  assign n41140 = n41139 ^ n38418;
  assign n41141 = n41140 ^ n41135;
  assign n41142 = ~n41136 & n41141;
  assign n41143 = n41142 ^ n40752;
  assign n41144 = n41143 ^ n40746;
  assign n41145 = ~n40751 & ~n41144;
  assign n41146 = n41145 ^ n40750;
  assign n41147 = n41146 ^ n40740;
  assign n41148 = n40745 & n41147;
  assign n41149 = n41148 ^ n40744;
  assign n41150 = n41149 ^ n40738;
  assign n41151 = ~n40739 & ~n41150;
  assign n41152 = n41151 ^ n40737;
  assign n41153 = n41152 ^ n40732;
  assign n41154 = n40733 & n41153;
  assign n41155 = n41154 ^ n40731;
  assign n41156 = n41155 ^ n40726;
  assign n41157 = n40727 & n41156;
  assign n41158 = n41157 ^ n40725;
  assign n41159 = n41158 ^ n40720;
  assign n41160 = n40721 & n41159;
  assign n41161 = n41160 ^ n40719;
  assign n41162 = n41161 ^ n40708;
  assign n41163 = ~n40714 & ~n41162;
  assign n41164 = n41163 ^ n40713;
  assign n41165 = n41164 ^ n40706;
  assign n41166 = ~n40707 & ~n41165;
  assign n41167 = n41166 ^ n40705;
  assign n41168 = n41167 ^ n40699;
  assign n41169 = n40700 & n41168;
  assign n41170 = n41169 ^ n40698;
  assign n41171 = n41170 ^ n40687;
  assign n41172 = n40693 & n41171;
  assign n41173 = n41172 ^ n40692;
  assign n41174 = n41173 ^ n40680;
  assign n41175 = n40686 & ~n41174;
  assign n41176 = n41175 ^ n40685;
  assign n41177 = n41176 ^ n40673;
  assign n41178 = ~n40679 & ~n41177;
  assign n41179 = n41178 ^ n40678;
  assign n41180 = n41179 ^ n40666;
  assign n41181 = ~n40672 & ~n41180;
  assign n41182 = n41181 ^ n40671;
  assign n41183 = n41182 ^ n40659;
  assign n41184 = ~n40665 & n41183;
  assign n41185 = n41184 ^ n40664;
  assign n41186 = n41185 ^ n40656;
  assign n41187 = n40657 & n41186;
  assign n41188 = n41187 ^ n40027;
  assign n41324 = n41189 ^ n41188;
  assign n41325 = ~n41194 & ~n41324;
  assign n41326 = n41325 ^ n41193;
  assign n41579 = n41332 ^ n41326;
  assign n41580 = ~n41578 & n41579;
  assign n41581 = n41580 ^ n41330;
  assign n41716 = n41582 ^ n41581;
  assign n41717 = n41587 & ~n41716;
  assign n41718 = n41717 ^ n41586;
  assign n41719 = n41718 ^ n41710;
  assign n41720 = ~n41715 & n41719;
  assign n41721 = n41720 ^ n41714;
  assign n41722 = n41721 ^ n41704;
  assign n41723 = ~n41709 & n41722;
  assign n41724 = n41723 ^ n41708;
  assign n41725 = n41724 ^ n41698;
  assign n41726 = ~n41703 & ~n41725;
  assign n41727 = n41726 ^ n41702;
  assign n41729 = n41728 ^ n41727;
  assign n41694 = n39596 ^ n38846;
  assign n41695 = n40326 ^ n39596;
  assign n41696 = n41694 & n41695;
  assign n41697 = n41696 ^ n38846;
  assign n41758 = n41728 ^ n41697;
  assign n41759 = ~n41729 & ~n41758;
  assign n41760 = n41759 ^ n41697;
  assign n41597 = n41050 ^ n41047;
  assign n41761 = n41760 ^ n41597;
  assign n41754 = n39428 ^ n38469;
  assign n41755 = n40320 ^ n39428;
  assign n41756 = ~n41754 & ~n41755;
  assign n41757 = n41756 ^ n38469;
  assign n41762 = n41761 ^ n41757;
  assign n41763 = n41762 ^ n37456;
  assign n41730 = n41729 ^ n41697;
  assign n41731 = n41730 ^ n38068;
  assign n41732 = n41724 ^ n41702;
  assign n41733 = n41732 ^ n41698;
  assign n41734 = n41733 ^ n38070;
  assign n41735 = n41721 ^ n41709;
  assign n41736 = n41735 ^ n38080;
  assign n41737 = n41718 ^ n41715;
  assign n41738 = n41737 ^ n38093;
  assign n41588 = n41587 ^ n41581;
  assign n41589 = n41588 ^ n38086;
  assign n41331 = n41330 ^ n41326;
  assign n41333 = n41332 ^ n41331;
  assign n41334 = n41333 ^ n38833;
  assign n41195 = n41194 ^ n41188;
  assign n41196 = n41195 ^ n38676;
  assign n41197 = n41185 ^ n40657;
  assign n41198 = n41197 ^ n38592;
  assign n41199 = n41182 ^ n40665;
  assign n41200 = n41199 ^ n38486;
  assign n41201 = n41179 ^ n40672;
  assign n41202 = n41201 ^ n38492;
  assign n41203 = n41176 ^ n40679;
  assign n41204 = n41203 ^ n38498;
  assign n41205 = n41173 ^ n40686;
  assign n41206 = n41205 ^ n38378;
  assign n41207 = n41170 ^ n40693;
  assign n41208 = n41207 ^ n38385;
  assign n41209 = n41167 ^ n40698;
  assign n41210 = n41209 ^ n40699;
  assign n41211 = n41210 ^ n38392;
  assign n41212 = n41164 ^ n40707;
  assign n41213 = n41212 ^ n38399;
  assign n41214 = n41161 ^ n40713;
  assign n41215 = n41214 ^ n40708;
  assign n41216 = n41215 ^ n38406;
  assign n41217 = n41158 ^ n40719;
  assign n41218 = n41217 ^ n40720;
  assign n41219 = n41218 ^ n38413;
  assign n41220 = n41155 ^ n40727;
  assign n41221 = n41220 ^ n38420;
  assign n41222 = n41152 ^ n40731;
  assign n41223 = n41222 ^ n40732;
  assign n41224 = n41223 ^ n38427;
  assign n41225 = n41149 ^ n40737;
  assign n41226 = n41225 ^ n40738;
  assign n41227 = n41226 ^ n38434;
  assign n41228 = n41146 ^ n40744;
  assign n41229 = n41228 ^ n40740;
  assign n41230 = n41229 ^ n38440;
  assign n41231 = n41143 ^ n40750;
  assign n41232 = n41231 ^ n40746;
  assign n41233 = n41232 ^ n38361;
  assign n41234 = n41132 ^ n40757;
  assign n41235 = n41234 ^ n40753;
  assign n41236 = n41235 ^ n38206;
  assign n41262 = n41129 ^ n40764;
  assign n41237 = n41126 ^ n41093;
  assign n41238 = n41237 ^ n37419;
  assign n41239 = n41123 ^ n41098;
  assign n41240 = n41239 ^ n41094;
  assign n41241 = n41240 ^ n37426;
  assign n41242 = n41120 ^ n41103;
  assign n41243 = n41242 ^ n41104;
  assign n41244 = n41243 ^ n37428;
  assign n41250 = n41249 ^ n41246;
  assign n41251 = ~n41247 & n41250;
  assign n41252 = n41251 ^ n37435;
  assign n41253 = n41252 ^ n41243;
  assign n41254 = n41244 & n41253;
  assign n41255 = n41254 ^ n37428;
  assign n41256 = n41255 ^ n41240;
  assign n41257 = n41241 & n41256;
  assign n41258 = n41257 ^ n37426;
  assign n41259 = n41258 ^ n41237;
  assign n41260 = n41238 & ~n41259;
  assign n41261 = n41260 ^ n37419;
  assign n41263 = n41262 ^ n41261;
  assign n41264 = n41262 ^ n38131;
  assign n41265 = ~n41263 & ~n41264;
  assign n41266 = n41265 ^ n38131;
  assign n41267 = n41266 ^ n41235;
  assign n41268 = n41236 & ~n41267;
  assign n41269 = n41268 ^ n38206;
  assign n41270 = n41269 ^ n38341;
  assign n41271 = n41140 ^ n40752;
  assign n41272 = n41271 ^ n41135;
  assign n41273 = n41272 ^ n41269;
  assign n41274 = n41270 & ~n41273;
  assign n41275 = n41274 ^ n38341;
  assign n41276 = n41275 ^ n41232;
  assign n41277 = ~n41233 & ~n41276;
  assign n41278 = n41277 ^ n38361;
  assign n41279 = n41278 ^ n41229;
  assign n41280 = ~n41230 & n41279;
  assign n41281 = n41280 ^ n38440;
  assign n41282 = n41281 ^ n41226;
  assign n41283 = n41227 & n41282;
  assign n41284 = n41283 ^ n38434;
  assign n41285 = n41284 ^ n41223;
  assign n41286 = ~n41224 & ~n41285;
  assign n41287 = n41286 ^ n38427;
  assign n41288 = n41287 ^ n41220;
  assign n41289 = n41221 & ~n41288;
  assign n41290 = n41289 ^ n38420;
  assign n41291 = n41290 ^ n41218;
  assign n41292 = n41219 & n41291;
  assign n41293 = n41292 ^ n38413;
  assign n41294 = n41293 ^ n41215;
  assign n41295 = ~n41216 & ~n41294;
  assign n41296 = n41295 ^ n38406;
  assign n41297 = n41296 ^ n41212;
  assign n41298 = ~n41213 & ~n41297;
  assign n41299 = n41298 ^ n38399;
  assign n41300 = n41299 ^ n41210;
  assign n41301 = ~n41211 & n41300;
  assign n41302 = n41301 ^ n38392;
  assign n41303 = n41302 ^ n41207;
  assign n41304 = n41208 & ~n41303;
  assign n41305 = n41304 ^ n38385;
  assign n41306 = n41305 ^ n41205;
  assign n41307 = n41206 & n41306;
  assign n41308 = n41307 ^ n38378;
  assign n41309 = n41308 ^ n41203;
  assign n41310 = ~n41204 & n41309;
  assign n41311 = n41310 ^ n38498;
  assign n41312 = n41311 ^ n41201;
  assign n41313 = n41202 & ~n41312;
  assign n41314 = n41313 ^ n38492;
  assign n41315 = n41314 ^ n41199;
  assign n41316 = ~n41200 & n41315;
  assign n41317 = n41316 ^ n38486;
  assign n41318 = n41317 ^ n41197;
  assign n41319 = n41198 & ~n41318;
  assign n41320 = n41319 ^ n38592;
  assign n41321 = n41320 ^ n41195;
  assign n41322 = n41196 & ~n41321;
  assign n41323 = n41322 ^ n38676;
  assign n41575 = n41333 ^ n41323;
  assign n41576 = ~n41334 & n41575;
  assign n41577 = n41576 ^ n38833;
  assign n41739 = n41588 ^ n41577;
  assign n41740 = ~n41589 & ~n41739;
  assign n41741 = n41740 ^ n38086;
  assign n41742 = n41741 ^ n41737;
  assign n41743 = n41738 & ~n41742;
  assign n41744 = n41743 ^ n38093;
  assign n41745 = n41744 ^ n41735;
  assign n41746 = ~n41736 & ~n41745;
  assign n41747 = n41746 ^ n38080;
  assign n41748 = n41747 ^ n41733;
  assign n41749 = n41734 & n41748;
  assign n41750 = n41749 ^ n38070;
  assign n41751 = n41750 ^ n41730;
  assign n41752 = ~n41731 & n41751;
  assign n41753 = n41752 ^ n38068;
  assign n41764 = n41763 ^ n41753;
  assign n41765 = n41744 ^ n41736;
  assign n41766 = n41741 ^ n41738;
  assign n41335 = n41334 ^ n41323;
  assign n41336 = n41317 ^ n41198;
  assign n41337 = n41314 ^ n41200;
  assign n41338 = n41299 ^ n41211;
  assign n41339 = n41293 ^ n38406;
  assign n41340 = n41339 ^ n41215;
  assign n41341 = n41281 ^ n41227;
  assign n41342 = n41275 ^ n41233;
  assign n41343 = n41272 ^ n38341;
  assign n41344 = n41343 ^ n41269;
  assign n41345 = n41263 ^ n38131;
  assign n41346 = n41258 ^ n41238;
  assign n41347 = n41252 ^ n41244;
  assign n41348 = n41255 ^ n41241;
  assign n41349 = n41347 & ~n41348;
  assign n41350 = n41346 & n41349;
  assign n41351 = n41345 & ~n41350;
  assign n41352 = n41266 ^ n41236;
  assign n41353 = ~n41351 & ~n41352;
  assign n41354 = ~n41344 & n41353;
  assign n41355 = ~n41342 & ~n41354;
  assign n41356 = n41278 ^ n41230;
  assign n41357 = n41355 & n41356;
  assign n41358 = n41341 & ~n41357;
  assign n41359 = n41284 ^ n41224;
  assign n41360 = n41358 & n41359;
  assign n41361 = n41287 ^ n41221;
  assign n41362 = n41360 & n41361;
  assign n41363 = n41290 ^ n41219;
  assign n41364 = n41362 & n41363;
  assign n41365 = ~n41340 & ~n41364;
  assign n41366 = n41296 ^ n41213;
  assign n41367 = ~n41365 & ~n41366;
  assign n41368 = n41338 & n41367;
  assign n41369 = n41302 ^ n41208;
  assign n41370 = n41368 & ~n41369;
  assign n41371 = n41305 ^ n41206;
  assign n41372 = ~n41370 & n41371;
  assign n41373 = n41308 ^ n41204;
  assign n41374 = ~n41372 & ~n41373;
  assign n41375 = n41311 ^ n41202;
  assign n41376 = n41374 & n41375;
  assign n41377 = n41337 & ~n41376;
  assign n41378 = ~n41336 & n41377;
  assign n41379 = n41320 ^ n41196;
  assign n41380 = n41378 & ~n41379;
  assign n41574 = ~n41335 & ~n41380;
  assign n41590 = n41589 ^ n41577;
  assign n41767 = n41574 & ~n41590;
  assign n41768 = ~n41766 & n41767;
  assign n41769 = n41765 & n41768;
  assign n41770 = n41747 ^ n41734;
  assign n41771 = ~n41769 & ~n41770;
  assign n41772 = n41750 ^ n41731;
  assign n41773 = n41771 & ~n41772;
  assign n41827 = n41764 & n41773;
  assign n41824 = n41053 ^ n40989;
  assign n41819 = n39426 ^ n38463;
  assign n41820 = n40314 ^ n39426;
  assign n41821 = n41819 & n41820;
  assign n41822 = n41821 ^ n38463;
  assign n41816 = n41757 ^ n41597;
  assign n41817 = n41761 & n41816;
  assign n41818 = n41817 ^ n41757;
  assign n41823 = n41822 ^ n41818;
  assign n41825 = n41824 ^ n41823;
  assign n41812 = n41762 ^ n41753;
  assign n41813 = n41763 & n41812;
  assign n41814 = n41813 ^ n37456;
  assign n41815 = n41814 ^ n37449;
  assign n41826 = n41825 ^ n41815;
  assign n41828 = n41827 ^ n41826;
  assign n41808 = n39542 ^ n30939;
  assign n41809 = n41808 ^ n35583;
  assign n41810 = n41809 ^ n2499;
  assign n41774 = n41773 ^ n41764;
  assign n2370 = n2369 ^ n2345;
  assign n2398 = n2397 ^ n2370;
  assign n2405 = n2404 ^ n2398;
  assign n41775 = n41774 ^ n2405;
  assign n41777 = n39549 ^ n30805;
  assign n41778 = n41777 ^ n35590;
  assign n41779 = n41778 ^ n2389;
  assign n41776 = n41772 ^ n41771;
  assign n41780 = n41779 ^ n41776;
  assign n41782 = n2302 ^ n1353;
  assign n41783 = n41782 ^ n35595;
  assign n41784 = n41783 ^ n29264;
  assign n41781 = n41770 ^ n41769;
  assign n41785 = n41784 ^ n41781;
  assign n41786 = n41768 ^ n41765;
  assign n1292 = n1252 ^ n1198;
  assign n1293 = n1292 ^ n1289;
  assign n1300 = n1299 ^ n1293;
  assign n41787 = n41786 ^ n1300;
  assign n41788 = n41767 ^ n41766;
  assign n1256 = n1237 ^ n1180;
  assign n1275 = n1274 ^ n1256;
  assign n1282 = n1281 ^ n1275;
  assign n41789 = n41788 ^ n1282;
  assign n41591 = n41590 ^ n41574;
  assign n41382 = n39138 ^ n1089;
  assign n41383 = n41382 ^ n35609;
  assign n41384 = n41383 ^ n29275;
  assign n41381 = n41380 ^ n41335;
  assign n41385 = n41384 ^ n41381;
  assign n41389 = n41379 ^ n41378;
  assign n41390 = n41389 ^ n41388;
  assign n41392 = n39148 ^ n30693;
  assign n41393 = n41392 ^ n35619;
  assign n41394 = n41393 ^ n773;
  assign n41391 = n41377 ^ n41336;
  assign n41395 = n41394 ^ n41391;
  assign n41399 = n41376 ^ n41337;
  assign n41396 = n39307 ^ n30688;
  assign n41397 = n41396 ^ n707;
  assign n41398 = n41397 ^ n29282;
  assign n41400 = n41399 ^ n41398;
  assign n41402 = n39153 ^ n30717;
  assign n41403 = n41402 ^ n35625;
  assign n41404 = n41403 ^ n699;
  assign n41401 = n41375 ^ n41374;
  assign n41405 = n41404 ^ n41401;
  assign n41551 = n41373 ^ n41372;
  assign n41409 = n41371 ^ n41370;
  assign n41406 = n39157 ^ n30712;
  assign n41407 = n41406 ^ n35636;
  assign n41408 = n41407 ^ n29294;
  assign n41410 = n41409 ^ n41408;
  assign n41411 = n41369 ^ n41368;
  assign n41415 = n41414 ^ n41411;
  assign n41537 = n41367 ^ n41338;
  assign n41419 = n41366 ^ n41365;
  assign n41416 = n39279 ^ n30573;
  assign n41417 = n41416 ^ n35650;
  assign n41418 = n41417 ^ n29309;
  assign n41420 = n41419 ^ n41418;
  assign n41526 = n41364 ^ n41340;
  assign n41422 = n39178 ^ n2262;
  assign n41423 = n41422 ^ n35661;
  assign n41424 = n41423 ^ n29319;
  assign n41421 = n41363 ^ n41362;
  assign n41425 = n41424 ^ n41421;
  assign n41515 = n41361 ^ n41360;
  assign n41507 = n41359 ^ n41358;
  assign n41427 = n39193 ^ n30594;
  assign n41428 = n41427 ^ n1847;
  assign n41429 = n41428 ^ n28866;
  assign n41426 = n41357 ^ n41341;
  assign n41430 = n41429 ^ n41426;
  assign n41434 = n41356 ^ n41355;
  assign n41431 = n39256 ^ n30589;
  assign n41432 = n41431 ^ n35677;
  assign n41433 = n41432 ^ n1839;
  assign n41435 = n41434 ^ n41433;
  assign n41496 = n41354 ^ n41342;
  assign n41439 = n41353 ^ n41344;
  assign n41436 = n39199 ^ n30608;
  assign n41437 = n41436 ^ n35684;
  assign n41438 = n41437 ^ n1729;
  assign n41440 = n41439 ^ n41438;
  assign n41444 = n41352 ^ n41351;
  assign n41445 = n41444 ^ n41443;
  assign n41447 = n39210 ^ n30613;
  assign n41448 = n41447 ^ n35056;
  assign n41449 = n41448 ^ n28799;
  assign n41446 = n41350 ^ n41345;
  assign n41450 = n41449 ^ n41446;
  assign n41451 = n41349 ^ n41346;
  assign n41455 = n41454 ^ n41451;
  assign n41457 = n39214 ^ n30634;
  assign n41458 = n41457 ^ n35065;
  assign n41459 = n41458 ^ n28807;
  assign n41456 = n41348 ^ n41347;
  assign n41460 = n41459 ^ n41456;
  assign n41461 = n39218 ^ n30626;
  assign n41462 = n41461 ^ n35069;
  assign n41463 = n41462 ^ n28816;
  assign n41464 = n41463 ^ n41347;
  assign n41475 = n41474 ^ n41472;
  assign n41476 = n41473 & ~n41475;
  assign n41477 = n41476 ^ n41469;
  assign n41478 = n41477 ^ n41347;
  assign n41479 = n41464 & ~n41478;
  assign n41480 = n41479 ^ n41463;
  assign n41481 = n41480 ^ n41456;
  assign n41482 = n41460 & ~n41481;
  assign n41483 = n41482 ^ n41459;
  assign n41484 = n41483 ^ n41451;
  assign n41485 = ~n41455 & n41484;
  assign n41486 = n41485 ^ n41454;
  assign n41487 = n41486 ^ n41446;
  assign n41488 = ~n41450 & n41487;
  assign n41489 = n41488 ^ n41449;
  assign n41490 = n41489 ^ n41444;
  assign n41491 = ~n41445 & n41490;
  assign n41492 = n41491 ^ n41443;
  assign n41493 = n41492 ^ n41439;
  assign n41494 = n41440 & ~n41493;
  assign n41495 = n41494 ^ n41438;
  assign n41497 = n41496 ^ n41495;
  assign n1710 = n1709 ^ n1685;
  assign n1738 = n1737 ^ n1710;
  assign n1745 = n1744 ^ n1738;
  assign n41498 = n41496 ^ n1745;
  assign n41499 = ~n41497 & n41498;
  assign n41500 = n41499 ^ n1745;
  assign n41501 = n41500 ^ n41434;
  assign n41502 = n41435 & ~n41501;
  assign n41503 = n41502 ^ n41433;
  assign n41504 = n41503 ^ n41426;
  assign n41505 = n41430 & ~n41504;
  assign n41506 = n41505 ^ n41429;
  assign n41508 = n41507 ^ n41506;
  assign n41512 = n41511 ^ n41507;
  assign n41513 = n41508 & ~n41512;
  assign n41514 = n41513 ^ n41511;
  assign n41516 = n41515 ^ n41514;
  assign n41517 = n39183 ^ n2244;
  assign n41518 = n41517 ^ n35666;
  assign n41519 = n41518 ^ n29324;
  assign n41520 = n41519 ^ n41515;
  assign n41521 = n41516 & ~n41520;
  assign n41522 = n41521 ^ n41519;
  assign n41523 = n41522 ^ n41421;
  assign n41524 = ~n41425 & n41523;
  assign n41525 = n41524 ^ n41424;
  assign n41527 = n41526 ^ n41525;
  assign n41531 = n41530 ^ n41526;
  assign n41532 = ~n41527 & n41531;
  assign n41533 = n41532 ^ n41530;
  assign n41534 = n41533 ^ n41419;
  assign n41535 = ~n41420 & n41534;
  assign n41536 = n41535 ^ n41418;
  assign n41538 = n41537 ^ n41536;
  assign n41539 = n39168 ^ n30568;
  assign n41540 = n41539 ^ n35646;
  assign n41541 = n41540 ^ n29304;
  assign n41542 = n41541 ^ n41537;
  assign n41543 = n41538 & ~n41542;
  assign n41544 = n41543 ^ n41541;
  assign n41545 = n41544 ^ n41411;
  assign n41546 = n41415 & ~n41545;
  assign n41547 = n41546 ^ n41414;
  assign n41548 = n41547 ^ n41409;
  assign n41549 = ~n41410 & n41548;
  assign n41550 = n41549 ^ n41408;
  assign n41552 = n41551 ^ n41550;
  assign n41553 = n39296 ^ n662;
  assign n41554 = n41553 ^ n35631;
  assign n41555 = n41554 ^ n29289;
  assign n41556 = n41555 ^ n41551;
  assign n41557 = n41552 & ~n41556;
  assign n41558 = n41557 ^ n41555;
  assign n41559 = n41558 ^ n41401;
  assign n41560 = ~n41405 & n41559;
  assign n41561 = n41560 ^ n41404;
  assign n41562 = n41561 ^ n41399;
  assign n41563 = ~n41400 & n41562;
  assign n41564 = n41563 ^ n41398;
  assign n41565 = n41564 ^ n41391;
  assign n41566 = ~n41395 & n41565;
  assign n41567 = n41566 ^ n41394;
  assign n41568 = n41567 ^ n41389;
  assign n41569 = ~n41390 & n41568;
  assign n41570 = n41569 ^ n41388;
  assign n41571 = n41570 ^ n41381;
  assign n41572 = ~n41385 & n41571;
  assign n41573 = n41572 ^ n41384;
  assign n41592 = n41591 ^ n41573;
  assign n41790 = n41595 ^ n41591;
  assign n41791 = ~n41592 & n41790;
  assign n41792 = n41791 ^ n41595;
  assign n41793 = n41792 ^ n41788;
  assign n41794 = n41789 & ~n41793;
  assign n41795 = n41794 ^ n1282;
  assign n41796 = n41795 ^ n41786;
  assign n41797 = ~n41787 & n41796;
  assign n41798 = n41797 ^ n1300;
  assign n41799 = n41798 ^ n41781;
  assign n41800 = n41785 & ~n41799;
  assign n41801 = n41800 ^ n41784;
  assign n41802 = n41801 ^ n41776;
  assign n41803 = ~n41780 & n41802;
  assign n41804 = n41803 ^ n41779;
  assign n41805 = n41804 ^ n41774;
  assign n41806 = n41775 & ~n41805;
  assign n41807 = n41806 ^ n2405;
  assign n41811 = n41810 ^ n41807;
  assign n41829 = n41828 ^ n41811;
  assign n41690 = n40050 ^ n39392;
  assign n41691 = n40740 ^ n40050;
  assign n41692 = n41690 & ~n41691;
  assign n41693 = n41692 ^ n39392;
  assign n41830 = n41829 ^ n41693;
  assign n41832 = n40056 ^ n39398;
  assign n41833 = n40746 ^ n40056;
  assign n41834 = ~n41832 & ~n41833;
  assign n41835 = n41834 ^ n39398;
  assign n41831 = n41804 ^ n41775;
  assign n41836 = n41835 ^ n41831;
  assign n41841 = n41801 ^ n41780;
  assign n41837 = n40058 ^ n39404;
  assign n41838 = n40752 ^ n40058;
  assign n41839 = ~n41837 & ~n41838;
  assign n41840 = n41839 ^ n39404;
  assign n41842 = n41841 ^ n41840;
  assign n41844 = n40064 ^ n39410;
  assign n41845 = n40753 ^ n40064;
  assign n41846 = ~n41844 & n41845;
  assign n41847 = n41846 ^ n39410;
  assign n41843 = n41798 ^ n41785;
  assign n41848 = n41847 ^ n41843;
  assign n41849 = n40070 ^ n39420;
  assign n41850 = n40763 ^ n40070;
  assign n41851 = ~n41849 & ~n41850;
  assign n41852 = n41851 ^ n39420;
  assign n41853 = n41795 ^ n41787;
  assign n41854 = ~n41852 & ~n41853;
  assign n41855 = n41854 ^ n41843;
  assign n41856 = ~n41848 & n41855;
  assign n41857 = n41856 ^ n41854;
  assign n41858 = n41857 ^ n41841;
  assign n41859 = ~n41842 & n41858;
  assign n41860 = n41859 ^ n41840;
  assign n41861 = n41860 ^ n41831;
  assign n41862 = n41836 & ~n41861;
  assign n41863 = n41862 ^ n41835;
  assign n41864 = n41863 ^ n41829;
  assign n41865 = ~n41830 & ~n41864;
  assign n41866 = n41865 ^ n41693;
  assign n41867 = n41866 ^ n41684;
  assign n41868 = n41689 & n41867;
  assign n41869 = n41868 ^ n41688;
  assign n41870 = n41869 ^ n41678;
  assign n41871 = ~n41683 & ~n41870;
  assign n41872 = n41871 ^ n41682;
  assign n41673 = n40032 ^ n39374;
  assign n41674 = n40726 ^ n40032;
  assign n41675 = ~n41673 & ~n41674;
  assign n41676 = n41675 ^ n39374;
  assign n41672 = n41477 ^ n41464;
  assign n41677 = n41676 ^ n41672;
  assign n41950 = n41872 ^ n41677;
  assign n41951 = n41950 ^ n38418;
  assign n41952 = n41869 ^ n41682;
  assign n41953 = n41952 ^ n41678;
  assign n41954 = n41953 ^ n38425;
  assign n41955 = n41866 ^ n41689;
  assign n41956 = n41955 ^ n38432;
  assign n41957 = n41863 ^ n41830;
  assign n41958 = n41957 ^ n38444;
  assign n41959 = n41860 ^ n41835;
  assign n41960 = n41959 ^ n41831;
  assign n41961 = n41960 ^ n38904;
  assign n41962 = n41857 ^ n41842;
  assign n41963 = n41962 ^ n38450;
  assign n41964 = n41853 ^ n41852;
  assign n41965 = n38458 & n41964;
  assign n41966 = n41965 ^ n38456;
  assign n41967 = n41854 ^ n41847;
  assign n41968 = n41967 ^ n41843;
  assign n41969 = n41968 ^ n41965;
  assign n41970 = n41966 & ~n41969;
  assign n41971 = n41970 ^ n38456;
  assign n41972 = n41971 ^ n41962;
  assign n41973 = n41963 & n41972;
  assign n41974 = n41973 ^ n38450;
  assign n41975 = n41974 ^ n41960;
  assign n41976 = ~n41961 & n41975;
  assign n41977 = n41976 ^ n38904;
  assign n41978 = n41977 ^ n41957;
  assign n41979 = n41958 & ~n41978;
  assign n41980 = n41979 ^ n38444;
  assign n41981 = n41980 ^ n41955;
  assign n41982 = ~n41956 & ~n41981;
  assign n41983 = n41982 ^ n38432;
  assign n41984 = n41983 ^ n41953;
  assign n41985 = ~n41954 & n41984;
  assign n41986 = n41985 ^ n38425;
  assign n41987 = n41986 ^ n41950;
  assign n41988 = ~n41951 & ~n41987;
  assign n41989 = n41988 ^ n38418;
  assign n41873 = n41872 ^ n41672;
  assign n41874 = ~n41677 & n41873;
  assign n41875 = n41874 ^ n41676;
  assign n41667 = n40386 ^ n39372;
  assign n41668 = n40720 ^ n40386;
  assign n41669 = ~n41667 & ~n41668;
  assign n41670 = n41669 ^ n39372;
  assign n41947 = n41875 ^ n41670;
  assign n41665 = n41480 ^ n41459;
  assign n41666 = n41665 ^ n41456;
  assign n41948 = n41947 ^ n41666;
  assign n41949 = n41948 ^ n38411;
  assign n42045 = n41989 ^ n41949;
  assign n42046 = n41986 ^ n41951;
  assign n42047 = n41980 ^ n41956;
  assign n42048 = n41971 ^ n41963;
  assign n42049 = n41974 ^ n41961;
  assign n42050 = ~n42048 & ~n42049;
  assign n42051 = n41977 ^ n41958;
  assign n42052 = n42050 & n42051;
  assign n42053 = n42047 & ~n42052;
  assign n42054 = n41983 ^ n41954;
  assign n42055 = ~n42053 & n42054;
  assign n42056 = n42046 & n42055;
  assign n42057 = n42045 & ~n42056;
  assign n41990 = n41989 ^ n41948;
  assign n41991 = ~n41949 & ~n41990;
  assign n41992 = n41991 ^ n38411;
  assign n41671 = n41670 ^ n41666;
  assign n41876 = n41875 ^ n41666;
  assign n41877 = n41671 & n41876;
  assign n41878 = n41877 ^ n41670;
  assign n41659 = n40476 ^ n39362;
  assign n41660 = n40708 ^ n40476;
  assign n41661 = n41659 & n41660;
  assign n41662 = n41661 ^ n39362;
  assign n41944 = n41878 ^ n41662;
  assign n41663 = n41483 ^ n41455;
  assign n41945 = n41944 ^ n41663;
  assign n41946 = n41945 ^ n38404;
  assign n42058 = n41992 ^ n41946;
  assign n42059 = n42057 & n42058;
  assign n41993 = n41992 ^ n41945;
  assign n41994 = n41946 & n41993;
  assign n41995 = n41994 ^ n38404;
  assign n41664 = n41663 ^ n41662;
  assign n41879 = n41878 ^ n41663;
  assign n41880 = ~n41664 & n41879;
  assign n41881 = n41880 ^ n41662;
  assign n41653 = n40646 ^ n39360;
  assign n41654 = n40706 ^ n40646;
  assign n41655 = ~n41653 & ~n41654;
  assign n41656 = n41655 ^ n39360;
  assign n41941 = n41881 ^ n41656;
  assign n41657 = n41486 ^ n41450;
  assign n41942 = n41941 ^ n41657;
  assign n41943 = n41942 ^ n38397;
  assign n42060 = n41995 ^ n41943;
  assign n42061 = ~n42059 & n42060;
  assign n41996 = n41995 ^ n41942;
  assign n41997 = n41943 & n41996;
  assign n41998 = n41997 ^ n38397;
  assign n41658 = n41657 ^ n41656;
  assign n41882 = n41881 ^ n41657;
  assign n41883 = n41658 & n41882;
  assign n41884 = n41883 ^ n41656;
  assign n41648 = n40716 ^ n39354;
  assign n41649 = n40716 ^ n40699;
  assign n41650 = n41648 & n41649;
  assign n41651 = n41650 ^ n39354;
  assign n41938 = n41884 ^ n41651;
  assign n41647 = n41489 ^ n41445;
  assign n41939 = n41938 ^ n41647;
  assign n41940 = n41939 ^ n38390;
  assign n42062 = n41998 ^ n41940;
  assign n42063 = n42061 & ~n42062;
  assign n41999 = n41998 ^ n41939;
  assign n42000 = n41940 & n41999;
  assign n42001 = n42000 ^ n38390;
  assign n41652 = n41651 ^ n41647;
  assign n41885 = n41884 ^ n41647;
  assign n41886 = n41652 & ~n41885;
  assign n41887 = n41886 ^ n41651;
  assign n41642 = n40710 ^ n39348;
  assign n41643 = n40710 ^ n40687;
  assign n41644 = n41642 & ~n41643;
  assign n41645 = n41644 ^ n39348;
  assign n41935 = n41887 ^ n41645;
  assign n41641 = n41492 ^ n41440;
  assign n41936 = n41935 ^ n41641;
  assign n41937 = n41936 ^ n38383;
  assign n42044 = n42001 ^ n41937;
  assign n42217 = n42063 ^ n42044;
  assign n42134 = n42062 ^ n42061;
  assign n42135 = n42134 ^ n42133;
  assign n42136 = n42060 ^ n42059;
  assign n1933 = n1923 ^ n1881;
  assign n1958 = n1957 ^ n1933;
  assign n1965 = n1964 ^ n1958;
  assign n42137 = n42136 ^ n1965;
  assign n42141 = n42058 ^ n42057;
  assign n42138 = n39886 ^ n1810;
  assign n42139 = n42138 ^ n35963;
  assign n42140 = n42139 ^ n1949;
  assign n42142 = n42141 ^ n42140;
  assign n42200 = n42056 ^ n42045;
  assign n42143 = n42055 ^ n42046;
  assign n42147 = n42146 ^ n42143;
  assign n42148 = n42054 ^ n42053;
  assign n42152 = n42151 ^ n42148;
  assign n42154 = n39907 ^ n31240;
  assign n42155 = n42154 ^ n35984;
  assign n42156 = n42155 ^ n29666;
  assign n42153 = n42052 ^ n42047;
  assign n42157 = n42156 ^ n42153;
  assign n42159 = n39933 ^ n31245;
  assign n42160 = n42159 ^ n35988;
  assign n42161 = n42160 ^ n1562;
  assign n42158 = n42051 ^ n42050;
  assign n42162 = n42161 ^ n42158;
  assign n42180 = n42049 ^ n42048;
  assign n42163 = n39920 ^ n30874;
  assign n42164 = n42163 ^ n35999;
  assign n42165 = n42164 ^ n29679;
  assign n42166 = n42165 ^ n42048;
  assign n42169 = n39915 ^ n30869;
  assign n42170 = n42169 ^ n2620;
  assign n42171 = n42170 ^ n29674;
  assign n2581 = n2578 ^ n2532;
  assign n2603 = n2602 ^ n2581;
  assign n2610 = n2609 ^ n2603;
  assign n42167 = n41964 ^ n38458;
  assign n42168 = n2610 & n42167;
  assign n42172 = n42171 ^ n42168;
  assign n42173 = n41968 ^ n41966;
  assign n42174 = n42173 ^ n42171;
  assign n42175 = n42172 & ~n42174;
  assign n42176 = n42175 ^ n42168;
  assign n42177 = n42176 ^ n42048;
  assign n42178 = ~n42166 & n42177;
  assign n42179 = n42178 ^ n42165;
  assign n42181 = n42180 ^ n42179;
  assign n42182 = n39911 ^ n30865;
  assign n42183 = n42182 ^ n35993;
  assign n42184 = n42183 ^ n29671;
  assign n42185 = n42184 ^ n42180;
  assign n42186 = n42181 & ~n42185;
  assign n42187 = n42186 ^ n42184;
  assign n42188 = n42187 ^ n42158;
  assign n42189 = ~n42162 & n42188;
  assign n42190 = n42189 ^ n42161;
  assign n42191 = n42190 ^ n42153;
  assign n42192 = ~n42157 & n42191;
  assign n42193 = n42192 ^ n42156;
  assign n42194 = n42193 ^ n42148;
  assign n42195 = n42152 & ~n42194;
  assign n42196 = n42195 ^ n42151;
  assign n42197 = n42196 ^ n42143;
  assign n42198 = ~n42147 & n42197;
  assign n42199 = n42198 ^ n42146;
  assign n42201 = n42200 ^ n42199;
  assign n42202 = n39891 ^ n1795;
  assign n42203 = n42202 ^ n35969;
  assign n42204 = n42203 ^ n29656;
  assign n42205 = n42204 ^ n42200;
  assign n42206 = n42201 & ~n42205;
  assign n42207 = n42206 ^ n42204;
  assign n42208 = n42207 ^ n42141;
  assign n42209 = n42142 & ~n42208;
  assign n42210 = n42209 ^ n42140;
  assign n42211 = n42210 ^ n42136;
  assign n42212 = n42137 & ~n42211;
  assign n42213 = n42212 ^ n1965;
  assign n42214 = n42213 ^ n42134;
  assign n42215 = n42135 & ~n42214;
  assign n42216 = n42215 ^ n42133;
  assign n42218 = n42217 ^ n42216;
  assign n2088 = n2087 ^ n2021;
  assign n2104 = n2103 ^ n2088;
  assign n2111 = n2110 ^ n2104;
  assign n42219 = n42217 ^ n2111;
  assign n42220 = n42218 & ~n42219;
  assign n42221 = n42220 ^ n2111;
  assign n42002 = n42001 ^ n41936;
  assign n42003 = n41937 & n42002;
  assign n42004 = n42003 ^ n38383;
  assign n41646 = n41645 ^ n41641;
  assign n41888 = n41887 ^ n41641;
  assign n41889 = ~n41646 & n41888;
  assign n41890 = n41889 ^ n41645;
  assign n41639 = n41497 ^ n1745;
  assign n41635 = n40702 ^ n39683;
  assign n41636 = n40702 ^ n40680;
  assign n41637 = ~n41635 & n41636;
  assign n41638 = n41637 ^ n39683;
  assign n41640 = n41639 ^ n41638;
  assign n41933 = n41890 ^ n41640;
  assign n41934 = n41933 ^ n38376;
  assign n42065 = n42004 ^ n41934;
  assign n42064 = n42044 & n42063;
  assign n42126 = n42065 ^ n42064;
  assign n42130 = n42129 ^ n42126;
  assign n42845 = n42221 ^ n42130;
  assign n41609 = n41522 ^ n41425;
  assign n43953 = n42845 ^ n41609;
  assign n42717 = n40534 ^ n2039;
  assign n42718 = n42717 ^ n36690;
  assign n42719 = n42718 ^ n30594;
  assign n42309 = n40708 ^ n40032;
  assign n42310 = n42309 ^ n41641;
  assign n42308 = n42176 ^ n42166;
  assign n42311 = n42310 ^ n42308;
  assign n42313 = n41647 ^ n40720;
  assign n42314 = n42313 ^ n40038;
  assign n42312 = n42173 ^ n42172;
  assign n42315 = n42314 ^ n42312;
  assign n42318 = n42167 ^ n2610;
  assign n42316 = n40726 ^ n40040;
  assign n42317 = n42316 ^ n41657;
  assign n42319 = n42318 ^ n42317;
  assign n42405 = n40314 ^ n39596;
  assign n42406 = n41104 ^ n40314;
  assign n42407 = n42405 & ~n42406;
  assign n42408 = n42407 ^ n39596;
  assign n42404 = n41570 ^ n41385;
  assign n42409 = n42408 ^ n42404;
  assign n42362 = n40320 ^ n39598;
  assign n42363 = n41110 ^ n40320;
  assign n42364 = n42362 & ~n42363;
  assign n42365 = n42364 ^ n39598;
  assign n42288 = n41567 ^ n41390;
  assign n42400 = n42365 ^ n42288;
  assign n42326 = n41564 ^ n41395;
  assign n42322 = n40326 ^ n39608;
  assign n42323 = n41112 ^ n40326;
  assign n42324 = ~n42322 & n42323;
  assign n42325 = n42324 ^ n39608;
  assign n42327 = n42326 ^ n42325;
  assign n42332 = n41561 ^ n41400;
  assign n42328 = n40332 ^ n39621;
  assign n42329 = n41824 ^ n40332;
  assign n42330 = ~n42328 & ~n42329;
  assign n42331 = n42330 ^ n39621;
  assign n42333 = n42332 ^ n42331;
  assign n42338 = n41558 ^ n41405;
  assign n42334 = n40338 ^ n39618;
  assign n42335 = n41597 ^ n40338;
  assign n42336 = n42334 & n42335;
  assign n42337 = n42336 ^ n39618;
  assign n42339 = n42338 ^ n42337;
  assign n42344 = n41555 ^ n41552;
  assign n42340 = n41087 ^ n40303;
  assign n42341 = n41728 ^ n41087;
  assign n42342 = n42340 & n42341;
  assign n42343 = n42342 ^ n40303;
  assign n42345 = n42344 ^ n42343;
  assign n42280 = n41547 ^ n41410;
  assign n42275 = n40968 ^ n40208;
  assign n42276 = n41698 ^ n40968;
  assign n42277 = ~n42275 & ~n42276;
  assign n42278 = n42277 ^ n40208;
  assign n42346 = n42280 ^ n42278;
  assign n42092 = n41544 ^ n41415;
  assign n42038 = n41541 ^ n41538;
  assign n42033 = n40914 ^ n40096;
  assign n42034 = n41710 ^ n40914;
  assign n42035 = ~n42033 & ~n42034;
  assign n42036 = n42035 ^ n40096;
  assign n42088 = n42038 ^ n42036;
  assign n41917 = n41533 ^ n41420;
  assign n41912 = n40102 ^ n40024;
  assign n41913 = n41582 ^ n40024;
  assign n41914 = n41912 & n41913;
  assign n41915 = n41914 ^ n40102;
  assign n42029 = n41917 ^ n41915;
  assign n41603 = n41530 ^ n41527;
  assign n41599 = n40661 ^ n40108;
  assign n41600 = n41332 ^ n40661;
  assign n41601 = ~n41599 & n41600;
  assign n41602 = n41601 ^ n40108;
  assign n41604 = n41603 ^ n41602;
  assign n41605 = n40668 ^ n40114;
  assign n41606 = n41189 ^ n40668;
  assign n41607 = n41605 & ~n41606;
  assign n41608 = n41607 ^ n40114;
  assign n41610 = n41609 ^ n41608;
  assign n41615 = n41519 ^ n41516;
  assign n41611 = n40675 ^ n40120;
  assign n41612 = n40675 ^ n40656;
  assign n41613 = n41611 & n41612;
  assign n41614 = n41613 ^ n40120;
  assign n41616 = n41615 ^ n41614;
  assign n41618 = n40682 ^ n40122;
  assign n41619 = n40682 ^ n40659;
  assign n41620 = n41618 & n41619;
  assign n41621 = n41620 ^ n40122;
  assign n41617 = n41511 ^ n41508;
  assign n41622 = n41621 ^ n41617;
  assign n41627 = n41503 ^ n41430;
  assign n41623 = n40689 ^ n40018;
  assign n41624 = n40689 ^ n40666;
  assign n41625 = ~n41623 & ~n41624;
  assign n41626 = n41625 ^ n40018;
  assign n41628 = n41627 ^ n41626;
  assign n41630 = n40695 ^ n39798;
  assign n41631 = n40695 ^ n40673;
  assign n41632 = ~n41630 & ~n41631;
  assign n41633 = n41632 ^ n39798;
  assign n41629 = n41500 ^ n41435;
  assign n41634 = n41633 ^ n41629;
  assign n41891 = n41890 ^ n41639;
  assign n41892 = ~n41640 & n41891;
  assign n41893 = n41892 ^ n41638;
  assign n41894 = n41893 ^ n41629;
  assign n41895 = n41634 & n41894;
  assign n41896 = n41895 ^ n41633;
  assign n41897 = n41896 ^ n41627;
  assign n41898 = ~n41628 & ~n41897;
  assign n41899 = n41898 ^ n41626;
  assign n41900 = n41899 ^ n41617;
  assign n41901 = n41622 & ~n41900;
  assign n41902 = n41901 ^ n41621;
  assign n41903 = n41902 ^ n41615;
  assign n41904 = n41616 & ~n41903;
  assign n41905 = n41904 ^ n41614;
  assign n41906 = n41905 ^ n41609;
  assign n41907 = ~n41610 & ~n41906;
  assign n41908 = n41907 ^ n41608;
  assign n41909 = n41908 ^ n41603;
  assign n41910 = n41604 & ~n41909;
  assign n41911 = n41910 ^ n41602;
  assign n42030 = n41917 ^ n41911;
  assign n42031 = ~n42029 & n42030;
  assign n42032 = n42031 ^ n41915;
  assign n42089 = n42038 ^ n42032;
  assign n42090 = n42088 & n42089;
  assign n42091 = n42090 ^ n42036;
  assign n42093 = n42092 ^ n42091;
  assign n42084 = n40952 ^ n39341;
  assign n42085 = n41704 ^ n40952;
  assign n42086 = n42084 & n42085;
  assign n42087 = n42086 ^ n39341;
  assign n42272 = n42092 ^ n42087;
  assign n42273 = n42093 & ~n42272;
  assign n42274 = n42273 ^ n42087;
  assign n42347 = n42280 ^ n42274;
  assign n42348 = ~n42346 & ~n42347;
  assign n42349 = n42348 ^ n42278;
  assign n42350 = n42349 ^ n42344;
  assign n42351 = n42345 & n42350;
  assign n42352 = n42351 ^ n42343;
  assign n42353 = n42352 ^ n42338;
  assign n42354 = n42339 & ~n42353;
  assign n42355 = n42354 ^ n42337;
  assign n42356 = n42355 ^ n42332;
  assign n42357 = n42333 & ~n42356;
  assign n42358 = n42357 ^ n42331;
  assign n42359 = n42358 ^ n42326;
  assign n42360 = n42327 & ~n42359;
  assign n42361 = n42360 ^ n42325;
  assign n42401 = n42361 ^ n42288;
  assign n42402 = n42400 & ~n42401;
  assign n42403 = n42402 ^ n42365;
  assign n42410 = n42409 ^ n42403;
  assign n42411 = n42410 ^ n38846;
  assign n42366 = n42365 ^ n42361;
  assign n42367 = n42366 ^ n42288;
  assign n42368 = n42367 ^ n38852;
  assign n42369 = n42358 ^ n42325;
  assign n42370 = n42369 ^ n42326;
  assign n42371 = n42370 ^ n38858;
  assign n42372 = n42355 ^ n42331;
  assign n42373 = n42372 ^ n42332;
  assign n42374 = n42373 ^ n38864;
  assign n42375 = n42352 ^ n42337;
  assign n42376 = n42375 ^ n42338;
  assign n42377 = n42376 ^ n38870;
  assign n42378 = n42349 ^ n42343;
  assign n42379 = n42378 ^ n42344;
  assign n42380 = n42379 ^ n39587;
  assign n42279 = n42278 ^ n42274;
  assign n42281 = n42280 ^ n42279;
  assign n42381 = n42281 ^ n39534;
  assign n42094 = n42093 ^ n42087;
  assign n42267 = n42094 ^ n39342;
  assign n42037 = n42036 ^ n42032;
  assign n42039 = n42038 ^ n42037;
  assign n42040 = n42039 ^ n39495;
  assign n41916 = n41915 ^ n41911;
  assign n41918 = n41917 ^ n41916;
  assign n41919 = n41918 ^ n39467;
  assign n41920 = n41908 ^ n41604;
  assign n41921 = n41920 ^ n39445;
  assign n41922 = n41905 ^ n41610;
  assign n41923 = n41922 ^ n39447;
  assign n41924 = n41902 ^ n41616;
  assign n41925 = n41924 ^ n39331;
  assign n41926 = n41899 ^ n41621;
  assign n41927 = n41926 ^ n41617;
  assign n41928 = n41927 ^ n39126;
  assign n41929 = n41896 ^ n41628;
  assign n41930 = n41929 ^ n39068;
  assign n41931 = n41893 ^ n41634;
  assign n41932 = n41931 ^ n38947;
  assign n42005 = n42004 ^ n41933;
  assign n42006 = ~n41934 & ~n42005;
  assign n42007 = n42006 ^ n38376;
  assign n42008 = n42007 ^ n41931;
  assign n42009 = ~n41932 & ~n42008;
  assign n42010 = n42009 ^ n38947;
  assign n42011 = n42010 ^ n41929;
  assign n42012 = n41930 & n42011;
  assign n42013 = n42012 ^ n39068;
  assign n42014 = n42013 ^ n41927;
  assign n42015 = ~n41928 & ~n42014;
  assign n42016 = n42015 ^ n39126;
  assign n42017 = n42016 ^ n41924;
  assign n42018 = n41925 & n42017;
  assign n42019 = n42018 ^ n39331;
  assign n42020 = n42019 ^ n41922;
  assign n42021 = ~n41923 & n42020;
  assign n42022 = n42021 ^ n39447;
  assign n42023 = n42022 ^ n41920;
  assign n42024 = n41921 & n42023;
  assign n42025 = n42024 ^ n39445;
  assign n42026 = n42025 ^ n41918;
  assign n42027 = n41919 & n42026;
  assign n42028 = n42027 ^ n39467;
  assign n42080 = n42039 ^ n42028;
  assign n42081 = ~n42040 & n42080;
  assign n42082 = n42081 ^ n39495;
  assign n42268 = n42094 ^ n42082;
  assign n42269 = n42267 & n42268;
  assign n42270 = n42269 ^ n39342;
  assign n42382 = n42281 ^ n42270;
  assign n42383 = ~n42381 & ~n42382;
  assign n42384 = n42383 ^ n39534;
  assign n42385 = n42384 ^ n42379;
  assign n42386 = ~n42380 & n42385;
  assign n42387 = n42386 ^ n39587;
  assign n42388 = n42387 ^ n42376;
  assign n42389 = n42377 & ~n42388;
  assign n42390 = n42389 ^ n38870;
  assign n42391 = n42390 ^ n42373;
  assign n42392 = n42374 & ~n42391;
  assign n42393 = n42392 ^ n38864;
  assign n42394 = n42393 ^ n42370;
  assign n42395 = n42371 & ~n42394;
  assign n42396 = n42395 ^ n38858;
  assign n42397 = n42396 ^ n42367;
  assign n42398 = ~n42368 & ~n42397;
  assign n42399 = n42398 ^ n38852;
  assign n42412 = n42411 ^ n42399;
  assign n42413 = n42384 ^ n42380;
  assign n42271 = n42270 ^ n39534;
  assign n42282 = n42281 ^ n42271;
  assign n42041 = n42040 ^ n42028;
  assign n42042 = n42010 ^ n41930;
  assign n42043 = n42007 ^ n41932;
  assign n42066 = n42064 & n42065;
  assign n42067 = n42043 & ~n42066;
  assign n42068 = ~n42042 & ~n42067;
  assign n42069 = n42013 ^ n41928;
  assign n42070 = n42068 & ~n42069;
  assign n42071 = n42016 ^ n41925;
  assign n42072 = n42070 & ~n42071;
  assign n42073 = n42019 ^ n41923;
  assign n42074 = ~n42072 & n42073;
  assign n42075 = n42022 ^ n41921;
  assign n42076 = ~n42074 & n42075;
  assign n42077 = n42025 ^ n41919;
  assign n42078 = n42076 & ~n42077;
  assign n42079 = n42041 & ~n42078;
  assign n42083 = n42082 ^ n39342;
  assign n42095 = n42094 ^ n42083;
  assign n42283 = n42079 & ~n42095;
  assign n42414 = ~n42282 & n42283;
  assign n42415 = ~n42413 & ~n42414;
  assign n42416 = n42387 ^ n42377;
  assign n42417 = n42415 & n42416;
  assign n42418 = n42390 ^ n42374;
  assign n42419 = n42417 & n42418;
  assign n42420 = n42393 ^ n42371;
  assign n42421 = n42419 & n42420;
  assign n42422 = n42396 ^ n42368;
  assign n42423 = ~n42421 & n42422;
  assign n42478 = n42412 & n42423;
  assign n42486 = n42404 ^ n42403;
  assign n42487 = n42409 & ~n42486;
  assign n42488 = n42487 ^ n42408;
  assign n41596 = n41595 ^ n41592;
  assign n42489 = n42488 ^ n41596;
  assign n42482 = n40082 ^ n39428;
  assign n42483 = n41094 ^ n40082;
  assign n42484 = ~n42482 & n42483;
  assign n42485 = n42484 ^ n39428;
  assign n42490 = n42489 ^ n42485;
  assign n42491 = n42490 ^ n38469;
  assign n42479 = n42410 ^ n42399;
  assign n42480 = n42411 & n42479;
  assign n42481 = n42480 ^ n38846;
  assign n42492 = n42491 ^ n42481;
  assign n42540 = n42478 & ~n42492;
  assign n42537 = n41792 ^ n41789;
  assign n42532 = n40076 ^ n39426;
  assign n42533 = n41092 ^ n40076;
  assign n42534 = ~n42532 & ~n42533;
  assign n42535 = n42534 ^ n39426;
  assign n42529 = n42485 ^ n41596;
  assign n42530 = n42489 & ~n42529;
  assign n42531 = n42530 ^ n42485;
  assign n42536 = n42535 ^ n42531;
  assign n42538 = n42537 ^ n42536;
  assign n42525 = n42490 ^ n42481;
  assign n42526 = n42491 & n42525;
  assign n42527 = n42526 ^ n38469;
  assign n42528 = n42527 ^ n38463;
  assign n42539 = n42538 ^ n42528;
  assign n42541 = n42540 ^ n42539;
  assign n42521 = n40231 ^ n2467;
  assign n42522 = n42521 ^ n36404;
  assign n42523 = n42522 ^ n2600;
  assign n42493 = n42492 ^ n42478;
  assign n42475 = n40235 ^ n2459;
  assign n42476 = n42475 ^ n36408;
  assign n42477 = n42476 ^ n30091;
  assign n42494 = n42493 ^ n42477;
  assign n42425 = n40241 ^ n31594;
  assign n42426 = n42425 ^ n36414;
  assign n42427 = n42426 ^ n30096;
  assign n42424 = n42423 ^ n42412;
  assign n42428 = n42427 ^ n42424;
  assign n42464 = n42422 ^ n42421;
  assign n42456 = n42420 ^ n42419;
  assign n42429 = n42418 ^ n42417;
  assign n42433 = n42432 ^ n42429;
  assign n42445 = n42416 ^ n42415;
  assign n42435 = n40260 ^ n31610;
  assign n42436 = n42435 ^ n36436;
  assign n42437 = n42436 ^ n969;
  assign n42434 = n42414 ^ n42413;
  assign n42438 = n42437 ^ n42434;
  assign n42284 = n42283 ^ n42282;
  assign n834 = n833 ^ n809;
  assign n862 = n861 ^ n834;
  assign n869 = n868 ^ n862;
  assign n42285 = n42284 ^ n869;
  assign n42097 = n39843 ^ n31617;
  assign n42098 = n42097 ^ n36443;
  assign n42099 = n42098 ^ n853;
  assign n42096 = n42095 ^ n42079;
  assign n42100 = n42099 ^ n42096;
  assign n42102 = n39999 ^ n751;
  assign n42103 = n42102 ^ n36448;
  assign n42104 = n42103 ^ n30119;
  assign n42101 = n42078 ^ n42041;
  assign n42105 = n42104 ^ n42101;
  assign n42107 = n39848 ^ n31624;
  assign n42108 = n42107 ^ n36453;
  assign n42109 = n42108 ^ n30137;
  assign n42106 = n42077 ^ n42076;
  assign n42110 = n42109 ^ n42106;
  assign n42112 = n39988 ^ n31629;
  assign n42113 = n42112 ^ n36458;
  assign n42114 = n42113 ^ n30124;
  assign n42111 = n42075 ^ n42074;
  assign n42115 = n42114 ^ n42111;
  assign n42247 = n42073 ^ n42072;
  assign n42119 = n42071 ^ n42070;
  assign n42116 = n39857 ^ n31192;
  assign n42117 = n42116 ^ n36489;
  assign n42118 = n42117 ^ n29762;
  assign n42120 = n42119 ^ n42118;
  assign n42236 = n42069 ^ n42068;
  assign n42121 = n42067 ^ n42042;
  assign n42125 = n42124 ^ n42121;
  assign n42225 = n42066 ^ n42043;
  assign n42222 = n42221 ^ n42126;
  assign n42223 = ~n42130 & n42222;
  assign n42224 = n42223 ^ n42129;
  assign n42226 = n42225 ^ n42224;
  assign n42227 = n39873 ^ n31207;
  assign n42228 = n42227 ^ n36040;
  assign n42229 = n42228 ^ n29641;
  assign n42230 = n42229 ^ n42225;
  assign n42231 = n42226 & ~n42230;
  assign n42232 = n42231 ^ n42229;
  assign n42233 = n42232 ^ n42121;
  assign n42234 = ~n42125 & n42233;
  assign n42235 = n42234 ^ n42124;
  assign n42237 = n42236 ^ n42235;
  assign n42241 = n42240 ^ n42236;
  assign n42242 = ~n42237 & n42241;
  assign n42243 = n42242 ^ n42240;
  assign n42244 = n42243 ^ n42119;
  assign n42245 = n42120 & ~n42244;
  assign n42246 = n42245 ^ n42118;
  assign n42248 = n42247 ^ n42246;
  assign n42249 = n39853 ^ n31634;
  assign n42250 = n42249 ^ n36463;
  assign n42251 = n42250 ^ n29768;
  assign n42252 = n42251 ^ n42247;
  assign n42253 = n42248 & ~n42252;
  assign n42254 = n42253 ^ n42251;
  assign n42255 = n42254 ^ n42111;
  assign n42256 = n42115 & ~n42255;
  assign n42257 = n42256 ^ n42114;
  assign n42258 = n42257 ^ n42106;
  assign n42259 = n42110 & ~n42258;
  assign n42260 = n42259 ^ n42109;
  assign n42261 = n42260 ^ n42101;
  assign n42262 = ~n42105 & n42261;
  assign n42263 = n42262 ^ n42104;
  assign n42264 = n42263 ^ n42096;
  assign n42265 = ~n42100 & n42264;
  assign n42266 = n42265 ^ n42099;
  assign n42439 = n42284 ^ n42266;
  assign n42440 = ~n42285 & n42439;
  assign n42441 = n42440 ^ n869;
  assign n42442 = n42441 ^ n42434;
  assign n42443 = ~n42438 & n42442;
  assign n42444 = n42443 ^ n42437;
  assign n42446 = n42445 ^ n42444;
  assign n42450 = n42449 ^ n42445;
  assign n42451 = n42446 & ~n42450;
  assign n42452 = n42451 ^ n42449;
  assign n42453 = n42452 ^ n42432;
  assign n42454 = ~n42433 & ~n42453;
  assign n42455 = n42454 ^ n42429;
  assign n42457 = n42456 ^ n42455;
  assign n42458 = n40245 ^ n1389;
  assign n42459 = n42458 ^ n36424;
  assign n42460 = n42459 ^ n30163;
  assign n42461 = n42460 ^ n42456;
  assign n42462 = ~n42457 & ~n42461;
  assign n42463 = n42462 ^ n42460;
  assign n42465 = n42464 ^ n42463;
  assign n42466 = n40282 ^ n1407;
  assign n42467 = n42466 ^ n36419;
  assign n42468 = n42467 ^ n30101;
  assign n42469 = n42468 ^ n42464;
  assign n42470 = n42465 & ~n42469;
  assign n42471 = n42470 ^ n42468;
  assign n42472 = n42471 ^ n42424;
  assign n42473 = n42428 & ~n42472;
  assign n42474 = n42473 ^ n42427;
  assign n42518 = n42493 ^ n42474;
  assign n42519 = ~n42494 & n42518;
  assign n42520 = n42519 ^ n42477;
  assign n42524 = n42523 ^ n42520;
  assign n42542 = n42541 ^ n42524;
  assign n42495 = n42494 ^ n42474;
  assign n42320 = n40738 ^ n40056;
  assign n42321 = n42320 ^ n41666;
  assign n42496 = n42495 ^ n42321;
  assign n42508 = n42471 ^ n42428;
  assign n42499 = n40752 ^ n40070;
  assign n42500 = n42499 ^ n41684;
  assign n42501 = n42460 ^ n42457;
  assign n42502 = ~n42500 & n42501;
  assign n42497 = n40746 ^ n40064;
  assign n42498 = n42497 ^ n41678;
  assign n42503 = n42502 ^ n42498;
  assign n42504 = n42468 ^ n42465;
  assign n42505 = n42504 ^ n42498;
  assign n42506 = n42503 & n42505;
  assign n42507 = n42506 ^ n42502;
  assign n42509 = n42508 ^ n42507;
  assign n42510 = n40740 ^ n40058;
  assign n42511 = n42510 ^ n41672;
  assign n42512 = n42511 ^ n42508;
  assign n42513 = ~n42509 & n42512;
  assign n42514 = n42513 ^ n42511;
  assign n42515 = n42514 ^ n42495;
  assign n42516 = ~n42496 & n42515;
  assign n42517 = n42516 ^ n42321;
  assign n42543 = n42542 ^ n42517;
  assign n42544 = n40732 ^ n40050;
  assign n42545 = n42544 ^ n41663;
  assign n42546 = n42545 ^ n42542;
  assign n42547 = ~n42543 & ~n42546;
  assign n42548 = n42547 ^ n42545;
  assign n42549 = n42548 ^ n42318;
  assign n42550 = n42319 & n42549;
  assign n42551 = n42550 ^ n42317;
  assign n42552 = n42551 ^ n42312;
  assign n42553 = n42315 & ~n42552;
  assign n42554 = n42553 ^ n42314;
  assign n42555 = n42554 ^ n42308;
  assign n42556 = n42311 & n42555;
  assign n42557 = n42556 ^ n42310;
  assign n42305 = n40706 ^ n40386;
  assign n42306 = n42305 ^ n41639;
  assign n42304 = n42184 ^ n42181;
  assign n42307 = n42306 ^ n42304;
  assign n42637 = n42557 ^ n42307;
  assign n42600 = n42554 ^ n42311;
  assign n42601 = n42600 ^ n39374;
  assign n42602 = n42551 ^ n42315;
  assign n42603 = n42602 ^ n39380;
  assign n42604 = n42548 ^ n42319;
  assign n42605 = n42604 ^ n39386;
  assign n42606 = n42545 ^ n42543;
  assign n42607 = n42606 ^ n39392;
  assign n42608 = n42514 ^ n42496;
  assign n42609 = n42608 ^ n39398;
  assign n42610 = n42511 ^ n42509;
  assign n42611 = n42610 ^ n39404;
  assign n42612 = n42501 ^ n42500;
  assign n42613 = ~n39420 & ~n42612;
  assign n42614 = n42613 ^ n39410;
  assign n42615 = n42504 ^ n42503;
  assign n42616 = n42615 ^ n42613;
  assign n42617 = n42614 & n42616;
  assign n42618 = n42617 ^ n39410;
  assign n42619 = n42618 ^ n42610;
  assign n42620 = n42611 & ~n42619;
  assign n42621 = n42620 ^ n39404;
  assign n42622 = n42621 ^ n42608;
  assign n42623 = ~n42609 & n42622;
  assign n42624 = n42623 ^ n39398;
  assign n42625 = n42624 ^ n42606;
  assign n42626 = n42607 & n42625;
  assign n42627 = n42626 ^ n39392;
  assign n42628 = n42627 ^ n42604;
  assign n42629 = ~n42605 & ~n42628;
  assign n42630 = n42629 ^ n39386;
  assign n42631 = n42630 ^ n42602;
  assign n42632 = ~n42603 & ~n42631;
  assign n42633 = n42632 ^ n39380;
  assign n42634 = n42633 ^ n42600;
  assign n42635 = ~n42601 & n42634;
  assign n42636 = n42635 ^ n39374;
  assign n42638 = n42637 ^ n42636;
  assign n42673 = n42638 ^ n39372;
  assign n42674 = n42633 ^ n42601;
  assign n42675 = n42621 ^ n42609;
  assign n42676 = n42615 ^ n42614;
  assign n42677 = n42618 ^ n42611;
  assign n42678 = n42676 & ~n42677;
  assign n42679 = ~n42675 & ~n42678;
  assign n42680 = n42624 ^ n42607;
  assign n42681 = ~n42679 & ~n42680;
  assign n42682 = n42627 ^ n42605;
  assign n42683 = ~n42681 & n42682;
  assign n42684 = n42630 ^ n42603;
  assign n42685 = ~n42683 & n42684;
  assign n42686 = ~n42674 & n42685;
  assign n42687 = ~n42673 & n42686;
  assign n42639 = n42637 ^ n39372;
  assign n42640 = ~n42638 & ~n42639;
  assign n42641 = n42640 ^ n39372;
  assign n42563 = n40699 ^ n40476;
  assign n42564 = n42563 ^ n41629;
  assign n42561 = n42187 ^ n42162;
  assign n42558 = n42557 ^ n42304;
  assign n42559 = n42307 & ~n42558;
  assign n42560 = n42559 ^ n42306;
  assign n42562 = n42561 ^ n42560;
  assign n42598 = n42564 ^ n42562;
  assign n42599 = n42598 ^ n39362;
  assign n42688 = n42641 ^ n42599;
  assign n42689 = ~n42687 & n42688;
  assign n42642 = n42641 ^ n42598;
  assign n42643 = n42599 & ~n42642;
  assign n42644 = n42643 ^ n39362;
  assign n42565 = n42564 ^ n42561;
  assign n42566 = ~n42562 & ~n42565;
  assign n42567 = n42566 ^ n42564;
  assign n42302 = n42190 ^ n42157;
  assign n42300 = n40687 ^ n40646;
  assign n42301 = n42300 ^ n41627;
  assign n42303 = n42302 ^ n42301;
  assign n42596 = n42567 ^ n42303;
  assign n42597 = n42596 ^ n39360;
  assign n42672 = n42644 ^ n42597;
  assign n42716 = n42689 ^ n42672;
  assign n42720 = n42719 ^ n42716;
  assign n42789 = n42688 ^ n42687;
  assign n42724 = n42686 ^ n42673;
  assign n42721 = n40538 ^ n31889;
  assign n42722 = n42721 ^ n36694;
  assign n42723 = n42722 ^ n1709;
  assign n42725 = n42724 ^ n42723;
  assign n42778 = n42685 ^ n42674;
  assign n42729 = n42684 ^ n42683;
  assign n42726 = n40548 ^ n31898;
  assign n42727 = n42726 ^ n36701;
  assign n42728 = n42727 ^ n1619;
  assign n42730 = n42729 ^ n42728;
  assign n42767 = n42682 ^ n42681;
  assign n42732 = n40580 ^ n31905;
  assign n42733 = n42732 ^ n36733;
  assign n42734 = n42733 ^ n30643;
  assign n42731 = n42680 ^ n42679;
  assign n42735 = n42734 ^ n42731;
  assign n42736 = n42678 ^ n42675;
  assign n42740 = n42739 ^ n42736;
  assign n42744 = n42677 ^ n42676;
  assign n42741 = n40562 ^ n31919;
  assign n42742 = n42741 ^ n36720;
  assign n42743 = n42742 ^ n30626;
  assign n42745 = n42744 ^ n42743;
  assign n42751 = n40565 ^ n31914;
  assign n42752 = n42751 ^ n36715;
  assign n42753 = n42752 ^ n30621;
  assign n42746 = n42612 ^ n39420;
  assign n42747 = n40771 ^ n32538;
  assign n42748 = n42747 ^ n37292;
  assign n42749 = n42748 ^ n30976;
  assign n42750 = n42746 & n42749;
  assign n42754 = n42753 ^ n42750;
  assign n42755 = n42750 ^ n42676;
  assign n42756 = n42754 & ~n42755;
  assign n42757 = n42756 ^ n42753;
  assign n42758 = n42757 ^ n42744;
  assign n42759 = n42745 & ~n42758;
  assign n42760 = n42759 ^ n42743;
  assign n42761 = n42760 ^ n42736;
  assign n42762 = n42740 & ~n42761;
  assign n42763 = n42762 ^ n42739;
  assign n42764 = n42763 ^ n42731;
  assign n42765 = ~n42735 & n42764;
  assign n42766 = n42765 ^ n42734;
  assign n42768 = n42767 ^ n42766;
  assign n42769 = n40553 ^ n1565;
  assign n42770 = n42769 ^ n36706;
  assign n42771 = n42770 ^ n30613;
  assign n42772 = n42771 ^ n42767;
  assign n42773 = n42768 & ~n42772;
  assign n42774 = n42773 ^ n42771;
  assign n42775 = n42774 ^ n42729;
  assign n42776 = n42730 & ~n42775;
  assign n42777 = n42776 ^ n42728;
  assign n42779 = n42778 ^ n42777;
  assign n42780 = n40544 ^ n31894;
  assign n42781 = n42780 ^ n1637;
  assign n42782 = n42781 ^ n30608;
  assign n42783 = n42782 ^ n42778;
  assign n42784 = ~n42779 & n42783;
  assign n42785 = n42784 ^ n42782;
  assign n42786 = n42785 ^ n42724;
  assign n42787 = n42725 & ~n42786;
  assign n42788 = n42787 ^ n42723;
  assign n42790 = n42789 ^ n42788;
  assign n42791 = n40600 ^ n31884;
  assign n42792 = n42791 ^ n36753;
  assign n42793 = n42792 ^ n30589;
  assign n42794 = n42793 ^ n42789;
  assign n42795 = n42790 & ~n42794;
  assign n42796 = n42795 ^ n42793;
  assign n42797 = n42796 ^ n42716;
  assign n42798 = ~n42720 & n42797;
  assign n42799 = n42798 ^ n42719;
  assign n42712 = n40529 ^ n2054;
  assign n42713 = n42712 ^ n36685;
  assign n42714 = n42713 ^ n2229;
  assign n42645 = n42644 ^ n42596;
  assign n42646 = ~n42597 & ~n42645;
  assign n42647 = n42646 ^ n39360;
  assign n42568 = n42567 ^ n42302;
  assign n42569 = n42303 & n42568;
  assign n42570 = n42569 ^ n42301;
  assign n42298 = n42193 ^ n42152;
  assign n42296 = n40716 ^ n40680;
  assign n42297 = n42296 ^ n41617;
  assign n42299 = n42298 ^ n42297;
  assign n42594 = n42570 ^ n42299;
  assign n42595 = n42594 ^ n39354;
  assign n42691 = n42647 ^ n42595;
  assign n42690 = ~n42672 & n42689;
  assign n42711 = n42691 ^ n42690;
  assign n42715 = n42714 ^ n42711;
  assign n43271 = n42799 ^ n42715;
  assign n43954 = n43953 ^ n43271;
  assign n42930 = n41110 ^ n40332;
  assign n42931 = n42930 ^ n42537;
  assign n42867 = n41112 ^ n40338;
  assign n42868 = n42867 ^ n41596;
  assign n42866 = n42257 ^ n42110;
  assign n42869 = n42868 ^ n42866;
  assign n42871 = n41824 ^ n41087;
  assign n42872 = n42871 ^ n42404;
  assign n42870 = n42254 ^ n42115;
  assign n42873 = n42872 ^ n42870;
  assign n42876 = n41728 ^ n40952;
  assign n42877 = n42876 ^ n42326;
  assign n42875 = n42243 ^ n42120;
  assign n42878 = n42877 ^ n42875;
  assign n42907 = n42240 ^ n42237;
  assign n42900 = n42232 ^ n42125;
  assign n42879 = n41710 ^ n40661;
  assign n42880 = n42879 ^ n42344;
  assign n42840 = n42229 ^ n42226;
  assign n42881 = n42880 ^ n42840;
  assign n42882 = n41332 ^ n40675;
  assign n42883 = n42882 ^ n42092;
  assign n42850 = n42218 ^ n2111;
  assign n42884 = n42883 ^ n42850;
  assign n42822 = n41189 ^ n40682;
  assign n42823 = n42822 ^ n42038;
  assign n42821 = n42213 ^ n42135;
  assign n42824 = n42823 ^ n42821;
  assign n42665 = n42210 ^ n42137;
  assign n42585 = n40695 ^ n40659;
  assign n42586 = n42585 ^ n41603;
  assign n42584 = n42207 ^ n42142;
  assign n42587 = n42586 ^ n42584;
  assign n42577 = n42204 ^ n42201;
  assign n42293 = n40710 ^ n40673;
  assign n42294 = n42293 ^ n41615;
  assign n42292 = n42196 ^ n42147;
  assign n42295 = n42294 ^ n42292;
  assign n42571 = n42570 ^ n42298;
  assign n42572 = ~n42299 & n42571;
  assign n42573 = n42572 ^ n42297;
  assign n42574 = n42573 ^ n42292;
  assign n42575 = n42295 & ~n42574;
  assign n42576 = n42575 ^ n42294;
  assign n42578 = n42577 ^ n42576;
  assign n42579 = n40702 ^ n40666;
  assign n42580 = n42579 ^ n41609;
  assign n42581 = n42580 ^ n42577;
  assign n42582 = ~n42578 & n42581;
  assign n42583 = n42582 ^ n42580;
  assign n42662 = n42584 ^ n42583;
  assign n42663 = ~n42587 & n42662;
  assign n42664 = n42663 ^ n42586;
  assign n42666 = n42665 ^ n42664;
  assign n42660 = n40689 ^ n40656;
  assign n42661 = n42660 ^ n41917;
  assign n42818 = n42665 ^ n42661;
  assign n42819 = n42666 & ~n42818;
  assign n42820 = n42819 ^ n42661;
  assign n42885 = n42821 ^ n42820;
  assign n42886 = n42824 & n42885;
  assign n42887 = n42886 ^ n42823;
  assign n42888 = n42887 ^ n42850;
  assign n42889 = n42884 & n42888;
  assign n42890 = n42889 ^ n42883;
  assign n42891 = n42890 ^ n42845;
  assign n42892 = n41582 ^ n40668;
  assign n42893 = n42892 ^ n42280;
  assign n42894 = n42893 ^ n42845;
  assign n42895 = ~n42891 & ~n42894;
  assign n42896 = n42895 ^ n42893;
  assign n42897 = n42896 ^ n42840;
  assign n42898 = ~n42881 & n42897;
  assign n42899 = n42898 ^ n42880;
  assign n42901 = n42900 ^ n42899;
  assign n42902 = n41704 ^ n40024;
  assign n42903 = n42902 ^ n42338;
  assign n42904 = n42903 ^ n42900;
  assign n42905 = n42901 & n42904;
  assign n42906 = n42905 ^ n42903;
  assign n42908 = n42907 ^ n42906;
  assign n42909 = n41698 ^ n40914;
  assign n42910 = n42909 ^ n42332;
  assign n42911 = n42910 ^ n42907;
  assign n42912 = n42908 & n42911;
  assign n42913 = n42912 ^ n42910;
  assign n42914 = n42913 ^ n42875;
  assign n42915 = n42878 & ~n42914;
  assign n42916 = n42915 ^ n42877;
  assign n42874 = n42251 ^ n42248;
  assign n42917 = n42916 ^ n42874;
  assign n42918 = n41597 ^ n40968;
  assign n42919 = n42918 ^ n42288;
  assign n42920 = n42919 ^ n42874;
  assign n42921 = n42917 & ~n42920;
  assign n42922 = n42921 ^ n42919;
  assign n42923 = n42922 ^ n42870;
  assign n42924 = n42873 & ~n42923;
  assign n42925 = n42924 ^ n42872;
  assign n42926 = n42925 ^ n42866;
  assign n42927 = n42869 & ~n42926;
  assign n42928 = n42927 ^ n42868;
  assign n42290 = n42260 ^ n42105;
  assign n42929 = n42928 ^ n42290;
  assign n42947 = n42931 ^ n42929;
  assign n42948 = n42947 ^ n39621;
  assign n42949 = n42925 ^ n42869;
  assign n42950 = n42949 ^ n39618;
  assign n42951 = n42922 ^ n42873;
  assign n42952 = n42951 ^ n40303;
  assign n42953 = n42919 ^ n42917;
  assign n42954 = n42953 ^ n40208;
  assign n42955 = n42913 ^ n42878;
  assign n42956 = n42955 ^ n39341;
  assign n42980 = n42910 ^ n42908;
  assign n42957 = n42903 ^ n42901;
  assign n42958 = n42957 ^ n40102;
  assign n42959 = n42896 ^ n42881;
  assign n42960 = n42959 ^ n40108;
  assign n42961 = n42893 ^ n42891;
  assign n42962 = n42961 ^ n40114;
  assign n42963 = n42887 ^ n42884;
  assign n42964 = n42963 ^ n40120;
  assign n42825 = n42824 ^ n42820;
  assign n42826 = n42825 ^ n40122;
  assign n42667 = n42666 ^ n42661;
  assign n42668 = n42667 ^ n40018;
  assign n42588 = n42587 ^ n42583;
  assign n42589 = n42588 ^ n39798;
  assign n42590 = n42580 ^ n42578;
  assign n42591 = n42590 ^ n39683;
  assign n42592 = n42573 ^ n42295;
  assign n42593 = n42592 ^ n39348;
  assign n42648 = n42647 ^ n42594;
  assign n42649 = ~n42595 & n42648;
  assign n42650 = n42649 ^ n39354;
  assign n42651 = n42650 ^ n42592;
  assign n42652 = n42593 & ~n42651;
  assign n42653 = n42652 ^ n39348;
  assign n42654 = n42653 ^ n42590;
  assign n42655 = n42591 & ~n42654;
  assign n42656 = n42655 ^ n39683;
  assign n42657 = n42656 ^ n42588;
  assign n42658 = n42589 & n42657;
  assign n42659 = n42658 ^ n39798;
  assign n42815 = n42667 ^ n42659;
  assign n42816 = ~n42668 & ~n42815;
  assign n42817 = n42816 ^ n40018;
  assign n42965 = n42825 ^ n42817;
  assign n42966 = n42826 & ~n42965;
  assign n42967 = n42966 ^ n40122;
  assign n42968 = n42967 ^ n42963;
  assign n42969 = ~n42964 & n42968;
  assign n42970 = n42969 ^ n40120;
  assign n42971 = n42970 ^ n42961;
  assign n42972 = n42962 & n42971;
  assign n42973 = n42972 ^ n40114;
  assign n42974 = n42973 ^ n42959;
  assign n42975 = ~n42960 & n42974;
  assign n42976 = n42975 ^ n40108;
  assign n42977 = n42976 ^ n42957;
  assign n42978 = n42958 & ~n42977;
  assign n42979 = n42978 ^ n40102;
  assign n42981 = n42980 ^ n42979;
  assign n42982 = n42980 ^ n40096;
  assign n42983 = n42981 & n42982;
  assign n42984 = n42983 ^ n40096;
  assign n42985 = n42984 ^ n42955;
  assign n42986 = ~n42956 & n42985;
  assign n42987 = n42986 ^ n39341;
  assign n42988 = n42987 ^ n42953;
  assign n42989 = ~n42954 & ~n42988;
  assign n42990 = n42989 ^ n40208;
  assign n42991 = n42990 ^ n42951;
  assign n42992 = ~n42952 & ~n42991;
  assign n42993 = n42992 ^ n40303;
  assign n42994 = n42993 ^ n42949;
  assign n42995 = ~n42950 & n42994;
  assign n42996 = n42995 ^ n39618;
  assign n42997 = n42996 ^ n42947;
  assign n42998 = ~n42948 & n42997;
  assign n42999 = n42998 ^ n39621;
  assign n42937 = n41104 ^ n40326;
  assign n42938 = n42937 ^ n41853;
  assign n42935 = n42263 ^ n42100;
  assign n42932 = n42931 ^ n42290;
  assign n42933 = n42929 & n42932;
  assign n42934 = n42933 ^ n42931;
  assign n42936 = n42935 ^ n42934;
  assign n42945 = n42938 ^ n42936;
  assign n42946 = n42945 ^ n39608;
  assign n43017 = n42999 ^ n42946;
  assign n43018 = n42993 ^ n42950;
  assign n43019 = n42987 ^ n42954;
  assign n43020 = n42981 ^ n40096;
  assign n43021 = n42970 ^ n42962;
  assign n43022 = n42967 ^ n42964;
  assign n42827 = n42826 ^ n42817;
  assign n42669 = n42668 ^ n42659;
  assign n42670 = n42653 ^ n42591;
  assign n42671 = n42650 ^ n42593;
  assign n42692 = n42690 & n42691;
  assign n42693 = ~n42671 & n42692;
  assign n42694 = ~n42670 & n42693;
  assign n42695 = n42656 ^ n42589;
  assign n42696 = ~n42694 & n42695;
  assign n42828 = n42669 & n42696;
  assign n43023 = ~n42827 & ~n42828;
  assign n43024 = ~n43022 & ~n43023;
  assign n43025 = ~n43021 & ~n43024;
  assign n43026 = n42973 ^ n42960;
  assign n43027 = n43025 & ~n43026;
  assign n43028 = n42976 ^ n42958;
  assign n43029 = n43027 & n43028;
  assign n43030 = ~n43020 & ~n43029;
  assign n43031 = n42984 ^ n42956;
  assign n43032 = n43030 & ~n43031;
  assign n43033 = n43019 & ~n43032;
  assign n43034 = n42990 ^ n42952;
  assign n43035 = n43033 & ~n43034;
  assign n43036 = ~n43018 & ~n43035;
  assign n43037 = n42996 ^ n42948;
  assign n43038 = ~n43036 & n43037;
  assign n43039 = ~n43017 & ~n43038;
  assign n43000 = n42999 ^ n42945;
  assign n43001 = ~n42946 & n43000;
  assign n43002 = n43001 ^ n39608;
  assign n42939 = n42938 ^ n42935;
  assign n42940 = ~n42936 & ~n42939;
  assign n42941 = n42940 ^ n42938;
  assign n42286 = n42285 ^ n42266;
  assign n42942 = n42941 ^ n42286;
  assign n42864 = n41094 ^ n40320;
  assign n42865 = n42864 ^ n41843;
  assign n42943 = n42942 ^ n42865;
  assign n42944 = n42943 ^ n39598;
  assign n43016 = n43002 ^ n42944;
  assign n43049 = n43039 ^ n43016;
  assign n43046 = n40985 ^ n32472;
  assign n43047 = n43046 ^ n37107;
  assign n43048 = n43047 ^ n2302;
  assign n43050 = n43049 ^ n43048;
  assign n43131 = n43038 ^ n43017;
  assign n43054 = n43037 ^ n43036;
  assign n43051 = n41050 ^ n32466;
  assign n43052 = n43051 ^ n1108;
  assign n43053 = n43052 ^ n1237;
  assign n43055 = n43054 ^ n43053;
  assign n43056 = n43035 ^ n43018;
  assign n1066 = n1063 ^ n1011;
  assign n1091 = n1090 ^ n1066;
  assign n1098 = n1097 ^ n1091;
  assign n43057 = n43056 ^ n1098;
  assign n43117 = n43034 ^ n43033;
  assign n43059 = n41000 ^ n932;
  assign n43060 = n43059 ^ n37123;
  assign n43061 = n43060 ^ n30699;
  assign n43058 = n43032 ^ n43019;
  assign n43062 = n43061 ^ n43058;
  assign n43106 = n43031 ^ n43030;
  assign n43064 = n41030 ^ n32420;
  assign n43065 = n43064 ^ n37132;
  assign n43066 = n43065 ^ n30688;
  assign n43063 = n43029 ^ n43020;
  assign n43067 = n43066 ^ n43063;
  assign n43071 = n43028 ^ n43027;
  assign n43068 = n41009 ^ n32404;
  assign n43069 = n43068 ^ n37137;
  assign n43070 = n43069 ^ n30717;
  assign n43072 = n43071 ^ n43070;
  assign n43076 = n43026 ^ n43025;
  assign n43073 = n41015 ^ n32387;
  assign n43074 = n43073 ^ n37142;
  assign n43075 = n43074 ^ n662;
  assign n43077 = n43076 ^ n43075;
  assign n43079 = n40654 ^ n32397;
  assign n43080 = n43079 ^ n37148;
  assign n43081 = n43080 ^ n30712;
  assign n43078 = n43024 ^ n43021;
  assign n43082 = n43081 ^ n43078;
  assign n43084 = n40512 ^ n32391;
  assign n43085 = n43084 ^ n37186;
  assign n43086 = n43085 ^ n30706;
  assign n43083 = n43023 ^ n43022;
  assign n43087 = n43086 ^ n43083;
  assign n42829 = n42828 ^ n42827;
  assign n42697 = n42696 ^ n42669;
  assign n42701 = n42700 ^ n42697;
  assign n42703 = n40522 ^ n31871;
  assign n42704 = n42703 ^ n37157;
  assign n42705 = n42704 ^ n30579;
  assign n42702 = n42695 ^ n42694;
  assign n42706 = n42705 ^ n42702;
  assign n42707 = n42693 ^ n42670;
  assign n2255 = n2215 ^ n2158;
  assign n2256 = n2255 ^ n2252;
  assign n2263 = n2262 ^ n2256;
  assign n42708 = n42707 ^ n2263;
  assign n42709 = n42692 ^ n42671;
  assign n2219 = n2200 ^ n2140;
  assign n2238 = n2237 ^ n2219;
  assign n2245 = n2244 ^ n2238;
  assign n42710 = n42709 ^ n2245;
  assign n42800 = n42799 ^ n42711;
  assign n42801 = n42715 & ~n42800;
  assign n42802 = n42801 ^ n42714;
  assign n42803 = n42802 ^ n42709;
  assign n42804 = ~n42710 & n42803;
  assign n42805 = n42804 ^ n2245;
  assign n42806 = n42805 ^ n42707;
  assign n42807 = ~n42708 & n42806;
  assign n42808 = n42807 ^ n2263;
  assign n42809 = n42808 ^ n42702;
  assign n42810 = n42706 & ~n42809;
  assign n42811 = n42810 ^ n42705;
  assign n42812 = n42811 ^ n42697;
  assign n42813 = ~n42701 & n42812;
  assign n42814 = n42813 ^ n42700;
  assign n42830 = n42829 ^ n42814;
  assign n43088 = n42833 ^ n42829;
  assign n43089 = ~n42830 & n43088;
  assign n43090 = n43089 ^ n42833;
  assign n43091 = n43090 ^ n43083;
  assign n43092 = ~n43087 & n43091;
  assign n43093 = n43092 ^ n43086;
  assign n43094 = n43093 ^ n43078;
  assign n43095 = n43082 & ~n43094;
  assign n43096 = n43095 ^ n43081;
  assign n43097 = n43096 ^ n43076;
  assign n43098 = ~n43077 & n43097;
  assign n43099 = n43098 ^ n43075;
  assign n43100 = n43099 ^ n43071;
  assign n43101 = n43072 & ~n43100;
  assign n43102 = n43101 ^ n43070;
  assign n43103 = n43102 ^ n43063;
  assign n43104 = ~n43067 & n43103;
  assign n43105 = n43104 ^ n43066;
  assign n43107 = n43106 ^ n43105;
  assign n43111 = n43110 ^ n43106;
  assign n43112 = ~n43107 & n43111;
  assign n43113 = n43112 ^ n43110;
  assign n43114 = n43113 ^ n43058;
  assign n43115 = ~n43062 & n43114;
  assign n43116 = n43115 ^ n43061;
  assign n43118 = n43117 ^ n43116;
  assign n43119 = n40995 ^ n940;
  assign n43120 = n43119 ^ n37118;
  assign n43121 = n43120 ^ n1089;
  assign n43122 = n43121 ^ n43117;
  assign n43123 = n43118 & ~n43122;
  assign n43124 = n43123 ^ n43121;
  assign n43125 = n43124 ^ n43056;
  assign n43126 = ~n43057 & n43125;
  assign n43127 = n43126 ^ n1098;
  assign n43128 = n43127 ^ n43054;
  assign n43129 = ~n43055 & n43128;
  assign n43130 = n43129 ^ n43053;
  assign n43132 = n43131 ^ n43130;
  assign n1230 = n1229 ^ n1154;
  assign n1246 = n1245 ^ n1230;
  assign n1253 = n1252 ^ n1246;
  assign n43133 = n43131 ^ n1253;
  assign n43134 = n43132 & ~n43133;
  assign n43135 = n43134 ^ n1253;
  assign n43136 = n43135 ^ n43049;
  assign n43137 = n43050 & ~n43136;
  assign n43138 = n43137 ^ n43048;
  assign n43042 = n41064 ^ n32494;
  assign n43043 = n43042 ^ n2303;
  assign n43044 = n43043 ^ n30805;
  assign n43040 = ~n43016 & ~n43039;
  assign n43009 = n42865 ^ n42286;
  assign n43010 = n42942 & ~n43009;
  assign n43011 = n43010 ^ n42865;
  assign n43008 = n42441 ^ n42438;
  assign n43012 = n43011 ^ n43008;
  assign n43006 = n41092 ^ n40314;
  assign n43007 = n43006 ^ n41841;
  assign n43013 = n43012 ^ n43007;
  assign n43014 = n43013 ^ n39596;
  assign n43003 = n43002 ^ n42943;
  assign n43004 = n42944 & ~n43003;
  assign n43005 = n43004 ^ n39598;
  assign n43015 = n43014 ^ n43005;
  assign n43041 = n43040 ^ n43015;
  assign n43045 = n43044 ^ n43041;
  assign n43176 = n43138 ^ n43045;
  assign n43167 = n43132 ^ n1253;
  assign n43168 = n41672 ^ n40752;
  assign n43169 = n43168 ^ n42318;
  assign n43170 = ~n43167 & ~n43169;
  assign n43165 = n41666 ^ n40746;
  assign n43166 = n43165 ^ n42312;
  assign n43171 = n43170 ^ n43166;
  assign n43172 = n43135 ^ n43050;
  assign n43173 = n43172 ^ n43166;
  assign n43174 = ~n43171 & n43173;
  assign n43175 = n43174 ^ n43170;
  assign n43177 = n43176 ^ n43175;
  assign n43178 = n41663 ^ n40740;
  assign n43179 = n43178 ^ n42308;
  assign n43180 = n43179 ^ n43176;
  assign n43181 = ~n43177 & ~n43180;
  assign n43182 = n43181 ^ n43179;
  assign n43162 = n41657 ^ n40738;
  assign n43163 = n43162 ^ n42304;
  assign n43158 = n40981 ^ n32499;
  assign n43159 = n43158 ^ n37102;
  assign n43160 = n43159 ^ n2369;
  assign n43155 = n43015 & n43040;
  assign n43150 = n40763 ^ n40082;
  assign n43151 = n43150 ^ n41831;
  assign n43148 = n42449 ^ n42446;
  assign n43145 = n43008 ^ n43007;
  assign n43146 = n43012 & n43145;
  assign n43147 = n43146 ^ n43007;
  assign n43149 = n43148 ^ n43147;
  assign n43152 = n43151 ^ n43149;
  assign n43153 = n43152 ^ n39428;
  assign n43142 = n43013 ^ n43005;
  assign n43143 = ~n43014 & n43142;
  assign n43144 = n43143 ^ n39596;
  assign n43154 = n43153 ^ n43144;
  assign n43156 = n43155 ^ n43154;
  assign n43139 = n43138 ^ n43041;
  assign n43140 = n43045 & ~n43139;
  assign n43141 = n43140 ^ n43044;
  assign n43157 = n43156 ^ n43141;
  assign n43161 = n43160 ^ n43157;
  assign n43164 = n43163 ^ n43161;
  assign n43351 = n43182 ^ n43164;
  assign n43352 = n43351 ^ n40056;
  assign n43353 = n43179 ^ n43177;
  assign n43354 = n43353 ^ n40058;
  assign n43355 = n43169 ^ n43167;
  assign n43356 = n40070 & n43355;
  assign n43357 = n43356 ^ n40064;
  assign n43358 = n43172 ^ n43171;
  assign n43359 = n43358 ^ n43356;
  assign n43360 = ~n43357 & n43359;
  assign n43361 = n43360 ^ n40064;
  assign n43362 = n43361 ^ n43353;
  assign n43363 = n43354 & ~n43362;
  assign n43364 = n43363 ^ n40058;
  assign n43365 = n43364 ^ n43351;
  assign n43366 = n43352 & ~n43365;
  assign n43367 = n43366 ^ n40056;
  assign n43210 = n41647 ^ n40732;
  assign n43211 = n43210 ^ n42561;
  assign n43206 = ~n43154 & ~n43155;
  assign n43202 = n40976 ^ n32369;
  assign n43203 = n43202 ^ n37252;
  assign n43204 = n43203 ^ n30939;
  assign n43197 = n40753 ^ n40076;
  assign n43198 = n43197 ^ n41829;
  assign n43196 = n42452 ^ n42433;
  assign n43199 = n43198 ^ n43196;
  assign n43193 = n43151 ^ n43148;
  assign n43194 = ~n43149 & ~n43193;
  assign n43195 = n43194 ^ n43151;
  assign n43200 = n43199 ^ n43195;
  assign n43189 = n43152 ^ n43144;
  assign n43190 = ~n43153 & n43189;
  assign n43191 = n43190 ^ n39428;
  assign n43192 = n43191 ^ n39426;
  assign n43201 = n43200 ^ n43192;
  assign n43205 = n43204 ^ n43201;
  assign n43207 = n43206 ^ n43205;
  assign n43186 = n43160 ^ n43156;
  assign n43187 = n43157 & ~n43186;
  assign n43188 = n43187 ^ n43160;
  assign n43208 = n43207 ^ n43188;
  assign n43183 = n43182 ^ n43161;
  assign n43184 = n43164 & ~n43183;
  assign n43185 = n43184 ^ n43163;
  assign n43209 = n43208 ^ n43185;
  assign n43349 = n43211 ^ n43209;
  assign n43350 = n43349 ^ n40050;
  assign n43451 = n43367 ^ n43350;
  assign n43452 = n43364 ^ n40056;
  assign n43453 = n43452 ^ n43351;
  assign n43454 = n43358 ^ n43357;
  assign n43455 = n43361 ^ n43354;
  assign n43456 = ~n43454 & n43455;
  assign n43457 = ~n43453 & ~n43456;
  assign n43458 = n43451 & ~n43457;
  assign n43212 = n43211 ^ n43208;
  assign n43213 = ~n43209 & n43212;
  assign n43214 = n43213 ^ n43211;
  assign n42862 = n42749 ^ n42746;
  assign n42860 = n41641 ^ n40726;
  assign n42861 = n42860 ^ n42302;
  assign n42863 = n42862 ^ n42861;
  assign n43371 = n43214 ^ n42863;
  assign n43368 = n43367 ^ n43349;
  assign n43369 = n43350 & ~n43368;
  assign n43370 = n43369 ^ n40050;
  assign n43372 = n43371 ^ n43370;
  assign n43450 = n43372 ^ n40040;
  assign n43612 = n43458 ^ n43450;
  assign n43577 = n41459 ^ n32687;
  assign n43578 = n43577 ^ n37369;
  assign n43579 = n43578 ^ n31245;
  assign n43576 = n43457 ^ n43451;
  assign n43580 = n43579 ^ n43576;
  assign n43582 = n41463 ^ n32691;
  assign n43583 = n43582 ^ n37373;
  assign n43584 = n43583 ^ n30865;
  assign n43581 = n43456 ^ n43453;
  assign n43585 = n43584 ^ n43581;
  assign n43587 = n41472 ^ n32700;
  assign n43588 = n43587 ^ n37379;
  assign n43589 = n43588 ^ n30874;
  assign n43586 = n43455 ^ n43454;
  assign n43590 = n43589 ^ n43586;
  assign n43596 = n41468 ^ n32696;
  assign n43597 = n43596 ^ n2579;
  assign n43598 = n43597 ^ n30869;
  assign n43591 = n41810 ^ n33369;
  assign n43592 = n43591 ^ n38048;
  assign n43593 = n43592 ^ n2578;
  assign n43594 = n43355 ^ n40070;
  assign n43595 = n43593 & n43594;
  assign n43599 = n43598 ^ n43595;
  assign n43600 = n43595 ^ n43454;
  assign n43601 = n43599 & n43600;
  assign n43602 = n43601 ^ n43598;
  assign n43603 = n43602 ^ n43586;
  assign n43604 = n43590 & ~n43603;
  assign n43605 = n43604 ^ n43589;
  assign n43606 = n43605 ^ n43581;
  assign n43607 = n43585 & ~n43606;
  assign n43608 = n43607 ^ n43584;
  assign n43609 = n43608 ^ n43576;
  assign n43610 = n43580 & ~n43609;
  assign n43611 = n43610 ^ n43579;
  assign n43613 = n43612 ^ n43611;
  assign n43617 = n43616 ^ n43612;
  assign n43618 = n43613 & ~n43617;
  assign n43619 = n43618 ^ n43616;
  assign n43572 = n41449 ^ n32680;
  assign n43573 = n43572 ^ n37359;
  assign n43574 = n43573 ^ n31234;
  assign n43459 = n43450 & ~n43458;
  assign n43373 = n43371 ^ n40040;
  assign n43374 = n43372 & ~n43373;
  assign n43375 = n43374 ^ n40040;
  assign n43215 = n43214 ^ n42862;
  assign n43216 = ~n42863 & n43215;
  assign n43217 = n43216 ^ n42861;
  assign n42857 = n41639 ^ n40720;
  assign n42858 = n42857 ^ n42298;
  assign n42855 = n42753 ^ n42676;
  assign n42856 = n42855 ^ n42750;
  assign n42859 = n42858 ^ n42856;
  assign n43347 = n43217 ^ n42859;
  assign n43348 = n43347 ^ n40038;
  assign n43449 = n43375 ^ n43348;
  assign n43571 = n43459 ^ n43449;
  assign n43575 = n43574 ^ n43571;
  assign n43951 = n43619 ^ n43575;
  assign n43800 = n42850 ^ n41615;
  assign n42838 = n42796 ^ n42720;
  assign n43801 = n43800 ^ n42838;
  assign n43755 = n43616 ^ n43613;
  assign n43802 = n43801 ^ n43755;
  assign n43805 = n42665 ^ n41627;
  assign n42844 = n42785 ^ n42725;
  assign n43806 = n43805 ^ n42844;
  assign n43804 = n43605 ^ n43585;
  assign n43807 = n43806 ^ n43804;
  assign n43932 = n43602 ^ n43590;
  assign n43810 = n42577 ^ n41639;
  assign n42854 = n42774 ^ n42730;
  assign n43811 = n43810 ^ n42854;
  assign n43808 = n43598 ^ n43454;
  assign n43809 = n43808 ^ n43595;
  assign n43812 = n43811 ^ n43809;
  assign n43815 = n43594 ^ n43593;
  assign n43813 = n42292 ^ n41641;
  assign n43243 = n42771 ^ n42768;
  assign n43814 = n43813 ^ n43243;
  assign n43816 = n43815 ^ n43814;
  assign n43832 = n43113 ^ n43062;
  assign n43737 = n43110 ^ n43107;
  assign n43715 = n43102 ^ n43067;
  assign n43439 = n43096 ^ n43077;
  assign n43314 = n43093 ^ n43082;
  assign n43307 = n43090 ^ n43087;
  assign n42834 = n42833 ^ n42830;
  assign n42289 = n42288 ^ n41698;
  assign n42291 = n42290 ^ n42289;
  assign n42835 = n42834 ^ n42291;
  assign n43297 = n42811 ^ n42701;
  assign n43290 = n42808 ^ n42706;
  assign n42841 = n42038 ^ n40659;
  assign n42842 = n42841 ^ n42840;
  assign n42839 = n42793 ^ n42790;
  assign n42843 = n42842 ^ n42839;
  assign n42846 = n41917 ^ n40666;
  assign n42847 = n42846 ^ n42845;
  assign n42848 = n42847 ^ n42844;
  assign n42851 = n41603 ^ n40673;
  assign n42852 = n42851 ^ n42850;
  assign n42849 = n42782 ^ n42779;
  assign n42853 = n42852 ^ n42849;
  assign n43236 = n42763 ^ n42735;
  assign n43229 = n42760 ^ n42740;
  assign n43221 = n42757 ^ n42743;
  assign n43222 = n43221 ^ n42744;
  assign n43218 = n43217 ^ n42856;
  assign n43219 = ~n42859 & n43218;
  assign n43220 = n43219 ^ n42858;
  assign n43223 = n43222 ^ n43220;
  assign n43224 = n41629 ^ n40708;
  assign n43225 = n43224 ^ n42292;
  assign n43226 = n43225 ^ n43222;
  assign n43227 = n43223 & n43226;
  assign n43228 = n43227 ^ n43225;
  assign n43230 = n43229 ^ n43228;
  assign n43231 = n41627 ^ n40706;
  assign n43232 = n43231 ^ n42577;
  assign n43233 = n43232 ^ n43229;
  assign n43234 = ~n43230 & ~n43233;
  assign n43235 = n43234 ^ n43232;
  assign n43237 = n43236 ^ n43235;
  assign n43238 = n41617 ^ n40699;
  assign n43239 = n43238 ^ n42584;
  assign n43240 = n43239 ^ n43236;
  assign n43241 = ~n43237 & n43240;
  assign n43242 = n43241 ^ n43239;
  assign n43244 = n43243 ^ n43242;
  assign n43245 = n41615 ^ n40687;
  assign n43246 = n43245 ^ n42665;
  assign n43247 = n43246 ^ n43243;
  assign n43248 = ~n43244 & ~n43247;
  assign n43249 = n43248 ^ n43246;
  assign n43250 = n43249 ^ n42854;
  assign n43251 = n41609 ^ n40680;
  assign n43252 = n43251 ^ n42821;
  assign n43253 = n43252 ^ n42854;
  assign n43254 = ~n43250 & n43253;
  assign n43255 = n43254 ^ n43252;
  assign n43256 = n43255 ^ n42849;
  assign n43257 = n42853 & ~n43256;
  assign n43258 = n43257 ^ n42852;
  assign n43259 = n43258 ^ n42844;
  assign n43260 = n42848 & ~n43259;
  assign n43261 = n43260 ^ n42847;
  assign n43262 = n43261 ^ n42839;
  assign n43263 = ~n42843 & n43262;
  assign n43264 = n43263 ^ n42842;
  assign n43265 = n43264 ^ n42838;
  assign n43266 = n42092 ^ n40656;
  assign n43267 = n43266 ^ n42900;
  assign n43268 = n43267 ^ n42838;
  assign n43269 = n43265 & n43268;
  assign n43270 = n43269 ^ n43267;
  assign n43272 = n43271 ^ n43270;
  assign n43273 = n42280 ^ n41189;
  assign n43274 = n43273 ^ n42907;
  assign n43275 = n43274 ^ n43271;
  assign n43276 = n43272 & ~n43275;
  assign n43277 = n43276 ^ n43274;
  assign n42837 = n42802 ^ n42710;
  assign n43278 = n43277 ^ n42837;
  assign n43279 = n42344 ^ n41332;
  assign n43280 = n43279 ^ n42875;
  assign n43281 = n43280 ^ n42837;
  assign n43282 = ~n43278 & n43281;
  assign n43283 = n43282 ^ n43280;
  assign n42836 = n42805 ^ n42708;
  assign n43284 = n43283 ^ n42836;
  assign n43285 = n42338 ^ n41582;
  assign n43286 = n43285 ^ n42874;
  assign n43287 = n43286 ^ n42836;
  assign n43288 = ~n43284 & n43287;
  assign n43289 = n43288 ^ n43286;
  assign n43291 = n43290 ^ n43289;
  assign n43292 = n42332 ^ n41710;
  assign n43293 = n43292 ^ n42870;
  assign n43294 = n43293 ^ n43290;
  assign n43295 = n43291 & ~n43294;
  assign n43296 = n43295 ^ n43293;
  assign n43298 = n43297 ^ n43296;
  assign n43299 = n42326 ^ n41704;
  assign n43300 = n43299 ^ n42866;
  assign n43301 = n43300 ^ n43297;
  assign n43302 = ~n43298 & n43301;
  assign n43303 = n43302 ^ n43300;
  assign n43304 = n43303 ^ n42834;
  assign n43305 = ~n42835 & n43304;
  assign n43306 = n43305 ^ n42291;
  assign n43308 = n43307 ^ n43306;
  assign n43309 = n42404 ^ n41728;
  assign n43310 = n43309 ^ n42935;
  assign n43311 = n43310 ^ n43307;
  assign n43312 = ~n43308 & ~n43311;
  assign n43313 = n43312 ^ n43310;
  assign n43315 = n43314 ^ n43313;
  assign n41598 = n41597 ^ n41596;
  assign n42287 = n42286 ^ n41598;
  assign n43436 = n43314 ^ n42287;
  assign n43437 = ~n43315 & ~n43436;
  assign n43438 = n43437 ^ n42287;
  assign n43440 = n43439 ^ n43438;
  assign n43434 = n42537 ^ n41824;
  assign n43435 = n43434 ^ n43008;
  assign n43499 = n43439 ^ n43435;
  assign n43500 = ~n43440 & n43499;
  assign n43501 = n43500 ^ n43435;
  assign n43498 = n43099 ^ n43072;
  assign n43502 = n43501 ^ n43498;
  assign n43496 = n41853 ^ n41112;
  assign n43497 = n43496 ^ n43148;
  assign n43712 = n43498 ^ n43497;
  assign n43713 = n43502 & ~n43712;
  assign n43714 = n43713 ^ n43497;
  assign n43716 = n43715 ^ n43714;
  assign n43710 = n41843 ^ n41110;
  assign n43711 = n43710 ^ n43196;
  assign n43734 = n43715 ^ n43711;
  assign n43735 = ~n43716 & ~n43734;
  assign n43736 = n43735 ^ n43711;
  assign n43738 = n43737 ^ n43736;
  assign n43732 = n41841 ^ n41104;
  assign n43733 = n43732 ^ n42501;
  assign n43829 = n43737 ^ n43733;
  assign n43830 = ~n43738 & n43829;
  assign n43831 = n43830 ^ n43733;
  assign n43833 = n43832 ^ n43831;
  assign n43827 = n41831 ^ n41094;
  assign n43828 = n43827 ^ n42504;
  assign n43834 = n43833 ^ n43828;
  assign n43835 = n43834 ^ n40320;
  assign n43739 = n43738 ^ n43733;
  assign n43740 = n43739 ^ n40326;
  assign n43717 = n43716 ^ n43711;
  assign n43718 = n43717 ^ n40332;
  assign n43503 = n43502 ^ n43497;
  assign n43504 = n43503 ^ n40338;
  assign n43441 = n43440 ^ n43435;
  assign n43442 = n43441 ^ n41087;
  assign n43316 = n43315 ^ n42287;
  assign n43317 = n43316 ^ n40968;
  assign n43318 = n43310 ^ n43308;
  assign n43319 = n43318 ^ n40952;
  assign n43320 = n43303 ^ n42291;
  assign n43321 = n43320 ^ n42834;
  assign n43322 = n43321 ^ n40914;
  assign n43323 = n43300 ^ n43298;
  assign n43324 = n43323 ^ n40024;
  assign n43325 = n43293 ^ n43291;
  assign n43326 = n43325 ^ n40661;
  assign n43327 = n43286 ^ n43284;
  assign n43328 = n43327 ^ n40668;
  assign n43329 = n43280 ^ n43278;
  assign n43330 = n43329 ^ n40675;
  assign n43331 = n43274 ^ n43272;
  assign n43332 = n43331 ^ n40682;
  assign n43333 = n43267 ^ n43265;
  assign n43334 = n43333 ^ n40689;
  assign n43335 = n43261 ^ n42843;
  assign n43336 = n43335 ^ n40695;
  assign n43337 = n43258 ^ n42848;
  assign n43338 = n43337 ^ n40702;
  assign n43339 = n43255 ^ n42853;
  assign n43340 = n43339 ^ n40710;
  assign n43393 = n43252 ^ n43250;
  assign n43341 = n43246 ^ n43244;
  assign n43342 = n43341 ^ n40646;
  assign n43385 = n43239 ^ n43237;
  assign n43343 = n43232 ^ n43230;
  assign n43344 = n43343 ^ n40386;
  assign n43345 = n43225 ^ n43223;
  assign n43346 = n43345 ^ n40032;
  assign n43376 = n43375 ^ n43347;
  assign n43377 = n43348 & n43376;
  assign n43378 = n43377 ^ n40038;
  assign n43379 = n43378 ^ n43345;
  assign n43380 = ~n43346 & n43379;
  assign n43381 = n43380 ^ n40032;
  assign n43382 = n43381 ^ n43343;
  assign n43383 = n43344 & n43382;
  assign n43384 = n43383 ^ n40386;
  assign n43386 = n43385 ^ n43384;
  assign n43387 = n43385 ^ n40476;
  assign n43388 = ~n43386 & ~n43387;
  assign n43389 = n43388 ^ n40476;
  assign n43390 = n43389 ^ n43341;
  assign n43391 = n43342 & ~n43390;
  assign n43392 = n43391 ^ n40646;
  assign n43394 = n43393 ^ n43392;
  assign n43395 = n43393 ^ n40716;
  assign n43396 = ~n43394 & ~n43395;
  assign n43397 = n43396 ^ n40716;
  assign n43398 = n43397 ^ n43339;
  assign n43399 = ~n43340 & n43398;
  assign n43400 = n43399 ^ n40710;
  assign n43401 = n43400 ^ n43337;
  assign n43402 = n43338 & n43401;
  assign n43403 = n43402 ^ n40702;
  assign n43404 = n43403 ^ n43335;
  assign n43405 = n43336 & n43404;
  assign n43406 = n43405 ^ n40695;
  assign n43407 = n43406 ^ n43333;
  assign n43408 = n43334 & n43407;
  assign n43409 = n43408 ^ n40689;
  assign n43410 = n43409 ^ n43331;
  assign n43411 = ~n43332 & ~n43410;
  assign n43412 = n43411 ^ n40682;
  assign n43413 = n43412 ^ n43329;
  assign n43414 = n43330 & ~n43413;
  assign n43415 = n43414 ^ n40675;
  assign n43416 = n43415 ^ n43327;
  assign n43417 = ~n43328 & ~n43416;
  assign n43418 = n43417 ^ n40668;
  assign n43419 = n43418 ^ n43325;
  assign n43420 = ~n43326 & ~n43419;
  assign n43421 = n43420 ^ n40661;
  assign n43422 = n43421 ^ n43323;
  assign n43423 = ~n43324 & ~n43422;
  assign n43424 = n43423 ^ n40024;
  assign n43425 = n43424 ^ n43321;
  assign n43426 = n43322 & ~n43425;
  assign n43427 = n43426 ^ n40914;
  assign n43428 = n43427 ^ n43318;
  assign n43429 = ~n43319 & ~n43428;
  assign n43430 = n43429 ^ n40952;
  assign n43431 = n43430 ^ n43316;
  assign n43432 = n43317 & ~n43431;
  assign n43433 = n43432 ^ n40968;
  assign n43493 = n43441 ^ n43433;
  assign n43494 = n43442 & ~n43493;
  assign n43495 = n43494 ^ n41087;
  assign n43707 = n43503 ^ n43495;
  assign n43708 = ~n43504 & n43707;
  assign n43709 = n43708 ^ n40338;
  assign n43729 = n43717 ^ n43709;
  assign n43730 = n43718 & n43729;
  assign n43731 = n43730 ^ n40332;
  assign n43824 = n43739 ^ n43731;
  assign n43825 = n43740 & ~n43824;
  assign n43826 = n43825 ^ n40326;
  assign n43836 = n43835 ^ n43826;
  assign n43741 = n43740 ^ n43731;
  assign n43719 = n43718 ^ n43709;
  assign n43443 = n43442 ^ n43433;
  assign n43444 = n43415 ^ n43328;
  assign n43445 = n43409 ^ n43332;
  assign n43446 = n43403 ^ n43336;
  assign n43447 = n43389 ^ n43342;
  assign n43448 = n43381 ^ n43344;
  assign n43460 = n43449 & ~n43459;
  assign n43461 = n43378 ^ n43346;
  assign n43462 = n43460 & n43461;
  assign n43463 = ~n43448 & n43462;
  assign n43464 = n43386 ^ n40476;
  assign n43465 = ~n43463 & n43464;
  assign n43466 = n43447 & n43465;
  assign n43467 = n43394 ^ n40716;
  assign n43468 = n43466 & ~n43467;
  assign n43469 = n43397 ^ n43340;
  assign n43470 = n43468 & n43469;
  assign n43471 = n43400 ^ n43338;
  assign n43472 = n43470 & ~n43471;
  assign n43473 = ~n43446 & ~n43472;
  assign n43474 = n43406 ^ n43334;
  assign n43475 = n43473 & n43474;
  assign n43476 = ~n43445 & ~n43475;
  assign n43477 = n43412 ^ n43330;
  assign n43478 = ~n43476 & n43477;
  assign n43479 = n43444 & ~n43478;
  assign n43480 = n43418 ^ n43326;
  assign n43481 = n43479 & ~n43480;
  assign n43482 = n43421 ^ n43324;
  assign n43483 = n43481 & n43482;
  assign n43484 = n43424 ^ n43322;
  assign n43485 = ~n43483 & ~n43484;
  assign n43486 = n43427 ^ n40952;
  assign n43487 = n43486 ^ n43318;
  assign n43488 = n43485 & n43487;
  assign n43489 = n43430 ^ n40968;
  assign n43490 = n43489 ^ n43316;
  assign n43491 = ~n43488 & ~n43490;
  assign n43492 = ~n43443 & n43491;
  assign n43505 = n43504 ^ n43495;
  assign n43720 = ~n43492 & ~n43505;
  assign n43742 = ~n43719 & ~n43720;
  assign n43837 = ~n43741 & ~n43742;
  assign n43850 = n43836 & ~n43837;
  assign n43856 = n43832 ^ n43828;
  assign n43857 = n43833 & ~n43856;
  assign n43858 = n43857 ^ n43828;
  assign n43767 = n43121 ^ n43118;
  assign n43859 = n43858 ^ n43767;
  assign n43854 = n41829 ^ n41092;
  assign n43855 = n43854 ^ n42508;
  assign n43860 = n43859 ^ n43855;
  assign n43861 = n43860 ^ n40314;
  assign n43851 = n43834 ^ n43826;
  assign n43852 = n43835 & n43851;
  assign n43853 = n43852 ^ n40320;
  assign n43862 = n43861 ^ n43853;
  assign n43878 = n43850 & n43862;
  assign n43886 = n41684 ^ n40763;
  assign n43887 = n43886 ^ n42495;
  assign n43882 = n43855 ^ n43767;
  assign n43883 = n43859 & n43882;
  assign n43884 = n43883 ^ n43855;
  assign n43763 = n43124 ^ n43057;
  assign n43885 = n43884 ^ n43763;
  assign n43888 = n43887 ^ n43885;
  assign n43879 = n43860 ^ n43853;
  assign n43880 = ~n43861 & n43879;
  assign n43881 = n43880 ^ n40314;
  assign n43889 = n43888 ^ n43881;
  assign n43890 = n43889 ^ n40082;
  assign n43916 = ~n43878 & ~n43890;
  assign n43913 = n43127 ^ n43055;
  assign n43910 = n41678 ^ n40753;
  assign n43911 = n43910 ^ n42542;
  assign n43907 = n43887 ^ n43763;
  assign n43908 = ~n43885 & n43907;
  assign n43909 = n43908 ^ n43887;
  assign n43912 = n43911 ^ n43909;
  assign n43914 = n43913 ^ n43912;
  assign n43903 = n43888 ^ n40082;
  assign n43904 = ~n43889 & ~n43903;
  assign n43905 = n43904 ^ n40082;
  assign n43906 = n43905 ^ n40076;
  assign n43915 = n43914 ^ n43906;
  assign n43917 = n43916 ^ n43915;
  assign n2433 = n2432 ^ n2405;
  assign n2461 = n2460 ^ n2433;
  assign n2468 = n2467 ^ n2461;
  assign n43918 = n43917 ^ n2468;
  assign n43891 = n43890 ^ n43878;
  assign n43875 = n41779 ^ n33189;
  assign n43876 = n43875 ^ n37874;
  assign n43877 = n43876 ^ n2459;
  assign n43892 = n43891 ^ n43877;
  assign n43863 = n43862 ^ n43850;
  assign n43847 = n41784 ^ n2337;
  assign n43848 = n43847 ^ n37878;
  assign n43849 = n43848 ^ n31594;
  assign n43864 = n43863 ^ n43849;
  assign n43838 = n43837 ^ n43836;
  assign n1400 = n1360 ^ n1300;
  assign n1401 = n1400 ^ n1397;
  assign n1408 = n1407 ^ n1401;
  assign n43839 = n43838 ^ n1408;
  assign n43743 = n43742 ^ n43741;
  assign n43721 = n43720 ^ n43719;
  assign n43507 = n41384 ^ n1172;
  assign n43508 = n43507 ^ n37888;
  assign n43509 = n43508 ^ n31605;
  assign n43506 = n43505 ^ n43492;
  assign n43510 = n43509 ^ n43506;
  assign n43514 = n43491 ^ n43443;
  assign n43515 = n43514 ^ n43513;
  assign n43517 = n41394 ^ n33270;
  assign n43518 = n43517 ^ n37898;
  assign n43519 = n43518 ^ n833;
  assign n43516 = n43490 ^ n43488;
  assign n43520 = n43519 ^ n43516;
  assign n43690 = n43487 ^ n43485;
  assign n43522 = n41404 ^ n33280;
  assign n43523 = n43522 ^ n37905;
  assign n43524 = n43523 ^ n751;
  assign n43521 = n43484 ^ n43483;
  assign n43525 = n43524 ^ n43521;
  assign n43527 = n41555 ^ n680;
  assign n43528 = n43527 ^ n37910;
  assign n43529 = n43528 ^ n31624;
  assign n43526 = n43482 ^ n43481;
  assign n43530 = n43529 ^ n43526;
  assign n43534 = n43480 ^ n43479;
  assign n43531 = n41408 ^ n33250;
  assign n43532 = n43531 ^ n37915;
  assign n43533 = n43532 ^ n31629;
  assign n43535 = n43534 ^ n43533;
  assign n43536 = n43478 ^ n43444;
  assign n43540 = n43539 ^ n43536;
  assign n43670 = n43477 ^ n43476;
  assign n43662 = n43475 ^ n43445;
  assign n43541 = n43474 ^ n43473;
  assign n43545 = n43544 ^ n43541;
  assign n43547 = n41424 ^ n33209;
  assign n43548 = n43547 ^ n37935;
  assign n43549 = n43548 ^ n31207;
  assign n43546 = n43472 ^ n43446;
  assign n43550 = n43549 ^ n43546;
  assign n43552 = n41519 ^ n33215;
  assign n43553 = n43552 ^ n37978;
  assign n43554 = n43553 ^ n31212;
  assign n43551 = n43471 ^ n43470;
  assign n43555 = n43554 ^ n43551;
  assign n43556 = n43469 ^ n43468;
  assign n43560 = n43559 ^ n43556;
  assign n43562 = n41429 ^ n33225;
  assign n43563 = n43562 ^ n1931;
  assign n43564 = n43563 ^ n31219;
  assign n43561 = n43467 ^ n43466;
  assign n43565 = n43564 ^ n43561;
  assign n43639 = n43465 ^ n43447;
  assign n43634 = n43464 ^ n43463;
  assign n43569 = n43462 ^ n43448;
  assign n43566 = n37949 ^ n32668;
  assign n43567 = n43566 ^ n41438;
  assign n43568 = n43567 ^ n1795;
  assign n43570 = n43569 ^ n43568;
  assign n43623 = n43461 ^ n43460;
  assign n43620 = n43619 ^ n43571;
  assign n43621 = n43575 & ~n43620;
  assign n43622 = n43621 ^ n43574;
  assign n43624 = n43623 ^ n43622;
  assign n43628 = n43627 ^ n43622;
  assign n43629 = n43624 & n43628;
  assign n43630 = n43629 ^ n43627;
  assign n43631 = n43630 ^ n43569;
  assign n43632 = n43570 & ~n43631;
  assign n43633 = n43632 ^ n43568;
  assign n43635 = n43634 ^ n43633;
  assign n1776 = n1775 ^ n1745;
  assign n1804 = n1803 ^ n1776;
  assign n1811 = n1810 ^ n1804;
  assign n43636 = n43634 ^ n1811;
  assign n43637 = n43635 & ~n43636;
  assign n43638 = n43637 ^ n1811;
  assign n43640 = n43639 ^ n43638;
  assign n43641 = n41433 ^ n32747;
  assign n43642 = n43641 ^ n37944;
  assign n43643 = n43642 ^ n1923;
  assign n43644 = n43643 ^ n43639;
  assign n43645 = ~n43640 & n43644;
  assign n43646 = n43645 ^ n43643;
  assign n43647 = n43646 ^ n43561;
  assign n43648 = ~n43565 & n43647;
  assign n43649 = n43648 ^ n43564;
  assign n43650 = n43649 ^ n43556;
  assign n43651 = n43560 & ~n43650;
  assign n43652 = n43651 ^ n43559;
  assign n43653 = n43652 ^ n43551;
  assign n43654 = ~n43555 & n43653;
  assign n43655 = n43654 ^ n43554;
  assign n43656 = n43655 ^ n43546;
  assign n43657 = ~n43550 & n43656;
  assign n43658 = n43657 ^ n43549;
  assign n43659 = n43658 ^ n43541;
  assign n43660 = ~n43545 & n43659;
  assign n43661 = n43660 ^ n43544;
  assign n43663 = n43662 ^ n43661;
  assign n43664 = n41418 ^ n33200;
  assign n43665 = n43664 ^ n37929;
  assign n43666 = n43665 ^ n31197;
  assign n43667 = n43666 ^ n43662;
  assign n43668 = ~n43663 & n43667;
  assign n43669 = n43668 ^ n43666;
  assign n43671 = n43670 ^ n43669;
  assign n43672 = n41541 ^ n33260;
  assign n43673 = n43672 ^ n37925;
  assign n43674 = n43673 ^ n31192;
  assign n43675 = n43674 ^ n43670;
  assign n43676 = ~n43671 & n43675;
  assign n43677 = n43676 ^ n43674;
  assign n43678 = n43677 ^ n43536;
  assign n43679 = ~n43540 & n43678;
  assign n43680 = n43679 ^ n43539;
  assign n43681 = n43680 ^ n43534;
  assign n43682 = ~n43535 & n43681;
  assign n43683 = n43682 ^ n43533;
  assign n43684 = n43683 ^ n43526;
  assign n43685 = n43530 & ~n43684;
  assign n43686 = n43685 ^ n43529;
  assign n43687 = n43686 ^ n43521;
  assign n43688 = ~n43525 & n43687;
  assign n43689 = n43688 ^ n43524;
  assign n43691 = n43690 ^ n43689;
  assign n43692 = n41398 ^ n33275;
  assign n43693 = n43692 ^ n752;
  assign n43694 = n43693 ^ n31617;
  assign n43695 = n43694 ^ n43690;
  assign n43696 = n43691 & ~n43695;
  assign n43697 = n43696 ^ n43694;
  assign n43698 = n43697 ^ n43516;
  assign n43699 = n43520 & ~n43698;
  assign n43700 = n43699 ^ n43519;
  assign n43701 = n43700 ^ n43514;
  assign n43702 = ~n43515 & n43701;
  assign n43703 = n43702 ^ n43513;
  assign n43704 = n43703 ^ n43506;
  assign n43705 = ~n43510 & n43704;
  assign n43706 = n43705 ^ n43509;
  assign n43722 = n43721 ^ n43706;
  assign n43726 = n43725 ^ n43721;
  assign n43727 = ~n43722 & n43726;
  assign n43728 = n43727 ^ n43725;
  assign n43744 = n43743 ^ n43728;
  assign n1364 = n1345 ^ n1282;
  assign n1383 = n1382 ^ n1364;
  assign n1390 = n1389 ^ n1383;
  assign n43821 = n43743 ^ n1390;
  assign n43822 = n43744 & ~n43821;
  assign n43823 = n43822 ^ n1390;
  assign n43844 = n43838 ^ n43823;
  assign n43845 = ~n43839 & n43844;
  assign n43846 = n43845 ^ n1408;
  assign n43872 = n43863 ^ n43846;
  assign n43873 = n43864 & ~n43872;
  assign n43874 = n43873 ^ n43849;
  assign n43900 = n43891 ^ n43874;
  assign n43901 = ~n43892 & n43900;
  assign n43902 = n43901 ^ n43877;
  assign n43919 = n43918 ^ n43902;
  assign n43893 = n43892 ^ n43874;
  assign n43865 = n43864 ^ n43846;
  assign n43745 = n43744 ^ n1390;
  assign n43746 = n42308 ^ n41672;
  assign n43747 = n43746 ^ n42862;
  assign n43819 = ~n43745 & ~n43747;
  assign n43817 = n42304 ^ n41666;
  assign n43818 = n43817 ^ n42856;
  assign n43820 = n43819 ^ n43818;
  assign n43840 = n43839 ^ n43823;
  assign n43841 = n43840 ^ n43818;
  assign n43842 = ~n43820 & ~n43841;
  assign n43843 = n43842 ^ n43819;
  assign n43866 = n43865 ^ n43843;
  assign n43867 = n42561 ^ n41663;
  assign n43868 = n43867 ^ n43222;
  assign n43869 = n43868 ^ n43865;
  assign n43870 = ~n43866 & n43869;
  assign n43871 = n43870 ^ n43868;
  assign n43894 = n43893 ^ n43871;
  assign n43895 = n42302 ^ n41657;
  assign n43896 = n43895 ^ n43229;
  assign n43897 = n43896 ^ n43893;
  assign n43898 = n43894 & ~n43897;
  assign n43899 = n43898 ^ n43896;
  assign n43920 = n43919 ^ n43899;
  assign n43921 = n42298 ^ n41647;
  assign n43922 = n43921 ^ n43236;
  assign n43923 = n43922 ^ n43919;
  assign n43924 = n43920 & ~n43923;
  assign n43925 = n43924 ^ n43922;
  assign n43926 = n43925 ^ n43815;
  assign n43927 = n43816 & ~n43926;
  assign n43928 = n43927 ^ n43814;
  assign n43929 = n43928 ^ n43809;
  assign n43930 = n43812 & n43929;
  assign n43931 = n43930 ^ n43811;
  assign n43933 = n43932 ^ n43931;
  assign n43934 = n42584 ^ n41629;
  assign n43935 = n43934 ^ n42849;
  assign n43936 = n43935 ^ n43932;
  assign n43937 = n43933 & n43936;
  assign n43938 = n43937 ^ n43935;
  assign n43939 = n43938 ^ n43804;
  assign n43940 = n43807 & ~n43939;
  assign n43941 = n43940 ^ n43806;
  assign n43803 = n43608 ^ n43580;
  assign n43942 = n43941 ^ n43803;
  assign n43943 = n42821 ^ n41617;
  assign n43944 = n43943 ^ n42839;
  assign n43945 = n43944 ^ n43803;
  assign n43946 = ~n43942 & n43945;
  assign n43947 = n43946 ^ n43944;
  assign n43948 = n43947 ^ n43755;
  assign n43949 = n43802 & n43948;
  assign n43950 = n43949 ^ n43801;
  assign n43952 = n43951 ^ n43950;
  assign n44067 = n43954 ^ n43952;
  assign n44068 = n44067 ^ n40680;
  assign n44069 = n43947 ^ n43802;
  assign n44070 = n44069 ^ n40687;
  assign n44071 = n43944 ^ n43942;
  assign n44072 = n44071 ^ n40699;
  assign n44073 = n43938 ^ n43807;
  assign n44074 = n44073 ^ n40706;
  assign n44107 = n43935 ^ n43933;
  assign n44075 = n43928 ^ n43812;
  assign n44076 = n44075 ^ n40720;
  assign n44077 = n43925 ^ n43814;
  assign n44078 = n44077 ^ n43815;
  assign n44079 = n44078 ^ n40726;
  assign n44080 = n43922 ^ n43920;
  assign n44081 = n44080 ^ n40732;
  assign n44082 = n43896 ^ n43894;
  assign n44083 = n44082 ^ n40738;
  assign n44084 = n43868 ^ n43866;
  assign n44085 = n44084 ^ n40740;
  assign n43748 = n43747 ^ n43745;
  assign n44086 = ~n40752 & n43748;
  assign n44087 = n44086 ^ n40746;
  assign n44088 = n43840 ^ n43820;
  assign n44089 = n44088 ^ n44086;
  assign n44090 = ~n44087 & ~n44089;
  assign n44091 = n44090 ^ n40746;
  assign n44092 = n44091 ^ n44084;
  assign n44093 = ~n44085 & n44092;
  assign n44094 = n44093 ^ n40740;
  assign n44095 = n44094 ^ n44082;
  assign n44096 = n44083 & ~n44095;
  assign n44097 = n44096 ^ n40738;
  assign n44098 = n44097 ^ n44080;
  assign n44099 = n44081 & ~n44098;
  assign n44100 = n44099 ^ n40732;
  assign n44101 = n44100 ^ n44078;
  assign n44102 = n44079 & n44101;
  assign n44103 = n44102 ^ n40726;
  assign n44104 = n44103 ^ n44075;
  assign n44105 = ~n44076 & ~n44104;
  assign n44106 = n44105 ^ n40720;
  assign n44108 = n44107 ^ n44106;
  assign n44109 = n44107 ^ n40708;
  assign n44110 = ~n44108 & n44109;
  assign n44111 = n44110 ^ n40708;
  assign n44112 = n44111 ^ n44073;
  assign n44113 = n44074 & n44112;
  assign n44114 = n44113 ^ n40706;
  assign n44115 = n44114 ^ n44071;
  assign n44116 = n44072 & ~n44115;
  assign n44117 = n44116 ^ n40699;
  assign n44118 = n44117 ^ n44069;
  assign n44119 = ~n44070 & ~n44118;
  assign n44120 = n44119 ^ n40687;
  assign n44121 = n44120 ^ n44067;
  assign n44122 = n44068 & ~n44121;
  assign n44123 = n44122 ^ n40680;
  assign n43955 = n43954 ^ n43951;
  assign n43956 = n43952 & n43955;
  assign n43957 = n43956 ^ n43954;
  assign n43797 = n42840 ^ n41603;
  assign n43798 = n43797 ^ n42837;
  assign n43796 = n43627 ^ n43624;
  assign n43799 = n43798 ^ n43796;
  assign n44065 = n43957 ^ n43799;
  assign n44066 = n44065 ^ n40673;
  assign n44217 = n44123 ^ n44066;
  assign n44196 = n44111 ^ n44074;
  assign n44197 = n44108 ^ n40708;
  assign n44198 = n44100 ^ n44079;
  assign n44199 = n44094 ^ n44083;
  assign n44200 = n44091 ^ n44085;
  assign n44201 = n44088 ^ n44087;
  assign n44202 = ~n44200 & n44201;
  assign n44203 = ~n44199 & ~n44202;
  assign n44204 = n44097 ^ n44081;
  assign n44205 = ~n44203 & n44204;
  assign n44206 = ~n44198 & ~n44205;
  assign n44207 = n44103 ^ n44076;
  assign n44208 = ~n44206 & n44207;
  assign n44209 = n44197 & n44208;
  assign n44210 = n44196 & n44209;
  assign n44211 = n44114 ^ n44072;
  assign n44212 = ~n44210 & n44211;
  assign n44213 = n44117 ^ n44070;
  assign n44214 = n44212 & ~n44213;
  assign n44215 = n44120 ^ n44068;
  assign n44216 = n44214 & ~n44215;
  assign n44310 = n44217 ^ n44216;
  assign n44314 = n44313 ^ n44310;
  assign n44315 = n44215 ^ n44214;
  assign n2023 = n2013 ^ n1965;
  assign n2048 = n2047 ^ n2023;
  assign n2055 = n2054 ^ n2048;
  assign n44316 = n44315 ^ n2055;
  assign n44318 = n42140 ^ n1891;
  assign n44319 = n44318 ^ n38244;
  assign n44320 = n44319 ^ n2039;
  assign n44317 = n44213 ^ n44212;
  assign n44321 = n44320 ^ n44317;
  assign n44386 = n44211 ^ n44210;
  assign n44378 = n44209 ^ n44196;
  assign n44370 = n44208 ^ n44197;
  assign n44323 = n42156 ^ n33673;
  assign n44324 = n44323 ^ n38259;
  assign n44325 = n44324 ^ n31898;
  assign n44322 = n44207 ^ n44206;
  assign n44326 = n44325 ^ n44322;
  assign n44359 = n44205 ^ n44198;
  assign n44328 = n42184 ^ n33683;
  assign n44329 = n44328 ^ n38290;
  assign n44330 = n44329 ^ n31905;
  assign n44327 = n44204 ^ n44203;
  assign n44331 = n44330 ^ n44327;
  assign n44333 = n42165 ^ n33687;
  assign n44334 = n44333 ^ n38268;
  assign n44335 = n44334 ^ n31910;
  assign n44332 = n44202 ^ n44199;
  assign n44336 = n44335 ^ n44332;
  assign n44338 = n42171 ^ n33696;
  assign n44339 = n44338 ^ n38277;
  assign n44340 = n44339 ^ n31919;
  assign n44337 = n44201 ^ n44200;
  assign n44341 = n44340 ^ n44337;
  assign n44343 = n33691 ^ n2610;
  assign n44344 = n44343 ^ n38272;
  assign n44345 = n44344 ^ n31914;
  assign n43749 = n43748 ^ n40752;
  assign n43750 = n42523 ^ n2542;
  assign n43751 = n43750 ^ n38827;
  assign n43752 = n43751 ^ n32538;
  assign n44342 = ~n43749 & n43752;
  assign n44346 = n44345 ^ n44342;
  assign n44347 = n44342 ^ n44201;
  assign n44348 = n44346 & ~n44347;
  assign n44349 = n44348 ^ n44345;
  assign n44350 = n44349 ^ n44337;
  assign n44351 = n44341 & ~n44350;
  assign n44352 = n44351 ^ n44340;
  assign n44353 = n44352 ^ n44332;
  assign n44354 = n44336 & ~n44353;
  assign n44355 = n44354 ^ n44335;
  assign n44356 = n44355 ^ n44327;
  assign n44357 = n44331 & ~n44356;
  assign n44358 = n44357 ^ n44330;
  assign n44360 = n44359 ^ n44358;
  assign n44361 = n42161 ^ n33678;
  assign n44362 = n44361 ^ n38263;
  assign n44363 = n44362 ^ n1565;
  assign n44364 = n44363 ^ n44359;
  assign n44365 = ~n44360 & n44364;
  assign n44366 = n44365 ^ n44363;
  assign n44367 = n44366 ^ n44322;
  assign n44368 = n44326 & ~n44367;
  assign n44369 = n44368 ^ n44325;
  assign n44371 = n44370 ^ n44369;
  assign n44375 = n44374 ^ n44370;
  assign n44376 = n44371 & ~n44375;
  assign n44377 = n44376 ^ n44374;
  assign n44379 = n44378 ^ n44377;
  assign n44383 = n44382 ^ n44378;
  assign n44384 = n44379 & ~n44383;
  assign n44385 = n44384 ^ n44382;
  assign n44387 = n44386 ^ n44385;
  assign n44388 = n42204 ^ n1873;
  assign n44389 = n44388 ^ n38310;
  assign n44390 = n44389 ^ n31884;
  assign n44391 = n44390 ^ n44386;
  assign n44392 = n44387 & ~n44391;
  assign n44393 = n44392 ^ n44390;
  assign n44394 = n44393 ^ n44317;
  assign n44395 = ~n44321 & n44394;
  assign n44396 = n44395 ^ n44320;
  assign n44397 = n44396 ^ n44315;
  assign n44398 = ~n44316 & n44397;
  assign n44399 = n44398 ^ n2055;
  assign n44400 = n44399 ^ n44310;
  assign n44401 = ~n44314 & n44400;
  assign n44402 = n44401 ^ n44313;
  assign n43958 = n43957 ^ n43796;
  assign n43959 = ~n43799 & n43958;
  assign n43960 = n43959 ^ n43798;
  assign n43793 = n42900 ^ n41917;
  assign n43794 = n43793 ^ n42836;
  assign n43792 = n43630 ^ n43570;
  assign n43795 = n43794 ^ n43792;
  assign n44128 = n43960 ^ n43795;
  assign n44219 = n44128 ^ n40666;
  assign n44124 = n44123 ^ n44065;
  assign n44125 = n44066 & ~n44124;
  assign n44126 = n44125 ^ n40673;
  assign n44220 = n44219 ^ n44126;
  assign n44218 = n44216 & ~n44217;
  assign n44308 = n44220 ^ n44218;
  assign n2193 = n2192 ^ n2111;
  assign n2209 = n2208 ^ n2193;
  assign n2216 = n2215 ^ n2209;
  assign n44309 = n44308 ^ n2216;
  assign n44762 = n44402 ^ n44309;
  assign n43979 = n43652 ^ n43555;
  assign n45707 = n44762 ^ n43979;
  assign n44741 = n42719 ^ n2132;
  assign n44742 = n44741 ^ n39188;
  assign n44743 = n44742 ^ n33225;
  assign n44544 = n42844 ^ n42577;
  assign n44545 = n44544 ^ n43951;
  assign n44542 = n44345 ^ n44201;
  assign n44543 = n44542 ^ n44342;
  assign n44546 = n44545 ^ n44543;
  assign n43754 = n42849 ^ n42292;
  assign n43756 = n43755 ^ n43754;
  assign n43753 = n43752 ^ n43749;
  assign n43757 = n43756 ^ n43753;
  assign n44474 = n43703 ^ n43510;
  assign n44472 = n42318 ^ n41684;
  assign n44473 = n44472 ^ n43161;
  assign n44475 = n44474 ^ n44473;
  assign n44184 = n43700 ^ n43515;
  assign n44034 = n42495 ^ n41831;
  assign n44035 = n44034 ^ n43172;
  assign n44033 = n43697 ^ n43520;
  assign n44036 = n44035 ^ n44033;
  assign n44026 = n43694 ^ n43691;
  assign n44019 = n43686 ^ n43525;
  assign n43762 = n42501 ^ n41853;
  assign n43764 = n43763 ^ n43762;
  assign n43761 = n43683 ^ n43530;
  assign n43765 = n43764 ^ n43761;
  assign n43769 = n43680 ^ n43535;
  assign n43766 = n43196 ^ n42537;
  assign n43768 = n43767 ^ n43766;
  assign n43770 = n43769 ^ n43768;
  assign n44006 = n43677 ^ n43540;
  assign n43773 = n43674 ^ n43671;
  assign n43771 = n43008 ^ n42404;
  assign n43772 = n43771 ^ n43737;
  assign n43774 = n43773 ^ n43772;
  assign n43996 = n43666 ^ n43663;
  assign n43989 = n43658 ^ n43545;
  assign n43776 = n42332 ^ n42290;
  assign n43777 = n43776 ^ n43439;
  assign n43775 = n43655 ^ n43550;
  assign n43778 = n43777 ^ n43775;
  assign n43780 = n42870 ^ n42344;
  assign n43781 = n43780 ^ n43307;
  assign n43779 = n43649 ^ n43560;
  assign n43782 = n43781 ^ n43779;
  assign n43784 = n42834 ^ n42280;
  assign n43785 = n43784 ^ n42874;
  assign n43783 = n43646 ^ n43565;
  assign n43786 = n43785 ^ n43783;
  assign n43790 = n43635 ^ n1811;
  assign n43788 = n42907 ^ n42038;
  assign n43789 = n43788 ^ n43290;
  assign n43791 = n43790 ^ n43789;
  assign n43961 = n43960 ^ n43792;
  assign n43962 = ~n43795 & ~n43961;
  assign n43963 = n43962 ^ n43794;
  assign n43964 = n43963 ^ n43790;
  assign n43965 = n43791 & ~n43964;
  assign n43966 = n43965 ^ n43789;
  assign n43787 = n43643 ^ n43640;
  assign n43967 = n43966 ^ n43787;
  assign n43968 = n42875 ^ n42092;
  assign n43969 = n43968 ^ n43297;
  assign n43970 = n43969 ^ n43787;
  assign n43971 = n43967 & ~n43970;
  assign n43972 = n43971 ^ n43969;
  assign n43973 = n43972 ^ n43783;
  assign n43974 = ~n43786 & ~n43973;
  assign n43975 = n43974 ^ n43785;
  assign n43976 = n43975 ^ n43779;
  assign n43977 = n43782 & ~n43976;
  assign n43978 = n43977 ^ n43781;
  assign n43980 = n43979 ^ n43978;
  assign n43981 = n42866 ^ n42338;
  assign n43982 = n43981 ^ n43314;
  assign n43983 = n43982 ^ n43979;
  assign n43984 = n43980 & n43983;
  assign n43985 = n43984 ^ n43982;
  assign n43986 = n43985 ^ n43775;
  assign n43987 = n43778 & ~n43986;
  assign n43988 = n43987 ^ n43777;
  assign n43990 = n43989 ^ n43988;
  assign n43991 = n43498 ^ n42326;
  assign n43992 = n43991 ^ n42935;
  assign n43993 = n43992 ^ n43989;
  assign n43994 = ~n43990 & ~n43993;
  assign n43995 = n43994 ^ n43992;
  assign n43997 = n43996 ^ n43995;
  assign n43998 = n42288 ^ n42286;
  assign n43999 = n43998 ^ n43715;
  assign n44000 = n43999 ^ n43996;
  assign n44001 = ~n43997 & ~n44000;
  assign n44002 = n44001 ^ n43999;
  assign n44003 = n44002 ^ n43772;
  assign n44004 = n43774 & n44003;
  assign n44005 = n44004 ^ n43773;
  assign n44007 = n44006 ^ n44005;
  assign n44008 = n43148 ^ n41596;
  assign n44009 = n44008 ^ n43832;
  assign n44010 = n44009 ^ n44006;
  assign n44011 = n44007 & ~n44010;
  assign n44012 = n44011 ^ n44009;
  assign n44013 = n44012 ^ n43769;
  assign n44014 = ~n43770 & n44013;
  assign n44015 = n44014 ^ n43768;
  assign n44016 = n44015 ^ n43761;
  assign n44017 = n43765 & ~n44016;
  assign n44018 = n44017 ^ n43764;
  assign n44020 = n44019 ^ n44018;
  assign n44021 = n43913 ^ n41843;
  assign n44022 = n44021 ^ n42504;
  assign n44023 = n44022 ^ n44019;
  assign n44024 = n44020 & ~n44023;
  assign n44025 = n44024 ^ n44022;
  assign n44027 = n44026 ^ n44025;
  assign n44028 = n43167 ^ n42508;
  assign n44029 = n44028 ^ n41841;
  assign n44030 = n44029 ^ n44026;
  assign n44031 = n44027 & ~n44030;
  assign n44032 = n44031 ^ n44029;
  assign n44181 = n44033 ^ n44032;
  assign n44182 = ~n44036 & ~n44181;
  assign n44183 = n44182 ^ n44035;
  assign n44185 = n44184 ^ n44183;
  assign n44179 = n42542 ^ n41829;
  assign n44180 = n44179 ^ n43176;
  assign n44469 = n44184 ^ n44180;
  assign n44470 = ~n44185 & ~n44469;
  assign n44471 = n44470 ^ n44180;
  assign n44526 = n44474 ^ n44471;
  assign n44527 = n44475 & n44526;
  assign n44528 = n44527 ^ n44473;
  assign n44476 = n44475 ^ n44471;
  assign n44477 = n44476 ^ n40763;
  assign n44186 = n44185 ^ n44180;
  assign n44187 = n44186 ^ n41092;
  assign n44037 = n44036 ^ n44032;
  assign n44038 = n44037 ^ n41094;
  assign n44039 = n44029 ^ n44027;
  assign n44040 = n44039 ^ n41104;
  assign n44041 = n44022 ^ n44020;
  assign n44042 = n44041 ^ n41110;
  assign n44043 = n44015 ^ n43765;
  assign n44044 = n44043 ^ n41112;
  assign n44045 = n44012 ^ n43770;
  assign n44046 = n44045 ^ n41824;
  assign n44047 = n44009 ^ n44007;
  assign n44048 = n44047 ^ n41597;
  assign n44049 = n43999 ^ n43997;
  assign n44050 = n44049 ^ n41698;
  assign n44051 = n43992 ^ n43990;
  assign n44052 = n44051 ^ n41704;
  assign n44053 = n43985 ^ n43778;
  assign n44054 = n44053 ^ n41710;
  assign n44055 = n43982 ^ n43980;
  assign n44056 = n44055 ^ n41582;
  assign n44057 = n43975 ^ n43782;
  assign n44058 = n44057 ^ n41332;
  assign n44059 = n43972 ^ n43786;
  assign n44060 = n44059 ^ n41189;
  assign n44061 = n43969 ^ n43967;
  assign n44062 = n44061 ^ n40656;
  assign n44063 = n43963 ^ n43791;
  assign n44064 = n44063 ^ n40659;
  assign n44127 = n44126 ^ n40666;
  assign n44129 = n44128 ^ n44126;
  assign n44130 = ~n44127 & ~n44129;
  assign n44131 = n44130 ^ n40666;
  assign n44132 = n44131 ^ n44063;
  assign n44133 = ~n44064 & n44132;
  assign n44134 = n44133 ^ n40659;
  assign n44135 = n44134 ^ n44061;
  assign n44136 = n44062 & ~n44135;
  assign n44137 = n44136 ^ n40656;
  assign n44138 = n44137 ^ n44059;
  assign n44139 = n44060 & ~n44138;
  assign n44140 = n44139 ^ n41189;
  assign n44141 = n44140 ^ n44057;
  assign n44142 = n44058 & ~n44141;
  assign n44143 = n44142 ^ n41332;
  assign n44144 = n44143 ^ n44055;
  assign n44145 = ~n44056 & ~n44144;
  assign n44146 = n44145 ^ n41582;
  assign n44147 = n44146 ^ n44053;
  assign n44148 = ~n44054 & ~n44147;
  assign n44149 = n44148 ^ n41710;
  assign n44150 = n44149 ^ n44051;
  assign n44151 = n44052 & ~n44150;
  assign n44152 = n44151 ^ n41704;
  assign n44153 = n44152 ^ n44049;
  assign n44154 = n44050 & n44153;
  assign n44155 = n44154 ^ n41698;
  assign n44156 = n44155 ^ n41728;
  assign n44157 = n44002 ^ n43774;
  assign n44158 = n44157 ^ n44155;
  assign n44159 = ~n44156 & ~n44158;
  assign n44160 = n44159 ^ n41728;
  assign n44161 = n44160 ^ n44047;
  assign n44162 = ~n44048 & n44161;
  assign n44163 = n44162 ^ n41597;
  assign n44164 = n44163 ^ n44045;
  assign n44165 = ~n44046 & n44164;
  assign n44166 = n44165 ^ n41824;
  assign n44167 = n44166 ^ n44043;
  assign n44168 = ~n44044 & ~n44167;
  assign n44169 = n44168 ^ n41112;
  assign n44170 = n44169 ^ n44041;
  assign n44171 = n44042 & ~n44170;
  assign n44172 = n44171 ^ n41110;
  assign n44173 = n44172 ^ n44039;
  assign n44174 = n44040 & ~n44173;
  assign n44175 = n44174 ^ n41104;
  assign n44176 = n44175 ^ n44037;
  assign n44177 = n44038 & ~n44176;
  assign n44178 = n44177 ^ n41094;
  assign n44466 = n44186 ^ n44178;
  assign n44467 = ~n44187 & n44466;
  assign n44468 = n44467 ^ n41092;
  assign n44478 = n44477 ^ n44468;
  assign n44188 = n44187 ^ n44178;
  assign n44189 = n44175 ^ n44038;
  assign n44190 = n44166 ^ n44044;
  assign n44191 = n44160 ^ n44048;
  assign n44192 = n44157 ^ n41728;
  assign n44193 = n44192 ^ n44155;
  assign n44194 = n44149 ^ n44052;
  assign n44195 = n44146 ^ n44054;
  assign n44221 = n44218 & n44220;
  assign n44222 = n44131 ^ n44064;
  assign n44223 = ~n44221 & n44222;
  assign n44224 = n44134 ^ n44062;
  assign n44225 = n44223 & ~n44224;
  assign n44226 = n44137 ^ n44060;
  assign n44227 = ~n44225 & n44226;
  assign n44228 = n44140 ^ n44058;
  assign n44229 = ~n44227 & ~n44228;
  assign n44230 = n44143 ^ n44056;
  assign n44231 = ~n44229 & ~n44230;
  assign n44232 = n44195 & n44231;
  assign n44233 = n44194 & n44232;
  assign n44234 = n44152 ^ n44050;
  assign n44235 = ~n44233 & ~n44234;
  assign n44236 = ~n44193 & n44235;
  assign n44237 = ~n44191 & ~n44236;
  assign n44238 = n44163 ^ n44046;
  assign n44239 = n44237 & ~n44238;
  assign n44240 = n44190 & ~n44239;
  assign n44241 = n44169 ^ n44042;
  assign n44242 = ~n44240 & ~n44241;
  assign n44243 = n44172 ^ n44040;
  assign n44244 = ~n44242 & n44243;
  assign n44245 = ~n44189 & ~n44244;
  assign n44479 = n44188 & n44245;
  assign n44521 = n44478 & ~n44479;
  assign n44518 = n42477 ^ n2524;
  assign n44519 = n44518 ^ n38477;
  assign n44520 = n44519 ^ n32369;
  assign n44522 = n44521 ^ n44520;
  assign n44523 = n44522 ^ n43910;
  assign n44517 = n43725 ^ n43722;
  assign n44524 = n44523 ^ n44517;
  assign n44525 = n44524 ^ n42312;
  assign n44529 = n44528 ^ n44525;
  assign n44514 = n44476 ^ n44468;
  assign n44515 = n44477 & n44514;
  assign n44516 = n44515 ^ n40763;
  assign n44530 = n44529 ^ n44516;
  assign n44531 = n44530 ^ n43208;
  assign n44480 = n44479 ^ n44478;
  assign n44246 = n44245 ^ n44188;
  assign n43758 = n42468 ^ n34136;
  assign n43759 = n43758 ^ n38815;
  assign n43760 = n43759 ^ n32494;
  assign n44247 = n44246 ^ n43760;
  assign n44249 = n42460 ^ n34142;
  assign n44250 = n44249 ^ n38721;
  assign n44251 = n44250 ^ n32472;
  assign n44248 = n44244 ^ n44189;
  assign n44252 = n44251 ^ n44248;
  assign n44256 = n44243 ^ n44242;
  assign n44253 = n42432 ^ n34147;
  assign n44254 = n44253 ^ n38725;
  assign n44255 = n44254 ^ n1229;
  assign n44257 = n44256 ^ n44255;
  assign n44444 = n44239 ^ n44190;
  assign n44261 = n44238 ^ n44237;
  assign n906 = n905 ^ n869;
  assign n934 = n933 ^ n906;
  assign n941 = n940 ^ n934;
  assign n44262 = n44261 ^ n941;
  assign n44264 = n38738 ^ n34174;
  assign n44265 = n44264 ^ n42099;
  assign n44266 = n44265 ^ n932;
  assign n44263 = n44236 ^ n44191;
  assign n44267 = n44266 ^ n44263;
  assign n44269 = n42104 ^ n801;
  assign n44270 = n44269 ^ n38743;
  assign n44271 = n44270 ^ n32415;
  assign n44268 = n44235 ^ n44193;
  assign n44272 = n44271 ^ n44268;
  assign n44274 = n42109 ^ n34154;
  assign n44275 = n44274 ^ n38747;
  assign n44276 = n44275 ^ n32420;
  assign n44273 = n44234 ^ n44233;
  assign n44277 = n44276 ^ n44273;
  assign n44281 = n44232 ^ n44194;
  assign n44278 = n42114 ^ n34167;
  assign n44279 = n44278 ^ n38752;
  assign n44280 = n44279 ^ n32404;
  assign n44282 = n44281 ^ n44280;
  assign n44421 = n44231 ^ n44195;
  assign n44286 = n44230 ^ n44229;
  assign n44283 = n42118 ^ n33775;
  assign n44284 = n44283 ^ n38758;
  assign n44285 = n44284 ^ n32397;
  assign n44287 = n44286 ^ n44285;
  assign n44289 = n42240 ^ n33634;
  assign n44290 = n44289 ^ n38767;
  assign n44291 = n44290 ^ n32391;
  assign n44288 = n44228 ^ n44227;
  assign n44292 = n44291 ^ n44288;
  assign n44293 = n44226 ^ n44225;
  assign n44297 = n44296 ^ n44293;
  assign n44299 = n42229 ^ n33644;
  assign n44300 = n44299 ^ n38351;
  assign n44301 = n44300 ^ n31980;
  assign n44298 = n44224 ^ n44223;
  assign n44302 = n44301 ^ n44298;
  assign n44303 = n44222 ^ n44221;
  assign n44307 = n44306 ^ n44303;
  assign n44403 = n44402 ^ n44308;
  assign n44404 = n44309 & ~n44403;
  assign n44405 = n44404 ^ n2216;
  assign n44406 = n44405 ^ n44303;
  assign n44407 = n44307 & ~n44406;
  assign n44408 = n44407 ^ n44306;
  assign n44409 = n44408 ^ n44298;
  assign n44410 = n44302 & ~n44409;
  assign n44411 = n44410 ^ n44301;
  assign n44412 = n44411 ^ n44293;
  assign n44413 = ~n44297 & n44412;
  assign n44414 = n44413 ^ n44296;
  assign n44415 = n44414 ^ n44291;
  assign n44416 = ~n44292 & ~n44415;
  assign n44417 = n44416 ^ n44288;
  assign n44418 = n44417 ^ n44286;
  assign n44419 = n44287 & n44418;
  assign n44420 = n44419 ^ n44285;
  assign n44422 = n44421 ^ n44420;
  assign n44423 = n42251 ^ n34159;
  assign n44424 = n44423 ^ n38778;
  assign n44425 = n44424 ^ n32387;
  assign n44426 = n44425 ^ n44421;
  assign n44427 = ~n44422 & n44426;
  assign n44428 = n44427 ^ n44425;
  assign n44429 = n44428 ^ n44281;
  assign n44430 = n44282 & ~n44429;
  assign n44431 = n44430 ^ n44280;
  assign n44432 = n44431 ^ n44273;
  assign n44433 = ~n44277 & n44432;
  assign n44434 = n44433 ^ n44276;
  assign n44435 = n44434 ^ n44268;
  assign n44436 = n44272 & ~n44435;
  assign n44437 = n44436 ^ n44271;
  assign n44438 = n44437 ^ n44263;
  assign n44439 = n44267 & ~n44438;
  assign n44440 = n44439 ^ n44266;
  assign n44441 = n44440 ^ n941;
  assign n44442 = ~n44262 & ~n44441;
  assign n44443 = n44442 ^ n44261;
  assign n44445 = n44444 ^ n44443;
  assign n44446 = n42437 ^ n34216;
  assign n44447 = n44446 ^ n38731;
  assign n44448 = n44447 ^ n1063;
  assign n44449 = n44448 ^ n44444;
  assign n44450 = n44445 & n44449;
  assign n44451 = n44450 ^ n44448;
  assign n44258 = n42449 ^ n34221;
  assign n44259 = n44258 ^ n1064;
  assign n44260 = n44259 ^ n32466;
  assign n44452 = n44451 ^ n44260;
  assign n44453 = n44241 ^ n44240;
  assign n44454 = n44453 ^ n44451;
  assign n44455 = n44452 & ~n44454;
  assign n44456 = n44455 ^ n44260;
  assign n44457 = n44456 ^ n44256;
  assign n44458 = n44257 & ~n44457;
  assign n44459 = n44458 ^ n44255;
  assign n44460 = n44459 ^ n44248;
  assign n44461 = n44252 & ~n44460;
  assign n44462 = n44461 ^ n44251;
  assign n44463 = n44462 ^ n44246;
  assign n44464 = n44247 & ~n44463;
  assign n44465 = n44464 ^ n43760;
  assign n44481 = n44480 ^ n44465;
  assign n44482 = n42427 ^ n34132;
  assign n44483 = n44482 ^ n38716;
  assign n44484 = n44483 ^ n32499;
  assign n44511 = n44484 ^ n44480;
  assign n44512 = ~n44481 & n44511;
  assign n44513 = n44512 ^ n44484;
  assign n44532 = n44531 ^ n44513;
  assign n44486 = n43243 ^ n42302;
  assign n44487 = n44486 ^ n43804;
  assign n44485 = n44484 ^ n44481;
  assign n44488 = n44487 ^ n44485;
  assign n44491 = n43932 ^ n43236;
  assign n44492 = n44491 ^ n42561;
  assign n44489 = n44462 ^ n43760;
  assign n44490 = n44489 ^ n44246;
  assign n44493 = n44492 ^ n44490;
  assign n44496 = n43222 ^ n42308;
  assign n44497 = n44496 ^ n43815;
  assign n44498 = n44456 ^ n44257;
  assign n44499 = ~n44497 & n44498;
  assign n44494 = n43229 ^ n42304;
  assign n44495 = n44494 ^ n43809;
  assign n44500 = n44499 ^ n44495;
  assign n44501 = n44459 ^ n44252;
  assign n44502 = n44501 ^ n44495;
  assign n44503 = n44500 & ~n44502;
  assign n44504 = n44503 ^ n44499;
  assign n44505 = n44504 ^ n44490;
  assign n44506 = n44493 & ~n44505;
  assign n44507 = n44506 ^ n44492;
  assign n44508 = n44507 ^ n44485;
  assign n44509 = n44488 & ~n44508;
  assign n44510 = n44509 ^ n44487;
  assign n44533 = n44532 ^ n44510;
  assign n44534 = n42854 ^ n42298;
  assign n44535 = n44534 ^ n43803;
  assign n44536 = n44535 ^ n44532;
  assign n44537 = ~n44533 & n44536;
  assign n44538 = n44537 ^ n44535;
  assign n44539 = n44538 ^ n43753;
  assign n44540 = ~n43757 & n44539;
  assign n44541 = n44540 ^ n43756;
  assign n44582 = n44543 ^ n44541;
  assign n44583 = ~n44546 & ~n44582;
  assign n44584 = n44583 ^ n44545;
  assign n44581 = n44349 ^ n44341;
  assign n44585 = n44584 ^ n44581;
  assign n44579 = n42839 ^ n42584;
  assign n44580 = n44579 ^ n43796;
  assign n44586 = n44585 ^ n44580;
  assign n44587 = n44586 ^ n41629;
  assign n44547 = n44546 ^ n44541;
  assign n44548 = n44547 ^ n41639;
  assign n44549 = n44538 ^ n43757;
  assign n44550 = n44549 ^ n41641;
  assign n44551 = n44535 ^ n44533;
  assign n44552 = n44551 ^ n41647;
  assign n44553 = n44507 ^ n44488;
  assign n44554 = n44553 ^ n41657;
  assign n44555 = n44504 ^ n44493;
  assign n44556 = n44555 ^ n41663;
  assign n44557 = n44498 ^ n44497;
  assign n44558 = n41672 & ~n44557;
  assign n44559 = n44558 ^ n41666;
  assign n44560 = n44501 ^ n44500;
  assign n44561 = n44560 ^ n44558;
  assign n44562 = n44559 & ~n44561;
  assign n44563 = n44562 ^ n41666;
  assign n44564 = n44563 ^ n44555;
  assign n44565 = ~n44556 & ~n44564;
  assign n44566 = n44565 ^ n41663;
  assign n44567 = n44566 ^ n44553;
  assign n44568 = ~n44554 & n44567;
  assign n44569 = n44568 ^ n41657;
  assign n44570 = n44569 ^ n44551;
  assign n44571 = ~n44552 & n44570;
  assign n44572 = n44571 ^ n41647;
  assign n44573 = n44572 ^ n44549;
  assign n44574 = ~n44550 & ~n44573;
  assign n44575 = n44574 ^ n41641;
  assign n44576 = n44575 ^ n44547;
  assign n44577 = ~n44548 & n44576;
  assign n44578 = n44577 ^ n41639;
  assign n44588 = n44587 ^ n44578;
  assign n44589 = n44572 ^ n44550;
  assign n44590 = n44569 ^ n44552;
  assign n44591 = n44566 ^ n44554;
  assign n44592 = n44563 ^ n44556;
  assign n44593 = n44560 ^ n44559;
  assign n44594 = n44592 & ~n44593;
  assign n44595 = n44591 & ~n44594;
  assign n44596 = ~n44590 & ~n44595;
  assign n44597 = n44589 & ~n44596;
  assign n44598 = n44575 ^ n44548;
  assign n44599 = ~n44597 & n44598;
  assign n44600 = n44588 & n44599;
  assign n44608 = n42838 ^ n42665;
  assign n44609 = n44608 ^ n43792;
  assign n44607 = n44352 ^ n44336;
  assign n44610 = n44609 ^ n44607;
  assign n44604 = n44581 ^ n44580;
  assign n44605 = n44585 & n44604;
  assign n44606 = n44605 ^ n44580;
  assign n44611 = n44610 ^ n44606;
  assign n44612 = n44611 ^ n41627;
  assign n44601 = n44586 ^ n44578;
  assign n44602 = ~n44587 & n44601;
  assign n44603 = n44602 ^ n41629;
  assign n44613 = n44612 ^ n44603;
  assign n44614 = n44600 & n44613;
  assign n44623 = n44355 ^ n44331;
  assign n44620 = n44607 ^ n44606;
  assign n44621 = ~n44610 & ~n44620;
  assign n44622 = n44621 ^ n44609;
  assign n44624 = n44623 ^ n44622;
  assign n44618 = n43271 ^ n42821;
  assign n44619 = n44618 ^ n43790;
  assign n44625 = n44624 ^ n44619;
  assign n44626 = n44625 ^ n41617;
  assign n44615 = n44611 ^ n44603;
  assign n44616 = ~n44612 & n44615;
  assign n44617 = n44616 ^ n41627;
  assign n44627 = n44626 ^ n44617;
  assign n44628 = ~n44614 & ~n44627;
  assign n44636 = n42850 ^ n42837;
  assign n44637 = n44636 ^ n43787;
  assign n44635 = n44363 ^ n44360;
  assign n44638 = n44637 ^ n44635;
  assign n44632 = n44623 ^ n44619;
  assign n44633 = n44624 & ~n44632;
  assign n44634 = n44633 ^ n44619;
  assign n44639 = n44638 ^ n44634;
  assign n44640 = n44639 ^ n41615;
  assign n44629 = n44625 ^ n44617;
  assign n44630 = ~n44626 & ~n44629;
  assign n44631 = n44630 ^ n41617;
  assign n44641 = n44640 ^ n44631;
  assign n44739 = n44628 & ~n44641;
  assign n44732 = n44635 ^ n44634;
  assign n44733 = n44638 & n44732;
  assign n44734 = n44733 ^ n44637;
  assign n44731 = n44366 ^ n44326;
  assign n44735 = n44734 ^ n44731;
  assign n44729 = n42845 ^ n42836;
  assign n44730 = n44729 ^ n43783;
  assign n44736 = n44735 ^ n44730;
  assign n44737 = n44736 ^ n41609;
  assign n44726 = n44639 ^ n44631;
  assign n44727 = n44640 & ~n44726;
  assign n44728 = n44727 ^ n41615;
  assign n44738 = n44737 ^ n44728;
  assign n44740 = n44739 ^ n44738;
  assign n44744 = n44743 ^ n44740;
  assign n44643 = n42793 ^ n34732;
  assign n44644 = n44643 ^ n39193;
  assign n44645 = n44644 ^ n32747;
  assign n44642 = n44641 ^ n44628;
  assign n44646 = n44645 ^ n44642;
  assign n44715 = n44627 ^ n44614;
  assign n44648 = n42782 ^ n34742;
  assign n44649 = n44648 ^ n1685;
  assign n44650 = n44649 ^ n32668;
  assign n44647 = n44613 ^ n44600;
  assign n44651 = n44650 ^ n44647;
  assign n44704 = n44599 ^ n44588;
  assign n44655 = n44598 ^ n44597;
  assign n44652 = n42771 ^ n1592;
  assign n44653 = n44652 ^ n39204;
  assign n44654 = n44653 ^ n32680;
  assign n44656 = n44655 ^ n44654;
  assign n44693 = n44596 ^ n44589;
  assign n44657 = n44595 ^ n44590;
  assign n44661 = n44660 ^ n44657;
  assign n44663 = n42743 ^ n34763;
  assign n44664 = n44663 ^ n39214;
  assign n44665 = n44664 ^ n32691;
  assign n44662 = n44594 ^ n44591;
  assign n44666 = n44665 ^ n44662;
  assign n44670 = n44593 ^ n44592;
  assign n44667 = n42753 ^ n34772;
  assign n44668 = n44667 ^ n39218;
  assign n44669 = n44668 ^ n32700;
  assign n44671 = n44670 ^ n44669;
  assign n44677 = n42749 ^ n34767;
  assign n44678 = n44677 ^ n39221;
  assign n44679 = n44678 ^ n32696;
  assign n44672 = n43204 ^ n35028;
  assign n44673 = n44672 ^ n39440;
  assign n44674 = n44673 ^ n33369;
  assign n44675 = n44557 ^ n41672;
  assign n44676 = n44674 & ~n44675;
  assign n44680 = n44679 ^ n44676;
  assign n44681 = n44676 ^ n44593;
  assign n44682 = n44680 & n44681;
  assign n44683 = n44682 ^ n44679;
  assign n44684 = n44683 ^ n44670;
  assign n44685 = n44671 & ~n44684;
  assign n44686 = n44685 ^ n44669;
  assign n44687 = n44686 ^ n44662;
  assign n44688 = ~n44666 & n44687;
  assign n44689 = n44688 ^ n44665;
  assign n44690 = n44689 ^ n44657;
  assign n44691 = ~n44661 & n44690;
  assign n44692 = n44691 ^ n44660;
  assign n44694 = n44693 ^ n44692;
  assign n44695 = n42734 ^ n34753;
  assign n44696 = n44695 ^ n39210;
  assign n44697 = n44696 ^ n32675;
  assign n44698 = n44697 ^ n44693;
  assign n44699 = n44694 & ~n44698;
  assign n44700 = n44699 ^ n44697;
  assign n44701 = n44700 ^ n44655;
  assign n44702 = n44656 & ~n44701;
  assign n44703 = n44702 ^ n44654;
  assign n44705 = n44704 ^ n44703;
  assign n44706 = n42728 ^ n34746;
  assign n44707 = n44706 ^ n39199;
  assign n44708 = n44707 ^ n1677;
  assign n44709 = n44708 ^ n44704;
  assign n44710 = n44705 & ~n44709;
  assign n44711 = n44710 ^ n44708;
  assign n44712 = n44711 ^ n44647;
  assign n44713 = ~n44651 & n44712;
  assign n44714 = n44713 ^ n44650;
  assign n44716 = n44715 ^ n44714;
  assign n44717 = n42723 ^ n34737;
  assign n44718 = n44717 ^ n39256;
  assign n44719 = n44718 ^ n1775;
  assign n44720 = n44719 ^ n44715;
  assign n44721 = ~n44716 & n44720;
  assign n44722 = n44721 ^ n44719;
  assign n44723 = n44722 ^ n44642;
  assign n44724 = ~n44646 & n44723;
  assign n44725 = n44724 ^ n44645;
  assign n44745 = n44744 ^ n44725;
  assign n45708 = n45707 ^ n44745;
  assign n44885 = n43763 ^ n43148;
  assign n44886 = n44885 ^ n44033;
  assign n44814 = n44414 ^ n44292;
  assign n44812 = n43767 ^ n43008;
  assign n44813 = n44812 ^ n44026;
  assign n44815 = n44814 ^ n44813;
  assign n44816 = n43832 ^ n42286;
  assign n44817 = n44816 ^ n44019;
  assign n44746 = n44411 ^ n44297;
  assign n44818 = n44817 ^ n44746;
  assign n44819 = n43715 ^ n42290;
  assign n44820 = n44819 ^ n43769;
  assign n44757 = n44405 ^ n44307;
  assign n44821 = n44820 ^ n44757;
  assign n44844 = n44393 ^ n44321;
  assign n44825 = n44374 ^ n44371;
  assign n44822 = n44731 ^ n44730;
  assign n44823 = ~n44735 & ~n44822;
  assign n44824 = n44823 ^ n44730;
  assign n44826 = n44825 ^ n44824;
  assign n44827 = n43290 ^ n42840;
  assign n44828 = n44827 ^ n43779;
  assign n44829 = n44828 ^ n44825;
  assign n44830 = ~n44826 & n44829;
  assign n44831 = n44830 ^ n44828;
  assign n44781 = n44382 ^ n44379;
  assign n44832 = n44831 ^ n44781;
  assign n44833 = n43297 ^ n42900;
  assign n44834 = n44833 ^ n43979;
  assign n44835 = n44834 ^ n44781;
  assign n44836 = ~n44832 & n44835;
  assign n44837 = n44836 ^ n44834;
  assign n44776 = n44390 ^ n44387;
  assign n44838 = n44837 ^ n44776;
  assign n44839 = n42907 ^ n42834;
  assign n44840 = n44839 ^ n43775;
  assign n44841 = n44840 ^ n44776;
  assign n44842 = ~n44838 & n44841;
  assign n44843 = n44842 ^ n44840;
  assign n44845 = n44844 ^ n44843;
  assign n44846 = n43307 ^ n42875;
  assign n44847 = n44846 ^ n43989;
  assign n44848 = n44847 ^ n44844;
  assign n44849 = ~n44845 & ~n44848;
  assign n44850 = n44849 ^ n44847;
  assign n44771 = n44396 ^ n44316;
  assign n44851 = n44850 ^ n44771;
  assign n44852 = n43314 ^ n42874;
  assign n44853 = n44852 ^ n43996;
  assign n44854 = n44853 ^ n44771;
  assign n44855 = n44851 & n44854;
  assign n44856 = n44855 ^ n44853;
  assign n44765 = n44399 ^ n44314;
  assign n44857 = n44856 ^ n44765;
  assign n44858 = n43439 ^ n42870;
  assign n44859 = n44858 ^ n43773;
  assign n44860 = n44859 ^ n44765;
  assign n44861 = ~n44857 & n44860;
  assign n44862 = n44861 ^ n44859;
  assign n44863 = n44862 ^ n44762;
  assign n44864 = n43498 ^ n42866;
  assign n44865 = n44864 ^ n44006;
  assign n44866 = n44865 ^ n44762;
  assign n44867 = n44863 & ~n44866;
  assign n44868 = n44867 ^ n44865;
  assign n44869 = n44868 ^ n44757;
  assign n44870 = ~n44821 & n44869;
  assign n44871 = n44870 ^ n44820;
  assign n44752 = n44408 ^ n44302;
  assign n44872 = n44871 ^ n44752;
  assign n44873 = n43737 ^ n42935;
  assign n44874 = n44873 ^ n43761;
  assign n44875 = n44874 ^ n44752;
  assign n44876 = n44872 & ~n44875;
  assign n44877 = n44876 ^ n44874;
  assign n44878 = n44877 ^ n44746;
  assign n44879 = n44818 & ~n44878;
  assign n44880 = n44879 ^ n44817;
  assign n44881 = n44880 ^ n44814;
  assign n44882 = n44815 & ~n44881;
  assign n44883 = n44882 ^ n44813;
  assign n44811 = n44417 ^ n44287;
  assign n44884 = n44883 ^ n44811;
  assign n44922 = n44886 ^ n44884;
  assign n44923 = n44922 ^ n41596;
  assign n44924 = n44880 ^ n44815;
  assign n44925 = n44924 ^ n42404;
  assign n44926 = n44877 ^ n44818;
  assign n44927 = n44926 ^ n42288;
  assign n44928 = n44874 ^ n44872;
  assign n44929 = n44928 ^ n42326;
  assign n44930 = n44868 ^ n44821;
  assign n44931 = n44930 ^ n42332;
  assign n44932 = n44865 ^ n44863;
  assign n44933 = n44932 ^ n42338;
  assign n44934 = n44859 ^ n44857;
  assign n44935 = n44934 ^ n42344;
  assign n44936 = n44853 ^ n44851;
  assign n44937 = n44936 ^ n42280;
  assign n44938 = n44847 ^ n44845;
  assign n44939 = n44938 ^ n42092;
  assign n44940 = n44840 ^ n44838;
  assign n44941 = n44940 ^ n42038;
  assign n44942 = n44834 ^ n44832;
  assign n44943 = n44942 ^ n41917;
  assign n44944 = n44828 ^ n44826;
  assign n44945 = n44944 ^ n41603;
  assign n44946 = n44736 ^ n44728;
  assign n44947 = n44737 & ~n44946;
  assign n44948 = n44947 ^ n41609;
  assign n44949 = n44948 ^ n44944;
  assign n44950 = ~n44945 & ~n44949;
  assign n44951 = n44950 ^ n41603;
  assign n44952 = n44951 ^ n44942;
  assign n44953 = n44943 & n44952;
  assign n44954 = n44953 ^ n41917;
  assign n44955 = n44954 ^ n44940;
  assign n44956 = n44941 & ~n44955;
  assign n44957 = n44956 ^ n42038;
  assign n44958 = n44957 ^ n44938;
  assign n44959 = n44939 & n44958;
  assign n44960 = n44959 ^ n42092;
  assign n44961 = n44960 ^ n44936;
  assign n44962 = ~n44937 & ~n44961;
  assign n44963 = n44962 ^ n42280;
  assign n44964 = n44963 ^ n44934;
  assign n44965 = n44935 & ~n44964;
  assign n44966 = n44965 ^ n42344;
  assign n44967 = n44966 ^ n44932;
  assign n44968 = ~n44933 & n44967;
  assign n44969 = n44968 ^ n42338;
  assign n44970 = n44969 ^ n44930;
  assign n44971 = ~n44931 & n44970;
  assign n44972 = n44971 ^ n42332;
  assign n44973 = n44972 ^ n44928;
  assign n44974 = ~n44929 & n44973;
  assign n44975 = n44974 ^ n42326;
  assign n44976 = n44975 ^ n44926;
  assign n44977 = n44927 & ~n44976;
  assign n44978 = n44977 ^ n42288;
  assign n44979 = n44978 ^ n44924;
  assign n44980 = n44925 & ~n44979;
  assign n44981 = n44980 ^ n42404;
  assign n44982 = n44981 ^ n44922;
  assign n44983 = n44923 & n44982;
  assign n44984 = n44983 ^ n41596;
  assign n44887 = n44886 ^ n44811;
  assign n44888 = ~n44884 & ~n44887;
  assign n44889 = n44888 ^ n44886;
  assign n44808 = n43913 ^ n43196;
  assign n44809 = n44808 ^ n44184;
  assign n44807 = n44425 ^ n44422;
  assign n44810 = n44809 ^ n44807;
  assign n44920 = n44889 ^ n44810;
  assign n44921 = n44920 ^ n42537;
  assign n45011 = n44984 ^ n44921;
  assign n45012 = n44981 ^ n44923;
  assign n45013 = n44978 ^ n44925;
  assign n45014 = n44975 ^ n44927;
  assign n45015 = n44969 ^ n44931;
  assign n45016 = n44957 ^ n42092;
  assign n45017 = n45016 ^ n44938;
  assign n45018 = n44954 ^ n42038;
  assign n45019 = n45018 ^ n44940;
  assign n45020 = n44948 ^ n44945;
  assign n45021 = ~n44738 & n44739;
  assign n45022 = n45020 & n45021;
  assign n45023 = n44951 ^ n44943;
  assign n45024 = n45022 & n45023;
  assign n45025 = n45019 & ~n45024;
  assign n45026 = n45017 & n45025;
  assign n45027 = n44960 ^ n44937;
  assign n45028 = ~n45026 & ~n45027;
  assign n45029 = n44963 ^ n44935;
  assign n45030 = ~n45028 & n45029;
  assign n45031 = n44966 ^ n44933;
  assign n45032 = ~n45030 & n45031;
  assign n45033 = n45015 & n45032;
  assign n45034 = n44972 ^ n44929;
  assign n45035 = n45033 & n45034;
  assign n45036 = n45014 & ~n45035;
  assign n45037 = n45013 & n45036;
  assign n45038 = ~n45012 & ~n45037;
  assign n45039 = ~n45011 & n45038;
  assign n44985 = n44984 ^ n44920;
  assign n44986 = ~n44921 & n44985;
  assign n44987 = n44986 ^ n42537;
  assign n44890 = n44889 ^ n44807;
  assign n44891 = ~n44810 & ~n44890;
  assign n44892 = n44891 ^ n44809;
  assign n44804 = n43167 ^ n42501;
  assign n44805 = n44804 ^ n44474;
  assign n44803 = n44428 ^ n44282;
  assign n44806 = n44805 ^ n44803;
  assign n44918 = n44892 ^ n44806;
  assign n44919 = n44918 ^ n41853;
  assign n45040 = n44987 ^ n44919;
  assign n45041 = ~n45039 & ~n45040;
  assign n44988 = n44987 ^ n44918;
  assign n44989 = n44919 & n44988;
  assign n44990 = n44989 ^ n41853;
  assign n44898 = n43172 ^ n42504;
  assign n44899 = n44898 ^ n44517;
  assign n44896 = n44431 ^ n44277;
  assign n44893 = n44892 ^ n44803;
  assign n44894 = n44806 & n44893;
  assign n44895 = n44894 ^ n44805;
  assign n44897 = n44896 ^ n44895;
  assign n44916 = n44899 ^ n44897;
  assign n44917 = n44916 ^ n41843;
  assign n45042 = n44990 ^ n44917;
  assign n45043 = ~n45041 & ~n45042;
  assign n44991 = n44990 ^ n44916;
  assign n44992 = n44917 & n44991;
  assign n44993 = n44992 ^ n41843;
  assign n44905 = n43176 ^ n42508;
  assign n44906 = n44905 ^ n43745;
  assign n44903 = n44434 ^ n44272;
  assign n44900 = n44899 ^ n44896;
  assign n44901 = n44897 & n44900;
  assign n44902 = n44901 ^ n44899;
  assign n44904 = n44903 ^ n44902;
  assign n44914 = n44906 ^ n44904;
  assign n44915 = n44914 ^ n41841;
  assign n45044 = n44993 ^ n44915;
  assign n45045 = ~n45043 & n45044;
  assign n44994 = n44993 ^ n44914;
  assign n44995 = ~n44915 & ~n44994;
  assign n44996 = n44995 ^ n41841;
  assign n44910 = n44437 ^ n44267;
  assign n44907 = n44906 ^ n44903;
  assign n44908 = n44904 & ~n44907;
  assign n44909 = n44908 ^ n44906;
  assign n44911 = n44910 ^ n44909;
  assign n44801 = n43161 ^ n42495;
  assign n44802 = n44801 ^ n43840;
  assign n44912 = n44911 ^ n44802;
  assign n44913 = n44912 ^ n41831;
  assign n45010 = n44996 ^ n44913;
  assign n45049 = n45045 ^ n45010;
  assign n1338 = n1337 ^ n1253;
  assign n1354 = n1353 ^ n1338;
  assign n1361 = n1360 ^ n1354;
  assign n45050 = n45049 ^ n1361;
  assign n45171 = n45044 ^ n45043;
  assign n45051 = n45042 ^ n45041;
  assign n1156 = n1146 ^ n1098;
  assign n1181 = n1180 ^ n1156;
  assign n1188 = n1187 ^ n1181;
  assign n45052 = n45051 ^ n1188;
  assign n45054 = n43121 ^ n1021;
  assign n45055 = n45054 ^ n39339;
  assign n45056 = n45055 ^ n1172;
  assign n45053 = n45040 ^ n45039;
  assign n45057 = n45056 ^ n45053;
  assign n45157 = n45038 ^ n45011;
  assign n45058 = n45037 ^ n45012;
  assign n45062 = n45061 ^ n45058;
  assign n45146 = n45036 ^ n45013;
  assign n45064 = n43070 ^ n34687;
  assign n45065 = n45064 ^ n39307;
  assign n45066 = n45065 ^ n33280;
  assign n45063 = n45035 ^ n45014;
  assign n45067 = n45066 ^ n45063;
  assign n45069 = n43075 ^ n34692;
  assign n45070 = n45069 ^ n39153;
  assign n45071 = n45070 ^ n680;
  assign n45068 = n45034 ^ n45033;
  assign n45072 = n45071 ^ n45068;
  assign n45132 = n45032 ^ n45015;
  assign n45124 = n45031 ^ n45030;
  assign n45116 = n45029 ^ n45028;
  assign n45073 = n45027 ^ n45026;
  assign n45077 = n45076 ^ n45073;
  assign n45079 = n42705 ^ n34713;
  assign n45080 = n45079 ^ n39279;
  assign n45081 = n45080 ^ n33205;
  assign n45078 = n45025 ^ n45017;
  assign n45082 = n45081 ^ n45078;
  assign n45084 = n34718 ^ n2263;
  assign n45085 = n45084 ^ n39173;
  assign n45086 = n45085 ^ n33209;
  assign n45083 = n45024 ^ n45019;
  assign n45087 = n45086 ^ n45083;
  assign n45089 = n34722 ^ n2245;
  assign n45090 = n45089 ^ n39178;
  assign n45091 = n45090 ^ n33215;
  assign n45088 = n45023 ^ n45022;
  assign n45092 = n45091 ^ n45088;
  assign n45094 = n42714 ^ n2147;
  assign n45095 = n45094 ^ n39183;
  assign n45096 = n45095 ^ n33220;
  assign n45093 = n45021 ^ n45020;
  assign n45097 = n45096 ^ n45093;
  assign n45098 = n44740 ^ n44725;
  assign n45099 = ~n44744 & n45098;
  assign n45100 = n45099 ^ n44743;
  assign n45101 = n45100 ^ n45093;
  assign n45102 = n45097 & ~n45101;
  assign n45103 = n45102 ^ n45096;
  assign n45104 = n45103 ^ n45088;
  assign n45105 = n45092 & ~n45104;
  assign n45106 = n45105 ^ n45091;
  assign n45107 = n45106 ^ n45083;
  assign n45108 = n45087 & ~n45107;
  assign n45109 = n45108 ^ n45086;
  assign n45110 = n45109 ^ n45078;
  assign n45111 = ~n45082 & n45110;
  assign n45112 = n45111 ^ n45081;
  assign n45113 = n45112 ^ n45073;
  assign n45114 = n45077 & ~n45113;
  assign n45115 = n45114 ^ n45076;
  assign n45117 = n45116 ^ n45115;
  assign n45121 = n45120 ^ n45116;
  assign n45122 = ~n45117 & n45121;
  assign n45123 = n45122 ^ n45120;
  assign n45125 = n45124 ^ n45123;
  assign n45126 = n43086 ^ n34703;
  assign n45127 = n45126 ^ n39157;
  assign n45128 = n45127 ^ n33255;
  assign n45129 = n45128 ^ n45124;
  assign n45130 = n45125 & ~n45129;
  assign n45131 = n45130 ^ n45128;
  assign n45133 = n45132 ^ n45131;
  assign n45134 = n43081 ^ n34697;
  assign n45135 = n45134 ^ n39296;
  assign n45136 = n45135 ^ n33250;
  assign n45137 = n45136 ^ n45132;
  assign n45138 = ~n45133 & n45137;
  assign n45139 = n45138 ^ n45136;
  assign n45140 = n45139 ^ n45068;
  assign n45141 = n45072 & ~n45140;
  assign n45142 = n45141 ^ n45071;
  assign n45143 = n45142 ^ n45063;
  assign n45144 = n45067 & ~n45143;
  assign n45145 = n45144 ^ n45066;
  assign n45147 = n45146 ^ n45145;
  assign n45148 = n43066 ^ n34683;
  assign n45149 = n45148 ^ n39148;
  assign n45150 = n45149 ^ n33275;
  assign n45151 = n45150 ^ n45146;
  assign n45152 = n45147 & ~n45151;
  assign n45153 = n45152 ^ n45150;
  assign n45154 = n45153 ^ n45058;
  assign n45155 = n45062 & ~n45154;
  assign n45156 = n45155 ^ n45061;
  assign n45158 = n45157 ^ n45156;
  assign n45159 = n43061 ^ n1003;
  assign n45160 = n45159 ^ n39138;
  assign n45161 = n45160 ^ n33286;
  assign n45162 = n45161 ^ n45157;
  assign n45163 = n45158 & ~n45162;
  assign n45164 = n45163 ^ n45161;
  assign n45165 = n45164 ^ n45053;
  assign n45166 = ~n45057 & n45165;
  assign n45167 = n45166 ^ n45056;
  assign n45168 = n45167 ^ n45051;
  assign n45169 = n45052 & ~n45168;
  assign n45170 = n45169 ^ n1188;
  assign n45172 = n45171 ^ n45170;
  assign n45173 = n43053 ^ n34667;
  assign n45174 = n45173 ^ n1198;
  assign n45175 = n45174 ^ n1345;
  assign n45176 = n45175 ^ n45171;
  assign n45177 = ~n45172 & n45176;
  assign n45178 = n45177 ^ n45175;
  assign n45179 = n45178 ^ n45049;
  assign n45180 = n45050 & ~n45179;
  assign n45181 = n45180 ^ n1361;
  assign n45046 = ~n45010 & ~n45045;
  assign n45005 = n44440 ^ n44262;
  assign n45002 = n44910 ^ n44802;
  assign n45003 = n44911 & ~n45002;
  assign n45004 = n45003 ^ n44802;
  assign n45006 = n45005 ^ n45004;
  assign n45000 = n43208 ^ n42542;
  assign n45001 = n45000 ^ n43865;
  assign n45007 = n45006 ^ n45001;
  assign n45008 = n45007 ^ n41829;
  assign n44997 = n44996 ^ n44912;
  assign n44998 = n44913 & n44997;
  assign n44999 = n44998 ^ n41831;
  assign n45009 = n45008 ^ n44999;
  assign n45047 = n45046 ^ n45009;
  assign n44798 = n43048 ^ n34913;
  assign n44799 = n44798 ^ n39549;
  assign n44800 = n44799 ^ n2337;
  assign n45048 = n45047 ^ n44800;
  assign n45216 = n45181 ^ n45048;
  assign n45207 = n43932 ^ n43222;
  assign n45208 = n45207 ^ n43753;
  assign n45209 = n45175 ^ n45172;
  assign n45210 = ~n45208 & n45209;
  assign n45205 = n43804 ^ n43229;
  assign n45206 = n45205 ^ n44543;
  assign n45211 = n45210 ^ n45206;
  assign n45212 = n45178 ^ n45050;
  assign n45213 = n45212 ^ n45206;
  assign n45214 = n45211 & ~n45213;
  assign n45215 = n45214 ^ n45210;
  assign n45217 = n45216 ^ n45215;
  assign n45218 = n43803 ^ n43236;
  assign n45219 = n45218 ^ n44581;
  assign n45220 = n45219 ^ n45216;
  assign n45221 = n45217 & n45220;
  assign n45222 = n45221 ^ n45219;
  assign n45202 = n43755 ^ n43243;
  assign n45203 = n45202 ^ n44607;
  assign n45198 = ~n45009 & n45046;
  assign n45193 = n42862 ^ n42318;
  assign n45194 = n45193 ^ n43893;
  assign n45191 = n44448 ^ n44445;
  assign n45188 = n45005 ^ n45001;
  assign n45189 = ~n45006 & n45188;
  assign n45190 = n45189 ^ n45001;
  assign n45192 = n45191 ^ n45190;
  assign n45195 = n45194 ^ n45192;
  assign n45196 = n45195 ^ n41684;
  assign n45185 = n45007 ^ n44999;
  assign n45186 = ~n45008 & n45185;
  assign n45187 = n45186 ^ n41829;
  assign n45197 = n45196 ^ n45187;
  assign n45199 = n45198 ^ n45197;
  assign n45182 = n45181 ^ n45047;
  assign n45183 = ~n45048 & n45182;
  assign n45184 = n45183 ^ n44800;
  assign n45200 = n45199 ^ n45184;
  assign n44795 = n43044 ^ n34939;
  assign n44796 = n44795 ^ n2345;
  assign n44797 = n44796 ^ n33189;
  assign n45201 = n45200 ^ n44797;
  assign n45204 = n45203 ^ n45201;
  assign n45318 = n45222 ^ n45204;
  assign n45319 = n45318 ^ n42302;
  assign n45327 = n45219 ^ n45217;
  assign n45320 = n45209 ^ n45208;
  assign n45321 = ~n42308 & ~n45320;
  assign n45322 = n45321 ^ n42304;
  assign n45323 = n45212 ^ n45211;
  assign n45324 = n45323 ^ n45321;
  assign n45325 = ~n45322 & ~n45324;
  assign n45326 = n45325 ^ n42304;
  assign n45328 = n45327 ^ n45326;
  assign n45329 = n45327 ^ n42561;
  assign n45330 = n45328 & ~n45329;
  assign n45331 = n45330 ^ n42561;
  assign n45332 = n45331 ^ n45318;
  assign n45333 = n45319 & ~n45332;
  assign n45334 = n45333 ^ n42302;
  assign n45251 = n43951 ^ n42854;
  assign n45252 = n45251 ^ n44623;
  assign n45245 = n43160 ^ n35004;
  assign n45246 = n45245 ^ n39542;
  assign n45247 = n45246 ^ n2432;
  assign n45243 = n45197 & ~n45198;
  assign n45239 = n44453 ^ n44260;
  assign n45240 = n45239 ^ n44451;
  assign n45236 = n42856 ^ n42312;
  assign n45237 = n45236 ^ n43919;
  assign n45233 = n45194 ^ n45191;
  assign n45234 = ~n45192 & n45233;
  assign n45235 = n45234 ^ n45194;
  assign n45238 = n45237 ^ n45235;
  assign n45241 = n45240 ^ n45238;
  assign n45229 = n45195 ^ n45187;
  assign n45230 = ~n45196 & n45229;
  assign n45231 = n45230 ^ n41684;
  assign n45232 = n45231 ^ n41678;
  assign n45242 = n45241 ^ n45232;
  assign n45244 = n45243 ^ n45242;
  assign n45248 = n45247 ^ n45244;
  assign n45226 = n45199 ^ n44797;
  assign n45227 = ~n45200 & n45226;
  assign n45228 = n45227 ^ n44797;
  assign n45249 = n45248 ^ n45228;
  assign n45223 = n45222 ^ n45201;
  assign n45224 = n45204 & n45223;
  assign n45225 = n45224 ^ n45203;
  assign n45250 = n45249 ^ n45225;
  assign n45316 = n45252 ^ n45250;
  assign n45317 = n45316 ^ n42298;
  assign n45405 = n45334 ^ n45317;
  assign n45406 = n45328 ^ n42561;
  assign n45407 = n45323 ^ n45322;
  assign n45408 = ~n45406 & n45407;
  assign n45409 = n45331 ^ n45319;
  assign n45410 = ~n45408 & ~n45409;
  assign n45411 = n45405 & ~n45410;
  assign n45335 = n45334 ^ n45316;
  assign n45336 = n45317 & n45335;
  assign n45337 = n45336 ^ n42298;
  assign n45253 = n45252 ^ n45249;
  assign n45254 = ~n45250 & n45253;
  assign n45255 = n45254 ^ n45252;
  assign n44792 = n43796 ^ n42849;
  assign n44793 = n44792 ^ n44635;
  assign n44791 = n44675 ^ n44674;
  assign n44794 = n44793 ^ n44791;
  assign n45314 = n45255 ^ n44794;
  assign n45315 = n45314 ^ n42292;
  assign n45404 = n45337 ^ n45315;
  assign n45571 = n45411 ^ n45404;
  assign n45539 = n43584 ^ n35061;
  assign n45540 = n45539 ^ n39933;
  assign n45541 = n45540 ^ n33683;
  assign n45538 = n45410 ^ n45405;
  assign n45542 = n45541 ^ n45538;
  assign n45544 = n43589 ^ n35065;
  assign n45545 = n45544 ^ n39911;
  assign n45546 = n45545 ^ n33687;
  assign n45543 = n45409 ^ n45408;
  assign n45547 = n45546 ^ n45543;
  assign n45557 = n43598 ^ n35069;
  assign n45558 = n45557 ^ n39920;
  assign n45559 = n45558 ^ n33696;
  assign n45550 = n43593 ^ n35072;
  assign n45551 = n45550 ^ n39915;
  assign n45552 = n45551 ^ n33691;
  assign n2502 = n2501 ^ n2468;
  assign n2533 = n2532 ^ n2502;
  assign n2543 = n2542 ^ n2533;
  assign n45548 = n45320 ^ n42308;
  assign n45549 = n2543 & n45548;
  assign n45553 = n45552 ^ n45549;
  assign n45554 = n45549 ^ n45407;
  assign n45555 = n45553 & ~n45554;
  assign n45556 = n45555 ^ n45552;
  assign n45560 = n45559 ^ n45556;
  assign n45561 = n45407 ^ n45406;
  assign n45562 = n45561 ^ n45556;
  assign n45563 = n45560 & ~n45562;
  assign n45564 = n45563 ^ n45559;
  assign n45565 = n45564 ^ n45543;
  assign n45566 = n45547 & ~n45565;
  assign n45567 = n45566 ^ n45546;
  assign n45568 = n45567 ^ n45538;
  assign n45569 = n45542 & ~n45568;
  assign n45570 = n45569 ^ n45541;
  assign n45572 = n45571 ^ n45570;
  assign n45573 = n43579 ^ n35056;
  assign n45574 = n45573 ^ n39907;
  assign n45575 = n45574 ^ n33678;
  assign n45576 = n45575 ^ n45571;
  assign n45577 = ~n45572 & n45576;
  assign n45578 = n45577 ^ n45575;
  assign n45338 = n45337 ^ n45314;
  assign n45339 = ~n45315 & ~n45338;
  assign n45340 = n45339 ^ n42292;
  assign n45256 = n45255 ^ n44791;
  assign n45257 = n44794 & n45256;
  assign n45258 = n45257 ^ n44793;
  assign n44788 = n43792 ^ n42844;
  assign n44789 = n44788 ^ n44731;
  assign n44786 = n44679 ^ n44593;
  assign n44787 = n44786 ^ n44676;
  assign n44790 = n44789 ^ n44787;
  assign n45312 = n45258 ^ n44790;
  assign n45313 = n45312 ^ n42577;
  assign n45413 = n45340 ^ n45313;
  assign n45412 = ~n45404 & ~n45411;
  assign n45533 = n45413 ^ n45412;
  assign n45537 = n45536 ^ n45533;
  assign n45706 = n45578 ^ n45537;
  assign n45709 = n45708 ^ n45706;
  assign n45711 = n44765 ^ n43779;
  assign n44750 = n44722 ^ n44646;
  assign n45712 = n45711 ^ n44750;
  assign n45710 = n45575 ^ n45572;
  assign n45713 = n45712 ^ n45710;
  assign n45715 = n44771 ^ n43783;
  assign n44755 = n44719 ^ n44716;
  assign n45716 = n45715 ^ n44755;
  assign n45714 = n45567 ^ n45542;
  assign n45717 = n45716 ^ n45714;
  assign n45719 = n44844 ^ n43787;
  assign n44760 = n44711 ^ n44651;
  assign n45720 = n45719 ^ n44760;
  assign n45718 = n45564 ^ n45547;
  assign n45721 = n45720 ^ n45718;
  assign n45724 = n44776 ^ n43790;
  assign n44768 = n44708 ^ n44705;
  assign n45725 = n45724 ^ n44768;
  assign n45722 = n45561 ^ n45559;
  assign n45723 = n45722 ^ n45556;
  assign n45726 = n45725 ^ n45723;
  assign n45729 = n45552 ^ n45407;
  assign n45730 = n45729 ^ n45549;
  assign n45727 = n44781 ^ n43792;
  assign n44773 = n44700 ^ n44656;
  assign n45728 = n45727 ^ n44773;
  assign n45731 = n45730 ^ n45728;
  assign n45817 = n43815 ^ n42862;
  assign n45818 = n45817 ^ n44485;
  assign n45686 = n45164 ^ n45057;
  assign n45819 = n45818 ^ n45686;
  assign n45779 = n45161 ^ n45158;
  assign n45776 = n43919 ^ n43208;
  assign n45777 = n45776 ^ n44490;
  assign n45813 = n45779 ^ n45777;
  assign n45739 = n43893 ^ n43161;
  assign n45740 = n45739 ^ n44501;
  assign n45738 = n45153 ^ n45062;
  assign n45741 = n45740 ^ n45738;
  assign n45743 = n43865 ^ n43176;
  assign n45744 = n45743 ^ n44498;
  assign n45742 = n45150 ^ n45147;
  assign n45745 = n45744 ^ n45742;
  assign n45747 = n43840 ^ n43172;
  assign n45748 = n45747 ^ n45240;
  assign n45746 = n45142 ^ n45067;
  assign n45749 = n45748 ^ n45746;
  assign n45751 = n45191 ^ n43167;
  assign n45752 = n45751 ^ n43745;
  assign n45750 = n45139 ^ n45072;
  assign n45753 = n45752 ^ n45750;
  assign n45756 = n45136 ^ n45133;
  assign n45754 = n45005 ^ n44517;
  assign n45755 = n45754 ^ n43913;
  assign n45757 = n45756 ^ n45755;
  assign n45677 = n44474 ^ n43763;
  assign n45678 = n45677 ^ n44910;
  assign n45676 = n45128 ^ n45125;
  assign n45679 = n45678 ^ n45676;
  assign n45652 = n44903 ^ n43767;
  assign n45653 = n45652 ^ n44184;
  assign n45651 = n45120 ^ n45117;
  assign n45654 = n45653 ^ n45651;
  assign n45472 = n44033 ^ n43832;
  assign n45473 = n45472 ^ n44896;
  assign n45470 = n45112 ^ n45076;
  assign n45471 = n45470 ^ n45073;
  assign n45474 = n45473 ^ n45471;
  assign n45396 = n45103 ^ n45092;
  assign n45300 = n43769 ^ n43439;
  assign n45301 = n45300 ^ n44814;
  assign n45299 = n45100 ^ n45097;
  assign n45302 = n45301 ^ n45299;
  assign n44747 = n44006 ^ n43314;
  assign n44748 = n44747 ^ n44746;
  assign n44749 = n44748 ^ n44745;
  assign n44751 = n43773 ^ n43307;
  assign n44753 = n44752 ^ n44751;
  assign n44754 = n44753 ^ n44750;
  assign n44756 = n43996 ^ n42834;
  assign n44758 = n44757 ^ n44756;
  assign n44759 = n44758 ^ n44755;
  assign n44761 = n43989 ^ n43297;
  assign n44763 = n44762 ^ n44761;
  assign n44764 = n44763 ^ n44760;
  assign n44766 = n44765 ^ n43290;
  assign n44767 = n44766 ^ n43775;
  assign n44769 = n44768 ^ n44767;
  assign n44770 = n43979 ^ n42836;
  assign n44772 = n44771 ^ n44770;
  assign n44774 = n44773 ^ n44772;
  assign n45274 = n44697 ^ n44694;
  assign n44778 = n44689 ^ n44661;
  assign n44775 = n43783 ^ n43271;
  assign n44777 = n44776 ^ n44775;
  assign n44779 = n44778 ^ n44777;
  assign n44783 = n44686 ^ n44666;
  assign n44780 = n43787 ^ n42838;
  assign n44782 = n44781 ^ n44780;
  assign n44784 = n44783 ^ n44782;
  assign n45259 = n45258 ^ n44787;
  assign n45260 = ~n44790 & ~n45259;
  assign n45261 = n45260 ^ n44789;
  assign n44785 = n44683 ^ n44671;
  assign n45262 = n45261 ^ n44785;
  assign n45263 = n43790 ^ n42839;
  assign n45264 = n45263 ^ n44825;
  assign n45265 = n45264 ^ n44785;
  assign n45266 = ~n45262 & ~n45265;
  assign n45267 = n45266 ^ n45264;
  assign n45268 = n45267 ^ n44783;
  assign n45269 = ~n44784 & ~n45268;
  assign n45270 = n45269 ^ n44782;
  assign n45271 = n45270 ^ n44777;
  assign n45272 = ~n44779 & ~n45271;
  assign n45273 = n45272 ^ n44778;
  assign n45275 = n45274 ^ n45273;
  assign n45276 = n43779 ^ n42837;
  assign n45277 = n45276 ^ n44844;
  assign n45278 = n45277 ^ n45274;
  assign n45279 = ~n45275 & ~n45278;
  assign n45280 = n45279 ^ n45277;
  assign n45281 = n45280 ^ n44773;
  assign n45282 = ~n44774 & ~n45281;
  assign n45283 = n45282 ^ n44772;
  assign n45284 = n45283 ^ n44768;
  assign n45285 = ~n44769 & ~n45284;
  assign n45286 = n45285 ^ n44767;
  assign n45287 = n45286 ^ n44760;
  assign n45288 = ~n44764 & n45287;
  assign n45289 = n45288 ^ n44763;
  assign n45290 = n45289 ^ n44758;
  assign n45291 = n44759 & ~n45290;
  assign n45292 = n45291 ^ n44755;
  assign n45293 = n45292 ^ n44753;
  assign n45294 = n44754 & n45293;
  assign n45295 = n45294 ^ n44750;
  assign n45296 = n45295 ^ n44745;
  assign n45297 = ~n44749 & ~n45296;
  assign n45298 = n45297 ^ n44748;
  assign n45393 = n45299 ^ n45298;
  assign n45394 = ~n45302 & ~n45393;
  assign n45395 = n45394 ^ n45301;
  assign n45397 = n45396 ^ n45395;
  assign n45391 = n43761 ^ n43498;
  assign n45392 = n45391 ^ n44811;
  assign n45442 = n45396 ^ n45392;
  assign n45443 = n45397 & ~n45442;
  assign n45444 = n45443 ^ n45392;
  assign n45441 = n45106 ^ n45087;
  assign n45445 = n45444 ^ n45441;
  assign n45439 = n44019 ^ n43715;
  assign n45440 = n45439 ^ n44807;
  assign n45456 = n45441 ^ n45440;
  assign n45457 = n45445 & n45456;
  assign n45458 = n45457 ^ n45440;
  assign n45455 = n45109 ^ n45082;
  assign n45459 = n45458 ^ n45455;
  assign n45453 = n44803 ^ n44026;
  assign n45454 = n45453 ^ n43737;
  assign n45467 = n45455 ^ n45454;
  assign n45468 = n45459 & n45467;
  assign n45469 = n45468 ^ n45454;
  assign n45648 = n45471 ^ n45469;
  assign n45649 = n45474 & n45648;
  assign n45650 = n45649 ^ n45473;
  assign n45673 = n45651 ^ n45650;
  assign n45674 = n45654 & ~n45673;
  assign n45675 = n45674 ^ n45653;
  assign n45758 = n45676 ^ n45675;
  assign n45759 = ~n45679 & n45758;
  assign n45760 = n45759 ^ n45678;
  assign n45761 = n45760 ^ n45755;
  assign n45762 = n45757 & ~n45761;
  assign n45763 = n45762 ^ n45756;
  assign n45764 = n45763 ^ n45750;
  assign n45765 = ~n45753 & ~n45764;
  assign n45766 = n45765 ^ n45752;
  assign n45767 = n45766 ^ n45746;
  assign n45768 = ~n45749 & n45767;
  assign n45769 = n45768 ^ n45748;
  assign n45770 = n45769 ^ n45742;
  assign n45771 = ~n45745 & ~n45770;
  assign n45772 = n45771 ^ n45744;
  assign n45773 = n45772 ^ n45738;
  assign n45774 = n45741 & ~n45773;
  assign n45775 = n45774 ^ n45740;
  assign n45814 = n45779 ^ n45775;
  assign n45815 = ~n45813 & n45814;
  assign n45816 = n45815 ^ n45777;
  assign n45905 = n45816 ^ n45686;
  assign n45906 = ~n45819 & n45905;
  assign n45907 = n45906 ^ n45818;
  assign n45908 = n45907 ^ n43809;
  assign n45902 = n45167 ^ n45052;
  assign n45903 = n45902 ^ n45236;
  assign n45820 = n45819 ^ n45816;
  assign n45821 = n45820 ^ n42318;
  assign n45778 = n45777 ^ n45775;
  assign n45780 = n45779 ^ n45778;
  assign n45781 = n45780 ^ n42542;
  assign n45782 = n45772 ^ n45741;
  assign n45783 = n45782 ^ n42495;
  assign n45784 = n45769 ^ n45745;
  assign n45785 = n45784 ^ n42508;
  assign n45786 = n45766 ^ n45749;
  assign n45787 = n45786 ^ n42504;
  assign n45796 = n45763 ^ n45753;
  assign n45791 = n45760 ^ n45757;
  assign n45680 = n45679 ^ n45675;
  assign n45655 = n45654 ^ n45650;
  assign n45475 = n45474 ^ n45469;
  assign n45460 = n45459 ^ n45454;
  assign n45461 = n45460 ^ n42935;
  assign n45446 = n45445 ^ n45440;
  assign n45447 = n45446 ^ n42290;
  assign n45398 = n45397 ^ n45392;
  assign n45435 = n45398 ^ n42866;
  assign n45303 = n45302 ^ n45298;
  assign n45304 = n45303 ^ n42870;
  assign n45382 = n45295 ^ n44749;
  assign n45305 = n45292 ^ n44754;
  assign n45306 = n45305 ^ n42875;
  assign n45307 = n45286 ^ n44764;
  assign n45308 = n45307 ^ n42900;
  assign n45366 = n45283 ^ n44769;
  assign n45361 = n45280 ^ n44774;
  assign n45356 = n45277 ^ n45275;
  assign n45347 = n45267 ^ n44784;
  assign n45310 = n45264 ^ n45262;
  assign n45311 = n45310 ^ n42584;
  assign n45341 = n45340 ^ n45312;
  assign n45342 = ~n45313 & n45341;
  assign n45343 = n45342 ^ n42577;
  assign n45344 = n45343 ^ n45310;
  assign n45345 = ~n45311 & ~n45344;
  assign n45346 = n45345 ^ n42584;
  assign n45348 = n45347 ^ n45346;
  assign n45349 = n45347 ^ n42665;
  assign n45350 = ~n45348 & n45349;
  assign n45351 = n45350 ^ n42665;
  assign n45309 = n45270 ^ n44779;
  assign n45352 = n45351 ^ n45309;
  assign n45353 = n45351 ^ n42821;
  assign n45354 = n45352 & n45353;
  assign n45355 = n45354 ^ n42821;
  assign n45357 = n45356 ^ n45355;
  assign n45358 = n45356 ^ n42850;
  assign n45359 = ~n45357 & ~n45358;
  assign n45360 = n45359 ^ n42850;
  assign n45362 = n45361 ^ n45360;
  assign n45363 = n45361 ^ n42845;
  assign n45364 = ~n45362 & n45363;
  assign n45365 = n45364 ^ n42845;
  assign n45367 = n45366 ^ n45365;
  assign n45368 = n45366 ^ n42840;
  assign n45369 = n45367 & ~n45368;
  assign n45370 = n45369 ^ n42840;
  assign n45371 = n45370 ^ n45307;
  assign n45372 = n45308 & ~n45371;
  assign n45373 = n45372 ^ n42900;
  assign n45374 = n45373 ^ n42907;
  assign n45375 = n45289 ^ n44759;
  assign n45376 = n45375 ^ n45373;
  assign n45377 = ~n45374 & n45376;
  assign n45378 = n45377 ^ n42907;
  assign n45379 = n45378 ^ n45305;
  assign n45380 = n45306 & ~n45379;
  assign n45381 = n45380 ^ n42875;
  assign n45383 = n45382 ^ n45381;
  assign n45384 = n45382 ^ n42874;
  assign n45385 = ~n45383 & ~n45384;
  assign n45386 = n45385 ^ n42874;
  assign n45387 = n45386 ^ n45303;
  assign n45388 = ~n45304 & ~n45387;
  assign n45389 = n45388 ^ n42870;
  assign n45436 = n45398 ^ n45389;
  assign n45437 = n45435 & ~n45436;
  assign n45438 = n45437 ^ n42866;
  assign n45450 = n45446 ^ n45438;
  assign n45451 = n45447 & n45450;
  assign n45452 = n45451 ^ n42290;
  assign n45464 = n45460 ^ n45452;
  assign n45465 = ~n45461 & n45464;
  assign n45466 = n45465 ^ n42935;
  assign n45476 = n45475 ^ n45466;
  assign n45645 = n45475 ^ n42286;
  assign n45646 = ~n45476 & n45645;
  assign n45647 = n45646 ^ n42286;
  assign n45656 = n45655 ^ n45647;
  assign n45670 = n45655 ^ n43008;
  assign n45671 = n45656 & ~n45670;
  assign n45672 = n45671 ^ n43008;
  assign n45681 = n45680 ^ n45672;
  assign n45788 = n45680 ^ n43148;
  assign n45789 = ~n45681 & n45788;
  assign n45790 = n45789 ^ n43148;
  assign n45792 = n45791 ^ n45790;
  assign n45793 = n45791 ^ n43196;
  assign n45794 = n45792 & ~n45793;
  assign n45795 = n45794 ^ n43196;
  assign n45797 = n45796 ^ n45795;
  assign n45798 = n45796 ^ n42501;
  assign n45799 = ~n45797 & ~n45798;
  assign n45800 = n45799 ^ n42501;
  assign n45801 = n45800 ^ n45786;
  assign n45802 = ~n45787 & ~n45801;
  assign n45803 = n45802 ^ n42504;
  assign n45804 = n45803 ^ n45784;
  assign n45805 = n45785 & n45804;
  assign n45806 = n45805 ^ n42508;
  assign n45807 = n45806 ^ n45782;
  assign n45808 = ~n45783 & ~n45807;
  assign n45809 = n45808 ^ n42495;
  assign n45810 = n45809 ^ n45780;
  assign n45811 = ~n45781 & ~n45810;
  assign n45812 = n45811 ^ n42542;
  assign n45898 = n45820 ^ n45812;
  assign n45899 = ~n45821 & n45898;
  assign n45900 = n45899 ^ n42318;
  assign n45901 = n45900 ^ n44532;
  assign n45904 = n45903 ^ n45901;
  assign n45909 = n45908 ^ n45904;
  assign n45822 = n45821 ^ n45812;
  assign n45823 = n45809 ^ n45781;
  assign n45824 = n45803 ^ n45785;
  assign n45682 = n45681 ^ n43148;
  assign n45390 = n45389 ^ n42866;
  assign n45399 = n45398 ^ n45390;
  assign n45400 = n45375 ^ n45374;
  assign n45401 = n45367 ^ n42840;
  assign n45402 = n45362 ^ n42845;
  assign n45403 = n45343 ^ n45311;
  assign n45414 = ~n45412 & ~n45413;
  assign n45415 = ~n45403 & n45414;
  assign n45416 = n45348 ^ n42665;
  assign n45417 = n45415 & ~n45416;
  assign n45418 = n45352 ^ n42821;
  assign n45419 = ~n45417 & ~n45418;
  assign n45420 = n45357 ^ n42850;
  assign n45421 = n45419 & ~n45420;
  assign n45422 = ~n45402 & n45421;
  assign n45423 = n45401 & n45422;
  assign n45424 = n45370 ^ n45308;
  assign n45425 = n45423 & ~n45424;
  assign n45426 = n45400 & ~n45425;
  assign n45427 = n45378 ^ n45306;
  assign n45428 = n45426 & ~n45427;
  assign n45429 = n45383 ^ n42874;
  assign n45430 = ~n45428 & ~n45429;
  assign n45431 = n45386 ^ n42870;
  assign n45432 = n45431 ^ n45303;
  assign n45433 = ~n45430 & ~n45432;
  assign n45434 = n45399 & ~n45433;
  assign n45448 = n45447 ^ n45438;
  assign n45449 = n45434 & n45448;
  assign n45462 = n45461 ^ n45452;
  assign n45463 = n45449 & n45462;
  assign n45477 = n45476 ^ n42286;
  assign n45644 = ~n45463 & n45477;
  assign n45657 = n45656 ^ n43008;
  assign n45683 = n45644 & ~n45657;
  assign n45825 = ~n45682 & ~n45683;
  assign n45826 = n45792 ^ n43196;
  assign n45827 = n45825 & n45826;
  assign n45828 = n45797 ^ n42501;
  assign n45829 = ~n45827 & ~n45828;
  assign n45830 = n45800 ^ n45787;
  assign n45831 = ~n45829 & ~n45830;
  assign n45832 = n45824 & ~n45831;
  assign n45833 = n45806 ^ n45783;
  assign n45834 = ~n45832 & ~n45833;
  assign n45835 = n45823 & n45834;
  assign n45896 = n45822 & ~n45835;
  assign n45893 = n43877 ^ n35583;
  assign n45894 = n45893 ^ n40231;
  assign n45895 = n45894 ^ n2524;
  assign n45897 = n45896 ^ n45895;
  assign n45910 = n45909 ^ n45897;
  assign n45836 = n45835 ^ n45822;
  assign n45735 = n43849 ^ n2397;
  assign n45736 = n45735 ^ n40235;
  assign n45737 = n45736 ^ n34132;
  assign n45837 = n45836 ^ n45737;
  assign n45841 = n45834 ^ n45823;
  assign n45838 = n35590 ^ n1408;
  assign n45839 = n45838 ^ n40241;
  assign n45840 = n45839 ^ n34136;
  assign n45842 = n45841 ^ n45840;
  assign n45846 = n45833 ^ n45832;
  assign n45843 = n35595 ^ n1390;
  assign n45844 = n45843 ^ n40282;
  assign n45845 = n45844 ^ n34142;
  assign n45847 = n45846 ^ n45845;
  assign n45851 = n45831 ^ n45824;
  assign n45848 = n43725 ^ n1289;
  assign n45849 = n45848 ^ n40245;
  assign n45850 = n45849 ^ n34147;
  assign n45852 = n45851 ^ n45850;
  assign n45854 = n43509 ^ n1274;
  assign n45855 = n45854 ^ n40271;
  assign n45856 = n45855 ^ n34221;
  assign n45853 = n45830 ^ n45829;
  assign n45857 = n45856 ^ n45853;
  assign n45861 = n45828 ^ n45827;
  assign n45862 = n45861 ^ n45860;
  assign n45864 = n43519 ^ n35609;
  assign n45865 = n45864 ^ n40260;
  assign n45866 = n45865 ^ n905;
  assign n45863 = n45826 ^ n45825;
  assign n45867 = n45866 ^ n45863;
  assign n45684 = n45683 ^ n45682;
  assign n45666 = n43694 ^ n35613;
  assign n45667 = n45666 ^ n809;
  assign n45668 = n45667 ^ n34174;
  assign n45868 = n45684 ^ n45668;
  assign n45658 = n45657 ^ n45644;
  assign n45479 = n43529 ^ n707;
  assign n45480 = n45479 ^ n39999;
  assign n45481 = n45480 ^ n34154;
  assign n45478 = n45477 ^ n45463;
  assign n45482 = n45481 ^ n45478;
  assign n45633 = n45462 ^ n45449;
  assign n45484 = n43539 ^ n35631;
  assign n45485 = n45484 ^ n39988;
  assign n45486 = n45485 ^ n34159;
  assign n45483 = n45448 ^ n45434;
  assign n45487 = n45486 ^ n45483;
  assign n45489 = n43674 ^ n35636;
  assign n45490 = n45489 ^ n39853;
  assign n45491 = n45490 ^ n33775;
  assign n45488 = n45433 ^ n45399;
  assign n45492 = n45491 ^ n45488;
  assign n45496 = n45432 ^ n45430;
  assign n45493 = n43666 ^ n35641;
  assign n45494 = n45493 ^ n39857;
  assign n45495 = n45494 ^ n33634;
  assign n45497 = n45496 ^ n45495;
  assign n45498 = n45429 ^ n45428;
  assign n45502 = n45501 ^ n45498;
  assign n45613 = n43549 ^ n35650;
  assign n45614 = n45613 ^ n39868;
  assign n45615 = n45614 ^ n33644;
  assign n45504 = n43554 ^ n35656;
  assign n45505 = n45504 ^ n39873;
  assign n45506 = n45505 ^ n33737;
  assign n45503 = n45425 ^ n45400;
  assign n45507 = n45506 ^ n45503;
  assign n45509 = n43564 ^ n35666;
  assign n45510 = n45509 ^ n2021;
  assign n45511 = n45510 ^ n33656;
  assign n45508 = n45422 ^ n45401;
  assign n45512 = n45511 ^ n45508;
  assign n45516 = n45421 ^ n45402;
  assign n45513 = n43643 ^ n35671;
  assign n45514 = n45513 ^ n39879;
  assign n45515 = n45514 ^ n2013;
  assign n45517 = n45516 ^ n45515;
  assign n45591 = n45420 ^ n45419;
  assign n45521 = n45418 ^ n45417;
  assign n45518 = n43568 ^ n35677;
  assign n45519 = n45518 ^ n39886;
  assign n45520 = n45519 ^ n1873;
  assign n45522 = n45521 ^ n45520;
  assign n45526 = n45416 ^ n45415;
  assign n45527 = n45526 ^ n45525;
  assign n45531 = n45414 ^ n45403;
  assign n45528 = n43574 ^ n35684;
  assign n45529 = n45528 ^ n39897;
  assign n45530 = n45529 ^ n33667;
  assign n45532 = n45531 ^ n45530;
  assign n45579 = n45578 ^ n45536;
  assign n45580 = ~n45537 & ~n45579;
  assign n45581 = n45580 ^ n45533;
  assign n45582 = n45581 ^ n45530;
  assign n45583 = n45532 & n45582;
  assign n45584 = n45583 ^ n45531;
  assign n45585 = n45584 ^ n45526;
  assign n45586 = n45527 & ~n45585;
  assign n45587 = n45586 ^ n45525;
  assign n45588 = n45587 ^ n45521;
  assign n45589 = n45522 & ~n45588;
  assign n45590 = n45589 ^ n45520;
  assign n45592 = n45591 ^ n45590;
  assign n1848 = n1847 ^ n1811;
  assign n1882 = n1881 ^ n1848;
  assign n1892 = n1891 ^ n1882;
  assign n45593 = n45590 ^ n1892;
  assign n45594 = n45592 & n45593;
  assign n45595 = n45594 ^ n1892;
  assign n45596 = n45595 ^ n45515;
  assign n45597 = ~n45517 & ~n45596;
  assign n45598 = n45597 ^ n45516;
  assign n45599 = n45598 ^ n45511;
  assign n45600 = n45512 & n45599;
  assign n45601 = n45600 ^ n45508;
  assign n45605 = n45604 ^ n45601;
  assign n45606 = n45424 ^ n45423;
  assign n45607 = n45606 ^ n45601;
  assign n45608 = n45605 & n45607;
  assign n45609 = n45608 ^ n45604;
  assign n45610 = n45609 ^ n45503;
  assign n45611 = n45507 & ~n45610;
  assign n45612 = n45611 ^ n45506;
  assign n45616 = n45615 ^ n45612;
  assign n45617 = n45427 ^ n45426;
  assign n45618 = n45617 ^ n45612;
  assign n45619 = n45616 & ~n45618;
  assign n45620 = n45619 ^ n45615;
  assign n45621 = n45620 ^ n45498;
  assign n45622 = n45502 & ~n45621;
  assign n45623 = n45622 ^ n45501;
  assign n45624 = n45623 ^ n45495;
  assign n45625 = ~n45497 & ~n45624;
  assign n45626 = n45625 ^ n45496;
  assign n45627 = n45626 ^ n45488;
  assign n45628 = ~n45492 & ~n45627;
  assign n45629 = n45628 ^ n45491;
  assign n45630 = n45629 ^ n45483;
  assign n45631 = n45487 & ~n45630;
  assign n45632 = n45631 ^ n45486;
  assign n45634 = n45633 ^ n45632;
  assign n45635 = n43533 ^ n35625;
  assign n45636 = n45635 ^ n39848;
  assign n45637 = n45636 ^ n34167;
  assign n45638 = n45637 ^ n45633;
  assign n45639 = ~n45634 & n45638;
  assign n45640 = n45639 ^ n45637;
  assign n45641 = n45640 ^ n45478;
  assign n45642 = n45482 & ~n45641;
  assign n45643 = n45642 ^ n45481;
  assign n45659 = n45658 ^ n45643;
  assign n45660 = n43524 ^ n35619;
  assign n45661 = n45660 ^ n39843;
  assign n45662 = n45661 ^ n801;
  assign n45663 = n45662 ^ n45658;
  assign n45664 = ~n45659 & n45663;
  assign n45665 = n45664 ^ n45662;
  assign n45869 = n45684 ^ n45665;
  assign n45870 = n45868 & ~n45869;
  assign n45871 = n45870 ^ n45668;
  assign n45872 = n45871 ^ n45863;
  assign n45873 = n45867 & ~n45872;
  assign n45874 = n45873 ^ n45866;
  assign n45875 = n45874 ^ n45861;
  assign n45876 = ~n45862 & n45875;
  assign n45877 = n45876 ^ n45860;
  assign n45878 = n45877 ^ n45853;
  assign n45879 = n45857 & ~n45878;
  assign n45880 = n45879 ^ n45856;
  assign n45881 = n45880 ^ n45850;
  assign n45882 = n45852 & ~n45881;
  assign n45883 = n45882 ^ n45851;
  assign n45884 = n45883 ^ n45845;
  assign n45885 = n45847 & ~n45884;
  assign n45886 = n45885 ^ n45846;
  assign n45887 = n45886 ^ n45841;
  assign n45888 = n45842 & ~n45887;
  assign n45889 = n45888 ^ n45840;
  assign n45890 = n45889 ^ n45836;
  assign n45891 = n45837 & ~n45890;
  assign n45892 = n45891 ^ n45737;
  assign n45911 = n45910 ^ n45892;
  assign n45733 = n44731 ^ n43951;
  assign n45734 = n45733 ^ n44778;
  assign n45912 = n45911 ^ n45734;
  assign n45931 = n45889 ^ n45837;
  assign n45914 = n44623 ^ n43803;
  assign n45915 = n45914 ^ n44785;
  assign n45913 = n45886 ^ n45842;
  assign n45916 = n45915 ^ n45913;
  assign n45919 = n44581 ^ n43932;
  assign n45920 = n45919 ^ n44791;
  assign n45921 = n45880 ^ n45852;
  assign n45922 = ~n45920 & n45921;
  assign n45917 = n44607 ^ n43804;
  assign n45918 = n45917 ^ n44787;
  assign n45923 = n45922 ^ n45918;
  assign n45924 = n45883 ^ n45847;
  assign n45925 = n45924 ^ n45918;
  assign n45926 = ~n45923 & n45925;
  assign n45927 = n45926 ^ n45922;
  assign n45928 = n45927 ^ n45913;
  assign n45929 = n45916 & ~n45928;
  assign n45930 = n45929 ^ n45915;
  assign n45932 = n45931 ^ n45930;
  assign n45933 = n44635 ^ n43755;
  assign n45934 = n45933 ^ n44783;
  assign n45935 = n45934 ^ n45931;
  assign n45936 = ~n45932 & n45935;
  assign n45937 = n45936 ^ n45934;
  assign n45938 = n45937 ^ n45734;
  assign n45939 = n45912 & n45938;
  assign n45940 = n45939 ^ n45911;
  assign n45732 = n45548 ^ n2543;
  assign n45941 = n45940 ^ n45732;
  assign n45942 = n44825 ^ n43796;
  assign n45943 = n45942 ^ n45274;
  assign n45944 = n45943 ^ n45732;
  assign n45945 = n45941 & ~n45944;
  assign n45946 = n45945 ^ n45943;
  assign n45947 = n45946 ^ n45728;
  assign n45948 = ~n45731 & ~n45947;
  assign n45949 = n45948 ^ n45730;
  assign n45950 = n45949 ^ n45723;
  assign n45951 = ~n45726 & ~n45950;
  assign n45952 = n45951 ^ n45725;
  assign n45953 = n45952 ^ n45718;
  assign n45954 = n45721 & n45953;
  assign n45955 = n45954 ^ n45720;
  assign n45956 = n45955 ^ n45716;
  assign n45957 = n45717 & ~n45956;
  assign n45958 = n45957 ^ n45714;
  assign n45959 = n45958 ^ n45710;
  assign n45960 = n45713 & ~n45959;
  assign n45961 = n45960 ^ n45712;
  assign n45962 = n45961 ^ n45706;
  assign n45963 = ~n45709 & n45962;
  assign n45964 = n45963 ^ n45708;
  assign n45704 = n45581 ^ n45532;
  assign n45702 = n44757 ^ n43775;
  assign n45703 = n45702 ^ n45299;
  assign n45705 = n45704 ^ n45703;
  assign n46048 = n45964 ^ n45705;
  assign n46079 = n46048 ^ n43290;
  assign n45988 = n45961 ^ n45708;
  assign n45989 = n45988 ^ n45706;
  assign n45990 = n45989 ^ n42836;
  assign n45991 = n45958 ^ n45712;
  assign n45992 = n45991 ^ n45710;
  assign n45993 = n45992 ^ n42837;
  assign n46036 = n45955 ^ n45717;
  assign n45994 = n45952 ^ n45721;
  assign n45995 = n45994 ^ n42838;
  assign n45996 = n45949 ^ n45726;
  assign n45997 = n45996 ^ n42839;
  assign n45998 = n45943 ^ n45941;
  assign n45999 = n45998 ^ n42849;
  assign n46013 = n45934 ^ n45932;
  assign n46001 = n45927 ^ n45916;
  assign n46002 = n46001 ^ n43236;
  assign n46003 = n45921 ^ n45920;
  assign n46004 = n43222 & ~n46003;
  assign n46005 = n46004 ^ n43229;
  assign n46006 = n45924 ^ n45923;
  assign n46007 = n46006 ^ n46004;
  assign n46008 = n46005 & n46007;
  assign n46009 = n46008 ^ n43229;
  assign n46010 = n46009 ^ n46001;
  assign n46011 = ~n46002 & ~n46010;
  assign n46012 = n46011 ^ n43236;
  assign n46014 = n46013 ^ n46012;
  assign n46015 = n46013 ^ n43243;
  assign n46016 = n46014 & ~n46015;
  assign n46017 = n46016 ^ n43243;
  assign n46000 = n45937 ^ n45912;
  assign n46018 = n46017 ^ n46000;
  assign n46019 = n46017 ^ n42854;
  assign n46020 = n46018 & ~n46019;
  assign n46021 = n46020 ^ n42854;
  assign n46022 = n46021 ^ n45998;
  assign n46023 = n45999 & ~n46022;
  assign n46024 = n46023 ^ n42849;
  assign n46025 = n46024 ^ n42844;
  assign n46026 = n45946 ^ n45731;
  assign n46027 = n46026 ^ n46024;
  assign n46028 = n46025 & ~n46027;
  assign n46029 = n46028 ^ n42844;
  assign n46030 = n46029 ^ n45996;
  assign n46031 = n45997 & n46030;
  assign n46032 = n46031 ^ n42839;
  assign n46033 = n46032 ^ n45994;
  assign n46034 = n45995 & ~n46033;
  assign n46035 = n46034 ^ n42838;
  assign n46037 = n46036 ^ n46035;
  assign n46038 = n46036 ^ n43271;
  assign n46039 = n46037 & n46038;
  assign n46040 = n46039 ^ n43271;
  assign n46041 = n46040 ^ n45992;
  assign n46042 = ~n45993 & ~n46041;
  assign n46043 = n46042 ^ n42837;
  assign n46044 = n46043 ^ n45989;
  assign n46045 = n45990 & ~n46044;
  assign n46046 = n46045 ^ n42836;
  assign n46080 = n46079 ^ n46046;
  assign n46081 = n46043 ^ n45990;
  assign n46082 = n46009 ^ n46002;
  assign n46083 = n46006 ^ n46005;
  assign n46084 = n46082 & n46083;
  assign n46085 = n46014 ^ n43243;
  assign n46086 = ~n46084 & n46085;
  assign n46087 = n46018 ^ n42854;
  assign n46088 = ~n46086 & n46087;
  assign n46089 = n46021 ^ n45999;
  assign n46090 = ~n46088 & n46089;
  assign n46091 = n46026 ^ n42844;
  assign n46092 = n46091 ^ n46024;
  assign n46093 = ~n46090 & ~n46092;
  assign n46094 = n46029 ^ n42839;
  assign n46095 = n46094 ^ n45996;
  assign n46096 = n46093 & ~n46095;
  assign n46097 = n46032 ^ n45995;
  assign n46098 = n46096 & n46097;
  assign n46099 = n46037 ^ n43271;
  assign n46100 = ~n46098 & ~n46099;
  assign n46101 = n46040 ^ n45993;
  assign n46102 = n46100 & ~n46101;
  assign n46103 = ~n46081 & n46102;
  assign n46104 = ~n46080 & n46103;
  assign n46047 = n46046 ^ n43290;
  assign n46049 = n46048 ^ n46046;
  assign n46050 = ~n46047 & n46049;
  assign n46051 = n46050 ^ n43290;
  assign n46077 = n46051 ^ n43297;
  assign n45965 = n45964 ^ n45704;
  assign n45966 = n45705 & n45965;
  assign n45967 = n45966 ^ n45703;
  assign n45700 = n45584 ^ n45527;
  assign n45698 = n44752 ^ n43989;
  assign n45699 = n45698 ^ n45396;
  assign n45701 = n45700 ^ n45699;
  assign n45986 = n45967 ^ n45701;
  assign n46078 = n46077 ^ n45986;
  assign n46127 = n46104 ^ n46078;
  assign n46131 = n46130 ^ n46127;
  assign n46132 = n46103 ^ n46080;
  assign n2113 = n2103 ^ n2055;
  assign n2141 = n2140 ^ n2113;
  assign n2148 = n2147 ^ n2141;
  assign n46133 = n46132 ^ n2148;
  assign n46135 = n44320 ^ n1975;
  assign n46136 = n46135 ^ n40529;
  assign n46137 = n46136 ^ n2132;
  assign n46134 = n46102 ^ n46081;
  assign n46138 = n46137 ^ n46134;
  assign n46140 = n44390 ^ n1957;
  assign n46141 = n46140 ^ n40534;
  assign n46142 = n46141 ^ n34732;
  assign n46139 = n46101 ^ n46100;
  assign n46143 = n46142 ^ n46139;
  assign n46147 = n46099 ^ n46098;
  assign n46144 = n44382 ^ n35963;
  assign n46145 = n46144 ^ n40600;
  assign n46146 = n46145 ^ n34737;
  assign n46148 = n46147 ^ n46146;
  assign n46152 = n46097 ^ n46096;
  assign n46149 = n44374 ^ n35969;
  assign n46150 = n46149 ^ n40538;
  assign n46151 = n46150 ^ n34742;
  assign n46153 = n46152 ^ n46151;
  assign n46157 = n46095 ^ n46093;
  assign n46154 = n44325 ^ n35974;
  assign n46155 = n46154 ^ n40544;
  assign n46156 = n46155 ^ n34746;
  assign n46158 = n46157 ^ n46156;
  assign n46160 = n44363 ^ n35979;
  assign n46161 = n46160 ^ n40548;
  assign n46162 = n46161 ^ n1592;
  assign n46159 = n46092 ^ n46090;
  assign n46163 = n46162 ^ n46159;
  assign n46167 = n46089 ^ n46088;
  assign n46164 = n44330 ^ n35984;
  assign n46165 = n46164 ^ n40553;
  assign n46166 = n46165 ^ n34753;
  assign n46168 = n46167 ^ n46166;
  assign n46197 = n46087 ^ n46086;
  assign n46189 = n46085 ^ n46084;
  assign n46170 = n44345 ^ n35999;
  assign n46171 = n46170 ^ n40562;
  assign n46172 = n46171 ^ n34772;
  assign n46169 = n46083 ^ n46082;
  assign n46173 = n46172 ^ n46169;
  assign n46179 = n40565 ^ n2620;
  assign n46180 = n46179 ^ n43752;
  assign n46181 = n46180 ^ n34767;
  assign n46174 = n44520 ^ n2602;
  assign n46175 = n46174 ^ n40771;
  assign n46176 = n46175 ^ n35028;
  assign n46177 = n46003 ^ n43222;
  assign n46178 = n46176 & ~n46177;
  assign n46182 = n46181 ^ n46178;
  assign n46183 = n46178 ^ n46083;
  assign n46184 = n46182 & ~n46183;
  assign n46185 = n46184 ^ n46181;
  assign n46186 = n46185 ^ n46169;
  assign n46187 = ~n46173 & n46186;
  assign n46188 = n46187 ^ n46172;
  assign n46190 = n46189 ^ n46188;
  assign n46191 = n44340 ^ n35993;
  assign n46192 = n46191 ^ n40558;
  assign n46193 = n46192 ^ n34763;
  assign n46194 = n46193 ^ n46189;
  assign n46195 = n46190 & ~n46194;
  assign n46196 = n46195 ^ n46193;
  assign n46198 = n46197 ^ n46196;
  assign n46199 = n44335 ^ n35988;
  assign n46200 = n46199 ^ n40580;
  assign n46201 = n46200 ^ n34758;
  assign n46202 = n46201 ^ n46197;
  assign n46203 = ~n46198 & n46202;
  assign n46204 = n46203 ^ n46201;
  assign n46205 = n46204 ^ n46167;
  assign n46206 = ~n46168 & n46205;
  assign n46207 = n46206 ^ n46166;
  assign n46208 = n46207 ^ n46159;
  assign n46209 = ~n46163 & n46208;
  assign n46210 = n46209 ^ n46162;
  assign n46211 = n46210 ^ n46156;
  assign n46212 = n46158 & ~n46211;
  assign n46213 = n46212 ^ n46157;
  assign n46214 = n46213 ^ n46151;
  assign n46215 = ~n46153 & ~n46214;
  assign n46216 = n46215 ^ n46152;
  assign n46217 = n46216 ^ n46146;
  assign n46218 = n46148 & n46217;
  assign n46219 = n46218 ^ n46147;
  assign n46220 = n46219 ^ n46139;
  assign n46221 = ~n46143 & n46220;
  assign n46222 = n46221 ^ n46142;
  assign n46223 = n46222 ^ n46134;
  assign n46224 = ~n46138 & n46223;
  assign n46225 = n46224 ^ n46137;
  assign n46226 = n46225 ^ n2148;
  assign n46227 = ~n46133 & ~n46226;
  assign n46228 = n46227 ^ n46132;
  assign n46229 = n46228 ^ n46127;
  assign n46230 = ~n46131 & ~n46229;
  assign n46231 = n46230 ^ n46130;
  assign n46105 = ~n46078 & n46104;
  assign n45968 = n45967 ^ n45699;
  assign n45969 = ~n45701 & ~n45968;
  assign n45970 = n45969 ^ n45700;
  assign n45695 = n45587 ^ n45520;
  assign n45696 = n45695 ^ n45521;
  assign n45693 = n44746 ^ n43996;
  assign n45694 = n45693 ^ n45441;
  assign n45697 = n45696 ^ n45694;
  assign n46055 = n45970 ^ n45697;
  assign n45987 = n45986 ^ n43297;
  assign n46052 = n46051 ^ n45986;
  assign n46053 = ~n45987 & ~n46052;
  assign n46054 = n46053 ^ n43297;
  assign n46056 = n46055 ^ n46054;
  assign n46076 = n46056 ^ n42834;
  assign n46125 = n46105 ^ n46076;
  assign n46122 = n36040 ^ n2216;
  assign n46123 = n46122 ^ n40522;
  assign n46124 = n46123 ^ n34718;
  assign n46126 = n46125 ^ n46124;
  assign n46291 = n46231 ^ n46126;
  assign n47253 = n46291 ^ n45471;
  assign n46305 = n45620 ^ n45501;
  assign n46306 = n46305 ^ n45498;
  assign n47254 = n47253 ^ n46306;
  assign n46667 = n44844 ^ n44750;
  assign n46668 = n46667 ^ n45700;
  assign n46665 = n46193 ^ n46190;
  assign n46657 = n46185 ^ n46172;
  assign n46658 = n46657 ^ n46169;
  assign n46332 = n45706 ^ n44781;
  assign n46333 = n46332 ^ n44760;
  assign n46330 = n46181 ^ n46083;
  assign n46331 = n46330 ^ n46178;
  assign n46334 = n46333 ^ n46331;
  assign n46647 = n46177 ^ n46176;
  assign n46446 = n44485 ^ n43893;
  assign n46447 = n46446 ^ n45212;
  assign n45669 = n45668 ^ n45665;
  assign n45685 = n45684 ^ n45669;
  assign n46448 = n46447 ^ n45685;
  assign n46390 = n44490 ^ n43865;
  assign n46391 = n46390 ^ n45209;
  assign n46274 = n45662 ^ n45659;
  assign n46442 = n46391 ^ n46274;
  assign n46337 = n44501 ^ n43840;
  assign n46338 = n46337 ^ n45902;
  assign n46278 = n45640 ^ n45481;
  assign n46279 = n46278 ^ n45478;
  assign n46339 = n46338 ^ n46279;
  assign n46340 = n44498 ^ n43745;
  assign n46341 = n46340 ^ n45686;
  assign n46283 = n45637 ^ n45634;
  assign n46342 = n46341 ^ n46283;
  assign n46343 = n45240 ^ n44517;
  assign n46344 = n46343 ^ n45779;
  assign n46289 = n45629 ^ n45487;
  assign n46345 = n46344 ^ n46289;
  assign n46346 = n45191 ^ n44474;
  assign n46347 = n46346 ^ n45738;
  assign n46293 = n45626 ^ n45491;
  assign n46294 = n46293 ^ n45488;
  assign n46348 = n46347 ^ n46294;
  assign n46349 = n45005 ^ n44184;
  assign n46350 = n46349 ^ n45742;
  assign n46300 = n45623 ^ n45497;
  assign n46351 = n46350 ^ n46300;
  assign n46352 = n44910 ^ n44033;
  assign n46353 = n46352 ^ n45746;
  assign n46354 = n46353 ^ n46306;
  assign n46357 = n45617 ^ n45616;
  assign n46355 = n44903 ^ n44026;
  assign n46356 = n46355 ^ n45750;
  assign n46358 = n46357 ^ n46356;
  assign n46362 = n44896 ^ n44019;
  assign n46363 = n46362 ^ n45756;
  assign n46072 = n45598 ^ n45512;
  assign n46069 = n44807 ^ n43769;
  assign n46070 = n46069 ^ n45651;
  assign n46256 = n46072 ^ n46070;
  assign n45978 = n44811 ^ n44006;
  assign n45979 = n45978 ^ n45471;
  assign n45977 = n45595 ^ n45517;
  assign n45980 = n45979 ^ n45977;
  assign n45690 = n44814 ^ n43773;
  assign n45691 = n45690 ^ n45455;
  assign n45689 = n45592 ^ n1892;
  assign n45692 = n45691 ^ n45689;
  assign n45971 = n45970 ^ n45694;
  assign n45972 = ~n45697 & n45971;
  assign n45973 = n45972 ^ n45696;
  assign n45974 = n45973 ^ n45689;
  assign n45975 = ~n45692 & n45974;
  assign n45976 = n45975 ^ n45691;
  assign n46066 = n45977 ^ n45976;
  assign n46067 = ~n45980 & n46066;
  assign n46068 = n46067 ^ n45979;
  assign n46257 = n46072 ^ n46068;
  assign n46258 = n46256 & n46257;
  assign n46259 = n46258 ^ n46070;
  assign n46254 = n45606 ^ n45604;
  assign n46255 = n46254 ^ n45601;
  assign n46260 = n46259 ^ n46255;
  assign n46252 = n44803 ^ n43761;
  assign n46253 = n46252 ^ n45676;
  assign n46359 = n46255 ^ n46253;
  assign n46360 = ~n46260 & n46359;
  assign n46361 = n46360 ^ n46253;
  assign n46364 = n46363 ^ n46361;
  assign n46365 = n45609 ^ n45507;
  assign n46366 = n46365 ^ n46361;
  assign n46367 = ~n46364 & n46366;
  assign n46368 = n46367 ^ n46363;
  assign n46369 = n46368 ^ n46357;
  assign n46370 = ~n46358 & ~n46369;
  assign n46371 = n46370 ^ n46356;
  assign n46372 = n46371 ^ n46306;
  assign n46373 = n46354 & n46372;
  assign n46374 = n46373 ^ n46353;
  assign n46375 = n46374 ^ n46300;
  assign n46376 = n46351 & n46375;
  assign n46377 = n46376 ^ n46350;
  assign n46378 = n46377 ^ n46294;
  assign n46379 = n46348 & n46378;
  assign n46380 = n46379 ^ n46347;
  assign n46381 = n46380 ^ n46289;
  assign n46382 = ~n46345 & ~n46381;
  assign n46383 = n46382 ^ n46344;
  assign n46384 = n46383 ^ n46283;
  assign n46385 = n46342 & n46384;
  assign n46386 = n46385 ^ n46341;
  assign n46387 = n46386 ^ n46338;
  assign n46388 = ~n46339 & n46387;
  assign n46389 = n46388 ^ n46279;
  assign n46443 = n46389 ^ n46274;
  assign n46444 = n46442 & ~n46443;
  assign n46445 = n46444 ^ n46391;
  assign n46449 = n46448 ^ n46445;
  assign n46450 = n46449 ^ n43161;
  assign n46392 = n46391 ^ n46389;
  assign n46393 = n46392 ^ n46274;
  assign n46394 = n46393 ^ n43176;
  assign n46395 = n46386 ^ n46339;
  assign n46396 = n46395 ^ n43172;
  assign n46397 = n46383 ^ n46342;
  assign n46398 = n46397 ^ n43167;
  assign n46399 = n46380 ^ n46345;
  assign n46400 = n46399 ^ n43913;
  assign n46401 = n46377 ^ n46348;
  assign n46402 = n46401 ^ n43763;
  assign n46403 = n46374 ^ n46351;
  assign n46404 = n46403 ^ n43767;
  assign n46405 = n46371 ^ n46354;
  assign n46406 = n46405 ^ n43832;
  assign n46407 = n46368 ^ n46358;
  assign n46408 = n46407 ^ n43737;
  assign n46409 = n46365 ^ n46363;
  assign n46410 = n46409 ^ n46361;
  assign n46411 = n46410 ^ n43715;
  assign n46261 = n46260 ^ n46253;
  assign n46262 = n46261 ^ n43498;
  assign n46071 = n46070 ^ n46068;
  assign n46073 = n46072 ^ n46071;
  assign n45981 = n45980 ^ n45976;
  assign n45982 = n45981 ^ n43314;
  assign n45983 = n45973 ^ n45691;
  assign n45984 = n45983 ^ n45689;
  assign n45985 = n45984 ^ n43307;
  assign n46057 = n46055 ^ n42834;
  assign n46058 = ~n46056 & ~n46057;
  assign n46059 = n46058 ^ n42834;
  assign n46060 = n46059 ^ n45984;
  assign n46061 = n45985 & n46060;
  assign n46062 = n46061 ^ n43307;
  assign n46063 = n46062 ^ n45981;
  assign n46064 = ~n45982 & ~n46063;
  assign n46065 = n46064 ^ n43314;
  assign n46074 = n46073 ^ n46065;
  assign n46249 = n46073 ^ n43439;
  assign n46250 = ~n46074 & ~n46249;
  assign n46251 = n46250 ^ n43439;
  assign n46412 = n46261 ^ n46251;
  assign n46413 = ~n46262 & ~n46412;
  assign n46414 = n46413 ^ n43498;
  assign n46415 = n46414 ^ n46410;
  assign n46416 = n46411 & n46415;
  assign n46417 = n46416 ^ n43715;
  assign n46418 = n46417 ^ n46407;
  assign n46419 = ~n46408 & ~n46418;
  assign n46420 = n46419 ^ n43737;
  assign n46421 = n46420 ^ n46405;
  assign n46422 = n46406 & n46421;
  assign n46423 = n46422 ^ n43832;
  assign n46424 = n46423 ^ n46403;
  assign n46425 = ~n46404 & n46424;
  assign n46426 = n46425 ^ n43767;
  assign n46427 = n46426 ^ n46401;
  assign n46428 = n46402 & ~n46427;
  assign n46429 = n46428 ^ n43763;
  assign n46430 = n46429 ^ n46399;
  assign n46431 = n46400 & ~n46430;
  assign n46432 = n46431 ^ n43913;
  assign n46433 = n46432 ^ n46397;
  assign n46434 = n46398 & ~n46433;
  assign n46435 = n46434 ^ n43167;
  assign n46436 = n46435 ^ n46395;
  assign n46437 = ~n46396 & ~n46436;
  assign n46438 = n46437 ^ n43172;
  assign n46439 = n46438 ^ n46393;
  assign n46440 = n46394 & ~n46439;
  assign n46441 = n46440 ^ n43176;
  assign n46451 = n46450 ^ n46441;
  assign n46452 = n46432 ^ n46398;
  assign n46453 = n46423 ^ n46404;
  assign n46454 = n46420 ^ n43832;
  assign n46455 = n46454 ^ n46405;
  assign n46263 = n46262 ^ n46251;
  assign n46075 = n46074 ^ n43439;
  assign n46106 = ~n46076 & ~n46105;
  assign n46107 = n46059 ^ n45985;
  assign n46108 = n46106 & ~n46107;
  assign n46109 = n46062 ^ n43314;
  assign n46110 = n46109 ^ n45981;
  assign n46111 = ~n46108 & n46110;
  assign n46264 = n46075 & ~n46111;
  assign n46456 = n46263 & ~n46264;
  assign n46457 = n46414 ^ n46411;
  assign n46458 = n46456 & n46457;
  assign n46459 = n46417 ^ n46408;
  assign n46460 = n46458 & n46459;
  assign n46461 = ~n46455 & ~n46460;
  assign n46462 = ~n46453 & n46461;
  assign n46463 = n46426 ^ n43763;
  assign n46464 = n46463 ^ n46401;
  assign n46465 = ~n46462 & ~n46464;
  assign n46466 = n46429 ^ n46400;
  assign n46467 = n46465 & ~n46466;
  assign n46468 = n46452 & ~n46467;
  assign n46469 = n46435 ^ n43172;
  assign n46470 = n46469 ^ n46395;
  assign n46471 = ~n46468 & n46470;
  assign n46472 = n46438 ^ n46394;
  assign n46473 = ~n46471 & ~n46472;
  assign n46474 = n46451 & ~n46473;
  assign n46482 = n44532 ^ n43919;
  assign n46483 = n46482 ^ n45216;
  assign n46481 = n45871 ^ n45867;
  assign n46484 = n46483 ^ n46481;
  assign n46478 = n46445 ^ n45685;
  assign n46479 = ~n46448 & ~n46478;
  assign n46480 = n46479 ^ n46447;
  assign n46485 = n46484 ^ n46480;
  assign n46486 = n46485 ^ n43208;
  assign n46475 = n46449 ^ n46441;
  assign n46476 = n46450 & n46475;
  assign n46477 = n46476 ^ n43161;
  assign n46487 = n46486 ^ n46477;
  assign n46576 = n46474 & ~n46487;
  assign n46584 = n43815 ^ n43753;
  assign n46585 = n46584 ^ n45201;
  assign n46583 = n45874 ^ n45862;
  assign n46586 = n46585 ^ n46583;
  assign n46580 = n46481 ^ n46480;
  assign n46581 = n46484 & n46580;
  assign n46582 = n46581 ^ n46483;
  assign n46587 = n46586 ^ n46582;
  assign n46588 = n46587 ^ n42862;
  assign n46577 = n46485 ^ n46477;
  assign n46578 = n46486 & ~n46577;
  assign n46579 = n46578 ^ n43208;
  assign n46589 = n46588 ^ n46579;
  assign n46615 = ~n46576 & n46589;
  assign n46611 = n44484 ^ n36404;
  assign n46612 = n46611 ^ n40976;
  assign n46613 = n46612 ^ n35004;
  assign n46606 = n44543 ^ n43809;
  assign n46607 = n46606 ^ n45249;
  assign n46605 = n45877 ^ n45857;
  assign n46608 = n46607 ^ n46605;
  assign n46602 = n46583 ^ n46582;
  assign n46603 = n46586 & n46602;
  assign n46604 = n46603 ^ n46585;
  assign n46609 = n46608 ^ n46604;
  assign n46598 = n46587 ^ n46579;
  assign n46599 = n46588 & n46598;
  assign n46600 = n46599 ^ n42862;
  assign n46601 = n46600 ^ n42856;
  assign n46610 = n46609 ^ n46601;
  assign n46614 = n46613 ^ n46610;
  assign n46616 = n46615 ^ n46614;
  assign n46590 = n46589 ^ n46576;
  assign n46489 = n44251 ^ n36414;
  assign n46490 = n46489 ^ n41064;
  assign n46491 = n46490 ^ n34913;
  assign n46488 = n46487 ^ n46474;
  assign n46492 = n46491 ^ n46488;
  assign n46496 = n46473 ^ n46451;
  assign n46493 = n44255 ^ n36419;
  assign n46494 = n46493 ^ n40985;
  assign n46495 = n46494 ^ n1337;
  assign n46497 = n46496 ^ n46495;
  assign n46499 = n44260 ^ n36424;
  assign n46500 = n46499 ^ n1154;
  assign n46501 = n46500 ^ n34667;
  assign n46498 = n46472 ^ n46471;
  assign n46502 = n46501 ^ n46498;
  assign n46504 = n44448 ^ n36429;
  assign n46505 = n46504 ^ n41050;
  assign n46506 = n46505 ^ n1146;
  assign n46503 = n46470 ^ n46468;
  assign n46507 = n46506 ^ n46503;
  assign n46508 = n46467 ^ n46452;
  assign n978 = n977 ^ n941;
  assign n1012 = n1011 ^ n978;
  assign n1022 = n1021 ^ n1012;
  assign n46509 = n46508 ^ n1022;
  assign n46511 = n44266 ^ n36436;
  assign n46512 = n46511 ^ n40995;
  assign n46513 = n46512 ^ n1003;
  assign n46510 = n46466 ^ n46465;
  assign n46514 = n46513 ^ n46510;
  assign n46516 = n44271 ^ n861;
  assign n46517 = n46516 ^ n41000;
  assign n46518 = n46517 ^ n34678;
  assign n46515 = n46464 ^ n46462;
  assign n46519 = n46518 ^ n46515;
  assign n46523 = n46461 ^ n46453;
  assign n46520 = n44276 ^ n36443;
  assign n46521 = n46520 ^ n41005;
  assign n46522 = n46521 ^ n34683;
  assign n46524 = n46523 ^ n46522;
  assign n46526 = n44280 ^ n36448;
  assign n46527 = n46526 ^ n41030;
  assign n46528 = n46527 ^ n34687;
  assign n46525 = n46460 ^ n46455;
  assign n46529 = n46528 ^ n46525;
  assign n46541 = n46459 ^ n46458;
  assign n46533 = n46457 ^ n46456;
  assign n46530 = n44285 ^ n36458;
  assign n46531 = n46530 ^ n41015;
  assign n46532 = n46531 ^ n34697;
  assign n46534 = n46533 ^ n46532;
  assign n46265 = n46264 ^ n46263;
  assign n46112 = n46111 ^ n46075;
  assign n46116 = n46115 ^ n46112;
  assign n46238 = n46110 ^ n46108;
  assign n46117 = n46107 ^ n46106;
  assign n46121 = n46120 ^ n46117;
  assign n46232 = n46231 ^ n46124;
  assign n46233 = ~n46126 & ~n46232;
  assign n46234 = n46233 ^ n46125;
  assign n46235 = n46234 ^ n46117;
  assign n46236 = n46121 & n46235;
  assign n46237 = n46236 ^ n46120;
  assign n46239 = n46238 ^ n46237;
  assign n46240 = n44301 ^ n36468;
  assign n46241 = n46240 ^ n40517;
  assign n46242 = n46241 ^ n34708;
  assign n46243 = n46242 ^ n46238;
  assign n46244 = n46239 & ~n46243;
  assign n46245 = n46244 ^ n46242;
  assign n46246 = n46245 ^ n46112;
  assign n46247 = n46116 & ~n46246;
  assign n46248 = n46247 ^ n46115;
  assign n46266 = n46265 ^ n46248;
  assign n46267 = n44291 ^ n36463;
  assign n46268 = n46267 ^ n40654;
  assign n46269 = n46268 ^ n34703;
  assign n46535 = n46269 ^ n46265;
  assign n46536 = n46266 & ~n46535;
  assign n46537 = n46536 ^ n46269;
  assign n46538 = n46537 ^ n46533;
  assign n46539 = n46534 & ~n46538;
  assign n46540 = n46539 ^ n46532;
  assign n46542 = n46541 ^ n46540;
  assign n46543 = n44425 ^ n36453;
  assign n46544 = n46543 ^ n41009;
  assign n46545 = n46544 ^ n34692;
  assign n46546 = n46545 ^ n46541;
  assign n46547 = ~n46542 & n46546;
  assign n46548 = n46547 ^ n46545;
  assign n46549 = n46548 ^ n46525;
  assign n46550 = ~n46529 & n46549;
  assign n46551 = n46550 ^ n46528;
  assign n46552 = n46551 ^ n46522;
  assign n46553 = n46524 & ~n46552;
  assign n46554 = n46553 ^ n46523;
  assign n46555 = n46554 ^ n46515;
  assign n46556 = n46519 & ~n46555;
  assign n46557 = n46556 ^ n46518;
  assign n46558 = n46557 ^ n46510;
  assign n46559 = ~n46514 & n46558;
  assign n46560 = n46559 ^ n46513;
  assign n46561 = n46560 ^ n46508;
  assign n46562 = n46509 & ~n46561;
  assign n46563 = n46562 ^ n1022;
  assign n46564 = n46563 ^ n46503;
  assign n46565 = ~n46507 & n46564;
  assign n46566 = n46565 ^ n46506;
  assign n46567 = n46566 ^ n46498;
  assign n46568 = ~n46502 & n46567;
  assign n46569 = n46568 ^ n46501;
  assign n46570 = n46569 ^ n46495;
  assign n46571 = ~n46497 & ~n46570;
  assign n46572 = n46571 ^ n46496;
  assign n46573 = n46572 ^ n46488;
  assign n46574 = ~n46492 & ~n46573;
  assign n46575 = n46574 ^ n46491;
  assign n46591 = n46590 ^ n46575;
  assign n46592 = n43760 ^ n36408;
  assign n46593 = n46592 ^ n40981;
  assign n46594 = n46593 ^ n34939;
  assign n46595 = n46594 ^ n46590;
  assign n46596 = ~n46591 & n46595;
  assign n46597 = n46596 ^ n46594;
  assign n46617 = n46616 ^ n46597;
  assign n46335 = n44773 ^ n44731;
  assign n46336 = n46335 ^ n45714;
  assign n46618 = n46617 ^ n46336;
  assign n46620 = n45274 ^ n44635;
  assign n46621 = n46620 ^ n45718;
  assign n46619 = n46594 ^ n46591;
  assign n46622 = n46621 ^ n46619;
  assign n46634 = n46572 ^ n46492;
  assign n46625 = n46566 ^ n46502;
  assign n46626 = n44785 ^ n44581;
  assign n46627 = n46626 ^ n45732;
  assign n46628 = ~n46625 & n46627;
  assign n46623 = n44783 ^ n44607;
  assign n46624 = n46623 ^ n45730;
  assign n46629 = n46628 ^ n46624;
  assign n46630 = n46569 ^ n46497;
  assign n46631 = n46630 ^ n46624;
  assign n46632 = ~n46629 & ~n46631;
  assign n46633 = n46632 ^ n46628;
  assign n46635 = n46634 ^ n46633;
  assign n46636 = n44778 ^ n44623;
  assign n46637 = n46636 ^ n45723;
  assign n46638 = n46637 ^ n46634;
  assign n46639 = ~n46635 & ~n46638;
  assign n46640 = n46639 ^ n46637;
  assign n46641 = n46640 ^ n46619;
  assign n46642 = ~n46622 & n46641;
  assign n46643 = n46642 ^ n46621;
  assign n46644 = n46643 ^ n46336;
  assign n46645 = n46618 & n46644;
  assign n46646 = n46645 ^ n46617;
  assign n46648 = n46647 ^ n46646;
  assign n46649 = n45710 ^ n44768;
  assign n46650 = n46649 ^ n44825;
  assign n46651 = n46650 ^ n46647;
  assign n46652 = n46648 & ~n46651;
  assign n46653 = n46652 ^ n46650;
  assign n46654 = n46653 ^ n46331;
  assign n46655 = ~n46334 & ~n46654;
  assign n46656 = n46655 ^ n46333;
  assign n46659 = n46658 ^ n46656;
  assign n46660 = n45704 ^ n44755;
  assign n46661 = n46660 ^ n44776;
  assign n46662 = n46661 ^ n46658;
  assign n46663 = ~n46659 & ~n46662;
  assign n46664 = n46663 ^ n46661;
  assign n46666 = n46665 ^ n46664;
  assign n46797 = n46668 ^ n46666;
  assign n46760 = n46661 ^ n46659;
  assign n46761 = n46760 ^ n43790;
  assign n46789 = n46653 ^ n46334;
  assign n46762 = n46650 ^ n46648;
  assign n46763 = n46762 ^ n43796;
  assign n46764 = n46640 ^ n46622;
  assign n46765 = n46764 ^ n43755;
  assign n46773 = n46637 ^ n46635;
  assign n46766 = n46627 ^ n46625;
  assign n46767 = n43932 & ~n46766;
  assign n46768 = n46767 ^ n43804;
  assign n46769 = n46630 ^ n46629;
  assign n46770 = n46769 ^ n46767;
  assign n46771 = n46768 & ~n46770;
  assign n46772 = n46771 ^ n43804;
  assign n46774 = n46773 ^ n46772;
  assign n46775 = n46773 ^ n43803;
  assign n46776 = n46774 & ~n46775;
  assign n46777 = n46776 ^ n43803;
  assign n46778 = n46777 ^ n46764;
  assign n46779 = ~n46765 & ~n46778;
  assign n46780 = n46779 ^ n43755;
  assign n46781 = n46780 ^ n43951;
  assign n46782 = n46643 ^ n46618;
  assign n46783 = n46782 ^ n46780;
  assign n46784 = ~n46781 & ~n46783;
  assign n46785 = n46784 ^ n43951;
  assign n46786 = n46785 ^ n46762;
  assign n46787 = n46763 & n46786;
  assign n46788 = n46787 ^ n43796;
  assign n46790 = n46789 ^ n46788;
  assign n46791 = n46789 ^ n43792;
  assign n46792 = ~n46790 & ~n46791;
  assign n46793 = n46792 ^ n43792;
  assign n46794 = n46793 ^ n46760;
  assign n46795 = ~n46761 & ~n46794;
  assign n46796 = n46795 ^ n43790;
  assign n46798 = n46797 ^ n46796;
  assign n46903 = n46798 ^ n43787;
  assign n46890 = n46793 ^ n46761;
  assign n46891 = n46782 ^ n46781;
  assign n46892 = n46769 ^ n46768;
  assign n46893 = n46774 ^ n43803;
  assign n46894 = ~n46892 & n46893;
  assign n46895 = n46777 ^ n46765;
  assign n46896 = ~n46894 & ~n46895;
  assign n46897 = ~n46891 & ~n46896;
  assign n46898 = n46785 ^ n46763;
  assign n46899 = ~n46897 & n46898;
  assign n46900 = n46790 ^ n43792;
  assign n46901 = ~n46899 & ~n46900;
  assign n46902 = n46890 & n46901;
  assign n47014 = n46903 ^ n46902;
  assign n47011 = n44708 ^ n36694;
  assign n47012 = n47011 ^ n41438;
  assign n47013 = n47012 ^ n1737;
  assign n47015 = n47014 ^ n47013;
  assign n47019 = n46901 ^ n46890;
  assign n47016 = n44654 ^ n1637;
  assign n47017 = n47016 ^ n41443;
  assign n47018 = n47017 ^ n35684;
  assign n47020 = n47019 ^ n47018;
  assign n47022 = n44697 ^ n36701;
  assign n47023 = n47022 ^ n41449;
  assign n47024 = n47023 ^ n35091;
  assign n47021 = n46900 ^ n46899;
  assign n47025 = n47024 ^ n47021;
  assign n47026 = n46898 ^ n46897;
  assign n47030 = n47029 ^ n47026;
  assign n47059 = n46896 ^ n46891;
  assign n47051 = n46895 ^ n46894;
  assign n47043 = n46893 ^ n46892;
  assign n47034 = n45247 ^ n37292;
  assign n47035 = n47034 ^ n41810;
  assign n47036 = n47035 ^ n2501;
  assign n47037 = n46766 ^ n43932;
  assign n47038 = n47036 & ~n47037;
  assign n47031 = n44674 ^ n36715;
  assign n47032 = n47031 ^ n41468;
  assign n47033 = n47032 ^ n35072;
  assign n47039 = n47038 ^ n47033;
  assign n47040 = n47038 ^ n46892;
  assign n47041 = n47039 & n47040;
  assign n47042 = n47041 ^ n47033;
  assign n47044 = n47043 ^ n47042;
  assign n47045 = n44679 ^ n36720;
  assign n47046 = n47045 ^ n41472;
  assign n47047 = n47046 ^ n35069;
  assign n47048 = n47047 ^ n47042;
  assign n47049 = ~n47044 & n47048;
  assign n47050 = n47049 ^ n47047;
  assign n47052 = n47051 ^ n47050;
  assign n47053 = n44669 ^ n36711;
  assign n47054 = n47053 ^ n41463;
  assign n47055 = n47054 ^ n35065;
  assign n47056 = n47055 ^ n47051;
  assign n47057 = ~n47052 & n47056;
  assign n47058 = n47057 ^ n47055;
  assign n47060 = n47059 ^ n47058;
  assign n47061 = n44665 ^ n36733;
  assign n47062 = n47061 ^ n41459;
  assign n47063 = n47062 ^ n35061;
  assign n47064 = n47063 ^ n47059;
  assign n47065 = n47060 & ~n47064;
  assign n47066 = n47065 ^ n47063;
  assign n47067 = n47066 ^ n47026;
  assign n47068 = ~n47030 & n47067;
  assign n47069 = n47068 ^ n47029;
  assign n47070 = n47069 ^ n47021;
  assign n47071 = ~n47025 & n47070;
  assign n47072 = n47071 ^ n47024;
  assign n47073 = n47072 ^ n47019;
  assign n47074 = ~n47020 & n47073;
  assign n47075 = n47074 ^ n47018;
  assign n47076 = n47075 ^ n47014;
  assign n47077 = n47015 & ~n47076;
  assign n47078 = n47077 ^ n47013;
  assign n46904 = n46902 & ~n46903;
  assign n46799 = n46797 ^ n43787;
  assign n46800 = ~n46798 & ~n46799;
  assign n46801 = n46800 ^ n43787;
  assign n46674 = n45696 ^ n44771;
  assign n46675 = n46674 ^ n44745;
  assign n46672 = n46201 ^ n46198;
  assign n46669 = n46668 ^ n46665;
  assign n46670 = n46666 & ~n46669;
  assign n46671 = n46670 ^ n46668;
  assign n46673 = n46672 ^ n46671;
  assign n46758 = n46675 ^ n46673;
  assign n46759 = n46758 ^ n43783;
  assign n46889 = n46801 ^ n46759;
  assign n47009 = n46904 ^ n46889;
  assign n47006 = n44650 ^ n36753;
  assign n47007 = n47006 ^ n1745;
  assign n47008 = n47007 ^ n35677;
  assign n47010 = n47009 ^ n47008;
  assign n47252 = n47078 ^ n47010;
  assign n47255 = n47254 ^ n47252;
  assign n46297 = n46228 ^ n46130;
  assign n46298 = n46297 ^ n46127;
  assign n47257 = n46357 ^ n46298;
  assign n47258 = n47257 ^ n45455;
  assign n47256 = n47075 ^ n47015;
  assign n47259 = n47258 ^ n47256;
  assign n47262 = n47072 ^ n47018;
  assign n47263 = n47262 ^ n47019;
  assign n47260 = n46365 ^ n45441;
  assign n46303 = n46225 ^ n46133;
  assign n47261 = n47260 ^ n46303;
  assign n47264 = n47263 ^ n47261;
  assign n47392 = n47066 ^ n47030;
  assign n46691 = n46216 ^ n46148;
  assign n47266 = n46691 ^ n45977;
  assign n47267 = n47266 ^ n44745;
  assign n47265 = n47063 ^ n47060;
  assign n47268 = n47267 ^ n47265;
  assign n46314 = n46213 ^ n46153;
  assign n47271 = n46314 ^ n44750;
  assign n47272 = n47271 ^ n45689;
  assign n47269 = n47055 ^ n47050;
  assign n47270 = n47269 ^ n47051;
  assign n47273 = n47272 ^ n47270;
  assign n47276 = n47047 ^ n47044;
  assign n46318 = n46210 ^ n46158;
  assign n47274 = n46318 ^ n44755;
  assign n47275 = n47274 ^ n45696;
  assign n47277 = n47276 ^ n47275;
  assign n47280 = n45700 ^ n44760;
  assign n46322 = n46207 ^ n46162;
  assign n46323 = n46322 ^ n46159;
  assign n47281 = n47280 ^ n46323;
  assign n47278 = n47033 ^ n46892;
  assign n47279 = n47278 ^ n47038;
  assign n47282 = n47281 ^ n47279;
  assign n46327 = n46204 ^ n46166;
  assign n46328 = n46327 ^ n46167;
  assign n47284 = n46328 ^ n45704;
  assign n47285 = n47284 ^ n44768;
  assign n47283 = n47037 ^ n47036;
  assign n47286 = n47285 ^ n47283;
  assign n47353 = n45706 ^ n44773;
  assign n47354 = n47353 ^ n46672;
  assign n47180 = n46554 ^ n46519;
  assign n46877 = n46548 ^ n46528;
  assign n46878 = n46877 ^ n46525;
  assign n46875 = n45212 ^ n44501;
  assign n46876 = n46875 ^ n46605;
  assign n46879 = n46878 ^ n46876;
  assign n46865 = n46545 ^ n46542;
  assign n46863 = n46583 ^ n44498;
  assign n46864 = n46863 ^ n45209;
  assign n46866 = n46865 ^ n46864;
  assign n46732 = n46537 ^ n46534;
  assign n46730 = n46481 ^ n45240;
  assign n46731 = n46730 ^ n45902;
  assign n46733 = n46732 ^ n46731;
  assign n46270 = n46269 ^ n46266;
  assign n45687 = n45686 ^ n45685;
  assign n45688 = n45687 ^ n45191;
  assign n46271 = n46270 ^ n45688;
  assign n46273 = n45779 ^ n45005;
  assign n46275 = n46274 ^ n46273;
  assign n46272 = n46245 ^ n46116;
  assign n46276 = n46275 ^ n46272;
  assign n46280 = n46279 ^ n45738;
  assign n46281 = n46280 ^ n44910;
  assign n46277 = n46242 ^ n46239;
  assign n46282 = n46281 ^ n46277;
  assign n46286 = n46234 ^ n46121;
  assign n46284 = n46283 ^ n45742;
  assign n46285 = n46284 ^ n44903;
  assign n46287 = n46286 ^ n46285;
  assign n46288 = n45746 ^ n44896;
  assign n46290 = n46289 ^ n46288;
  assign n46292 = n46291 ^ n46290;
  assign n46295 = n46294 ^ n44803;
  assign n46296 = n46295 ^ n45750;
  assign n46299 = n46298 ^ n46296;
  assign n46301 = n46300 ^ n44807;
  assign n46302 = n46301 ^ n45756;
  assign n46304 = n46303 ^ n46302;
  assign n46309 = n46222 ^ n46137;
  assign n46310 = n46309 ^ n46134;
  assign n46307 = n46306 ^ n44811;
  assign n46308 = n46307 ^ n45676;
  assign n46311 = n46310 ^ n46308;
  assign n46698 = n46219 ^ n46142;
  assign n46699 = n46698 ^ n46139;
  assign n46312 = n45455 ^ n44752;
  assign n46313 = n46312 ^ n46255;
  assign n46315 = n46314 ^ n46313;
  assign n46316 = n46072 ^ n45441;
  assign n46317 = n46316 ^ n44757;
  assign n46319 = n46318 ^ n46317;
  assign n46320 = n45977 ^ n45396;
  assign n46321 = n46320 ^ n44762;
  assign n46324 = n46323 ^ n46321;
  assign n46325 = n45689 ^ n44765;
  assign n46326 = n46325 ^ n45299;
  assign n46329 = n46328 ^ n46326;
  assign n46676 = n46675 ^ n46672;
  assign n46677 = ~n46673 & n46676;
  assign n46678 = n46677 ^ n46675;
  assign n46679 = n46678 ^ n46328;
  assign n46680 = ~n46329 & n46679;
  assign n46681 = n46680 ^ n46326;
  assign n46682 = n46681 ^ n46323;
  assign n46683 = n46324 & n46682;
  assign n46684 = n46683 ^ n46321;
  assign n46685 = n46684 ^ n46317;
  assign n46686 = ~n46319 & ~n46685;
  assign n46687 = n46686 ^ n46318;
  assign n46688 = n46687 ^ n46313;
  assign n46689 = ~n46315 & ~n46688;
  assign n46690 = n46689 ^ n46314;
  assign n46692 = n46691 ^ n46690;
  assign n46693 = n45471 ^ n44746;
  assign n46694 = n46693 ^ n46365;
  assign n46695 = n46694 ^ n46691;
  assign n46696 = ~n46692 & n46695;
  assign n46697 = n46696 ^ n46694;
  assign n46700 = n46699 ^ n46697;
  assign n46701 = n46357 ^ n44814;
  assign n46702 = n46701 ^ n45651;
  assign n46703 = n46702 ^ n46699;
  assign n46704 = ~n46700 & n46703;
  assign n46705 = n46704 ^ n46702;
  assign n46706 = n46705 ^ n46310;
  assign n46707 = ~n46311 & ~n46706;
  assign n46708 = n46707 ^ n46308;
  assign n46709 = n46708 ^ n46303;
  assign n46710 = n46304 & n46709;
  assign n46711 = n46710 ^ n46302;
  assign n46712 = n46711 ^ n46296;
  assign n46713 = n46299 & n46712;
  assign n46714 = n46713 ^ n46298;
  assign n46715 = n46714 ^ n46291;
  assign n46716 = n46292 & n46715;
  assign n46717 = n46716 ^ n46290;
  assign n46718 = n46717 ^ n46286;
  assign n46719 = n46287 & ~n46718;
  assign n46720 = n46719 ^ n46285;
  assign n46721 = n46720 ^ n46277;
  assign n46722 = ~n46282 & ~n46721;
  assign n46723 = n46722 ^ n46281;
  assign n46724 = n46723 ^ n46272;
  assign n46725 = n46276 & ~n46724;
  assign n46726 = n46725 ^ n46275;
  assign n46727 = n46726 ^ n46270;
  assign n46728 = ~n46271 & n46727;
  assign n46729 = n46728 ^ n45688;
  assign n46860 = n46732 ^ n46729;
  assign n46861 = n46733 & ~n46860;
  assign n46862 = n46861 ^ n46731;
  assign n46872 = n46864 ^ n46862;
  assign n46873 = ~n46866 & n46872;
  assign n46874 = n46873 ^ n46865;
  assign n47154 = n46878 ^ n46874;
  assign n47155 = ~n46879 & n47154;
  assign n47156 = n47155 ^ n46876;
  assign n47151 = n45921 ^ n45216;
  assign n47152 = n47151 ^ n44490;
  assign n47176 = n47156 ^ n47152;
  assign n47150 = n46551 ^ n46524;
  assign n47177 = n47156 ^ n47150;
  assign n47178 = ~n47176 & ~n47177;
  assign n47179 = n47178 ^ n47152;
  assign n47181 = n47180 ^ n47179;
  assign n47174 = n45201 ^ n44485;
  assign n47175 = n47174 ^ n45924;
  assign n47182 = n47181 ^ n47175;
  assign n47183 = n47182 ^ n43893;
  assign n46880 = n46879 ^ n46874;
  assign n46881 = n46880 ^ n43840;
  assign n46867 = n46866 ^ n46862;
  assign n46734 = n46733 ^ n46729;
  assign n46735 = n46734 ^ n44517;
  assign n46736 = n46726 ^ n45688;
  assign n46737 = n46736 ^ n46270;
  assign n46738 = n46737 ^ n44474;
  assign n46849 = n46723 ^ n46276;
  assign n46739 = n46720 ^ n46282;
  assign n46740 = n46739 ^ n44033;
  assign n46741 = n46717 ^ n46285;
  assign n46742 = n46741 ^ n46286;
  assign n46743 = n46742 ^ n44026;
  assign n46744 = n46714 ^ n46290;
  assign n46745 = n46744 ^ n46291;
  assign n46746 = n46745 ^ n44019;
  assign n46835 = n46711 ^ n46299;
  assign n46747 = n46708 ^ n46304;
  assign n46748 = n46747 ^ n43769;
  assign n46749 = n46705 ^ n46311;
  assign n46750 = n46749 ^ n44006;
  assign n46751 = n46702 ^ n46700;
  assign n46752 = n46751 ^ n43773;
  assign n46821 = n46694 ^ n46692;
  assign n46816 = n46687 ^ n46315;
  assign n46753 = n46681 ^ n46321;
  assign n46754 = n46753 ^ n46323;
  assign n46755 = n46754 ^ n43979;
  assign n46756 = n46678 ^ n46329;
  assign n46757 = n46756 ^ n43779;
  assign n46802 = n46801 ^ n46758;
  assign n46803 = ~n46759 & ~n46802;
  assign n46804 = n46803 ^ n43783;
  assign n46805 = n46804 ^ n46756;
  assign n46806 = ~n46757 & ~n46805;
  assign n46807 = n46806 ^ n43779;
  assign n46808 = n46807 ^ n46754;
  assign n46809 = ~n46755 & ~n46808;
  assign n46810 = n46809 ^ n43979;
  assign n46811 = n46810 ^ n43775;
  assign n46812 = n46684 ^ n46319;
  assign n46813 = n46812 ^ n46810;
  assign n46814 = n46811 & n46813;
  assign n46815 = n46814 ^ n43775;
  assign n46817 = n46816 ^ n46815;
  assign n46818 = n46816 ^ n43989;
  assign n46819 = ~n46817 & n46818;
  assign n46820 = n46819 ^ n43989;
  assign n46822 = n46821 ^ n46820;
  assign n46823 = n46821 ^ n43996;
  assign n46824 = ~n46822 & ~n46823;
  assign n46825 = n46824 ^ n43996;
  assign n46826 = n46825 ^ n46751;
  assign n46827 = ~n46752 & n46826;
  assign n46828 = n46827 ^ n43773;
  assign n46829 = n46828 ^ n46749;
  assign n46830 = ~n46750 & ~n46829;
  assign n46831 = n46830 ^ n44006;
  assign n46832 = n46831 ^ n46747;
  assign n46833 = ~n46748 & n46832;
  assign n46834 = n46833 ^ n43769;
  assign n46836 = n46835 ^ n46834;
  assign n46837 = n46835 ^ n43761;
  assign n46838 = ~n46836 & ~n46837;
  assign n46839 = n46838 ^ n43761;
  assign n46840 = n46839 ^ n46745;
  assign n46841 = ~n46746 & ~n46840;
  assign n46842 = n46841 ^ n44019;
  assign n46843 = n46842 ^ n46742;
  assign n46844 = n46743 & ~n46843;
  assign n46845 = n46844 ^ n44026;
  assign n46846 = n46845 ^ n46739;
  assign n46847 = n46740 & n46846;
  assign n46848 = n46847 ^ n44033;
  assign n46850 = n46849 ^ n46848;
  assign n46851 = n46849 ^ n44184;
  assign n46852 = ~n46850 & ~n46851;
  assign n46853 = n46852 ^ n44184;
  assign n46854 = n46853 ^ n46737;
  assign n46855 = n46738 & ~n46854;
  assign n46856 = n46855 ^ n44474;
  assign n46857 = n46856 ^ n46734;
  assign n46858 = n46735 & n46857;
  assign n46859 = n46858 ^ n44517;
  assign n46868 = n46867 ^ n46859;
  assign n46869 = n46859 ^ n43745;
  assign n46870 = n46868 & ~n46869;
  assign n46871 = n46870 ^ n43745;
  assign n47159 = n46880 ^ n46871;
  assign n47160 = n46881 & ~n47159;
  assign n47161 = n47160 ^ n43840;
  assign n47170 = n47161 ^ n43865;
  assign n47153 = n47152 ^ n47150;
  assign n47157 = n47156 ^ n47153;
  assign n47171 = n47161 ^ n47157;
  assign n47172 = ~n47170 & ~n47171;
  assign n47173 = n47172 ^ n43865;
  assign n47184 = n47183 ^ n47173;
  assign n46882 = n46881 ^ n46871;
  assign n46883 = n46850 ^ n44184;
  assign n46884 = n46845 ^ n46740;
  assign n46885 = n46839 ^ n46746;
  assign n46886 = n46836 ^ n43761;
  assign n46887 = n46817 ^ n43989;
  assign n46888 = n46807 ^ n46755;
  assign n46905 = ~n46889 & ~n46904;
  assign n46906 = n46804 ^ n43779;
  assign n46907 = n46906 ^ n46756;
  assign n46908 = n46905 & n46907;
  assign n46909 = ~n46888 & n46908;
  assign n46910 = n46812 ^ n43775;
  assign n46911 = n46910 ^ n46810;
  assign n46912 = n46909 & n46911;
  assign n46913 = ~n46887 & n46912;
  assign n46914 = n46822 ^ n43996;
  assign n46915 = ~n46913 & ~n46914;
  assign n46916 = n46825 ^ n46752;
  assign n46917 = n46915 & n46916;
  assign n46918 = n46828 ^ n46750;
  assign n46919 = ~n46917 & ~n46918;
  assign n46920 = n46831 ^ n43769;
  assign n46921 = n46920 ^ n46747;
  assign n46922 = ~n46919 & ~n46921;
  assign n46923 = n46886 & ~n46922;
  assign n46924 = ~n46885 & n46923;
  assign n46925 = n46842 ^ n46743;
  assign n46926 = n46924 & ~n46925;
  assign n46927 = n46884 & ~n46926;
  assign n46928 = n46883 & n46927;
  assign n46929 = n46853 ^ n46738;
  assign n46930 = ~n46928 & ~n46929;
  assign n46931 = n46856 ^ n46735;
  assign n46932 = n46930 & ~n46931;
  assign n46933 = n46867 ^ n43745;
  assign n46934 = n46933 ^ n46859;
  assign n46935 = ~n46932 & ~n46934;
  assign n47149 = ~n46882 & ~n46935;
  assign n47158 = n47157 ^ n43865;
  assign n47162 = n47161 ^ n47158;
  assign n47185 = ~n47149 & ~n47162;
  assign n47290 = n47184 & ~n47185;
  assign n47299 = n46557 ^ n46514;
  assign n47296 = n47180 ^ n47175;
  assign n47297 = n47181 & n47296;
  assign n47298 = n47297 ^ n47175;
  assign n47300 = n47299 ^ n47298;
  assign n47294 = n45249 ^ n44532;
  assign n47295 = n47294 ^ n45913;
  assign n47301 = n47300 ^ n47295;
  assign n47302 = n47301 ^ n43919;
  assign n47291 = n47182 ^ n47173;
  assign n47292 = n47183 & n47291;
  assign n47293 = n47292 ^ n43893;
  assign n47303 = n47302 ^ n47293;
  assign n47304 = n47290 & ~n47303;
  assign n47313 = n45931 ^ n43753;
  assign n47314 = n47313 ^ n44791;
  assign n47309 = n47299 ^ n47295;
  assign n47310 = n47300 & ~n47309;
  assign n47311 = n47310 ^ n47295;
  assign n47217 = n46560 ^ n1022;
  assign n47218 = n47217 ^ n46508;
  assign n47312 = n47311 ^ n47218;
  assign n47315 = n47314 ^ n47312;
  assign n47305 = n47301 ^ n47293;
  assign n47306 = n47302 & ~n47305;
  assign n47307 = n47306 ^ n43919;
  assign n47308 = n47307 ^ n43815;
  assign n47316 = n47315 ^ n47308;
  assign n47350 = ~n47304 & n47316;
  assign n47345 = n46563 ^ n46507;
  assign n47340 = n44797 ^ n37252;
  assign n47341 = n47340 ^ n2405;
  assign n47342 = n47341 ^ n35583;
  assign n47343 = n47342 ^ n44787;
  assign n47344 = n47343 ^ n46606;
  assign n47346 = n47345 ^ n47344;
  assign n47336 = n47315 ^ n43815;
  assign n47337 = n47315 ^ n47307;
  assign n47338 = n47336 & n47337;
  assign n47339 = n47338 ^ n43815;
  assign n47347 = n47346 ^ n47339;
  assign n47333 = n47314 ^ n47218;
  assign n47334 = ~n47312 & n47333;
  assign n47335 = n47334 ^ n47314;
  assign n47348 = n47347 ^ n47335;
  assign n47349 = n47348 ^ n45911;
  assign n47351 = n47350 ^ n47349;
  assign n47317 = n47316 ^ n47304;
  assign n47287 = n44800 ^ n37102;
  assign n47288 = n47287 ^ n41779;
  assign n47289 = n47288 ^ n2397;
  assign n47318 = n47317 ^ n47289;
  assign n47320 = n2303 ^ n1361;
  assign n47321 = n47320 ^ n41784;
  assign n47322 = n47321 ^ n35590;
  assign n47319 = n47303 ^ n47290;
  assign n47323 = n47322 ^ n47319;
  assign n47186 = n47185 ^ n47184;
  assign n47167 = n45175 ^ n37107;
  assign n47168 = n47167 ^ n1300;
  assign n47169 = n47168 ^ n35595;
  assign n47187 = n47186 ^ n47169;
  assign n46937 = n45056 ^ n1108;
  assign n46938 = n46937 ^ n41595;
  assign n46939 = n46938 ^ n1274;
  assign n46936 = n46935 ^ n46882;
  assign n46940 = n46939 ^ n46936;
  assign n46942 = n45161 ^ n1090;
  assign n46943 = n46942 ^ n41384;
  assign n46944 = n46943 ^ n35604;
  assign n46941 = n46934 ^ n46932;
  assign n46945 = n46944 ^ n46941;
  assign n46946 = n46931 ^ n46930;
  assign n46950 = n46949 ^ n46946;
  assign n46952 = n45150 ^ n37123;
  assign n46953 = n46952 ^ n41394;
  assign n46954 = n46953 ^ n35613;
  assign n46951 = n46929 ^ n46928;
  assign n46955 = n46954 ^ n46951;
  assign n46957 = n45066 ^ n37127;
  assign n46958 = n46957 ^ n41398;
  assign n46959 = n46958 ^ n35619;
  assign n46956 = n46927 ^ n46883;
  assign n46960 = n46959 ^ n46956;
  assign n46962 = n45071 ^ n37132;
  assign n46963 = n46962 ^ n41404;
  assign n46964 = n46963 ^ n707;
  assign n46961 = n46926 ^ n46884;
  assign n46965 = n46964 ^ n46961;
  assign n46967 = n45136 ^ n37137;
  assign n46968 = n46967 ^ n41555;
  assign n46969 = n46968 ^ n35625;
  assign n46966 = n46925 ^ n46924;
  assign n46970 = n46969 ^ n46966;
  assign n46972 = n45128 ^ n37142;
  assign n46973 = n46972 ^ n41408;
  assign n46974 = n46973 ^ n35631;
  assign n46971 = n46923 ^ n46885;
  assign n46975 = n46974 ^ n46971;
  assign n46976 = n46922 ^ n46886;
  assign n46980 = n46979 ^ n46976;
  assign n46982 = n45076 ^ n37186;
  assign n46983 = n46982 ^ n41541;
  assign n46984 = n46983 ^ n35641;
  assign n46981 = n46921 ^ n46919;
  assign n46985 = n46984 ^ n46981;
  assign n47110 = n46918 ^ n46917;
  assign n46987 = n45086 ^ n37175;
  assign n46988 = n46987 ^ n41530;
  assign n46989 = n46988 ^ n35650;
  assign n46986 = n46916 ^ n46915;
  assign n46990 = n46989 ^ n46986;
  assign n46992 = n45091 ^ n37157;
  assign n46993 = n46992 ^ n41424;
  assign n46994 = n46993 ^ n35656;
  assign n46991 = n46914 ^ n46913;
  assign n46995 = n46994 ^ n46991;
  assign n46997 = n45096 ^ n2252;
  assign n46998 = n46997 ^ n41519;
  assign n46999 = n46998 ^ n35661;
  assign n46996 = n46912 ^ n46887;
  assign n47000 = n46999 ^ n46996;
  assign n47002 = n44743 ^ n2237;
  assign n47003 = n47002 ^ n41511;
  assign n47004 = n47003 ^ n35666;
  assign n47001 = n46911 ^ n46909;
  assign n47005 = n47004 ^ n47001;
  assign n47090 = n46908 ^ n46888;
  assign n47082 = n46907 ^ n46905;
  assign n47079 = n47078 ^ n47008;
  assign n47080 = n47010 & ~n47079;
  assign n47081 = n47080 ^ n47009;
  assign n47083 = n47082 ^ n47081;
  assign n47084 = n44719 ^ n36690;
  assign n47085 = n47084 ^ n41433;
  assign n47086 = n47085 ^ n1847;
  assign n47087 = n47086 ^ n47082;
  assign n47088 = ~n47083 & n47087;
  assign n47089 = n47088 ^ n47086;
  assign n47091 = n47090 ^ n47089;
  assign n47092 = n44645 ^ n36685;
  assign n47093 = n47092 ^ n41429;
  assign n47094 = n47093 ^ n35671;
  assign n47095 = n47094 ^ n47089;
  assign n47096 = n47091 & n47095;
  assign n47097 = n47096 ^ n47094;
  assign n47098 = n47097 ^ n47001;
  assign n47099 = n47005 & ~n47098;
  assign n47100 = n47099 ^ n47004;
  assign n47101 = n47100 ^ n46996;
  assign n47102 = ~n47000 & n47101;
  assign n47103 = n47102 ^ n46999;
  assign n47104 = n47103 ^ n46991;
  assign n47105 = ~n46995 & n47104;
  assign n47106 = n47105 ^ n46994;
  assign n47107 = n47106 ^ n46986;
  assign n47108 = ~n46990 & n47107;
  assign n47109 = n47108 ^ n46989;
  assign n47111 = n47110 ^ n47109;
  assign n47112 = n45081 ^ n37153;
  assign n47113 = n47112 ^ n41418;
  assign n47114 = n47113 ^ n35646;
  assign n47115 = n47114 ^ n47110;
  assign n47116 = ~n47111 & n47115;
  assign n47117 = n47116 ^ n47114;
  assign n47118 = n47117 ^ n46981;
  assign n47119 = ~n46985 & n47118;
  assign n47120 = n47119 ^ n46984;
  assign n47121 = n47120 ^ n46976;
  assign n47122 = ~n46980 & n47121;
  assign n47123 = n47122 ^ n46979;
  assign n47124 = n47123 ^ n46971;
  assign n47125 = ~n46975 & n47124;
  assign n47126 = n47125 ^ n46974;
  assign n47127 = n47126 ^ n46966;
  assign n47128 = ~n46970 & n47127;
  assign n47129 = n47128 ^ n46969;
  assign n47130 = n47129 ^ n46961;
  assign n47131 = n46965 & ~n47130;
  assign n47132 = n47131 ^ n46964;
  assign n47133 = n47132 ^ n46956;
  assign n47134 = ~n46960 & n47133;
  assign n47135 = n47134 ^ n46959;
  assign n47136 = n47135 ^ n46951;
  assign n47137 = n46955 & ~n47136;
  assign n47138 = n47137 ^ n46954;
  assign n47139 = n47138 ^ n46946;
  assign n47140 = ~n46950 & n47139;
  assign n47141 = n47140 ^ n46949;
  assign n47142 = n47141 ^ n46941;
  assign n47143 = ~n46945 & n47142;
  assign n47144 = n47143 ^ n46944;
  assign n47145 = n47144 ^ n46936;
  assign n47146 = n46940 & ~n47145;
  assign n47147 = n47146 ^ n46939;
  assign n1255 = n1245 ^ n1188;
  assign n1283 = n1282 ^ n1255;
  assign n1290 = n1289 ^ n1283;
  assign n47148 = n47147 ^ n1290;
  assign n47163 = n47162 ^ n47149;
  assign n47164 = n47163 ^ n47147;
  assign n47165 = n47148 & n47164;
  assign n47166 = n47165 ^ n1290;
  assign n47324 = n47186 ^ n47166;
  assign n47325 = ~n47187 & n47324;
  assign n47326 = n47325 ^ n47169;
  assign n47327 = n47326 ^ n47319;
  assign n47328 = ~n47323 & n47327;
  assign n47329 = n47328 ^ n47322;
  assign n47330 = n47329 ^ n47317;
  assign n47331 = n47318 & ~n47330;
  assign n47332 = n47331 ^ n47289;
  assign n47352 = n47351 ^ n47332;
  assign n47355 = n47354 ^ n47352;
  assign n47358 = n47329 ^ n47318;
  assign n47356 = n46665 ^ n45274;
  assign n47357 = n47356 ^ n45710;
  assign n47359 = n47358 ^ n47357;
  assign n47362 = n46658 ^ n44778;
  assign n47363 = n47362 ^ n45714;
  assign n47360 = n47326 ^ n47322;
  assign n47361 = n47360 ^ n47319;
  assign n47364 = n47363 ^ n47361;
  assign n47191 = n47163 ^ n1290;
  assign n47192 = n47191 ^ n47147;
  assign n47193 = n45723 ^ n44785;
  assign n47194 = n47193 ^ n46647;
  assign n47195 = ~n47192 & ~n47194;
  assign n47189 = n45718 ^ n44783;
  assign n47190 = n47189 ^ n46331;
  assign n47196 = n47195 ^ n47190;
  assign n47188 = n47187 ^ n47166;
  assign n47365 = n47190 ^ n47188;
  assign n47366 = ~n47196 & ~n47365;
  assign n47367 = n47366 ^ n47195;
  assign n47368 = n47367 ^ n47361;
  assign n47369 = ~n47364 & n47368;
  assign n47370 = n47369 ^ n47363;
  assign n47371 = n47370 ^ n47358;
  assign n47372 = n47359 & ~n47371;
  assign n47373 = n47372 ^ n47357;
  assign n47374 = n47373 ^ n47352;
  assign n47375 = ~n47355 & ~n47374;
  assign n47376 = n47375 ^ n47354;
  assign n47377 = n47376 ^ n47283;
  assign n47378 = n47286 & ~n47377;
  assign n47379 = n47378 ^ n47285;
  assign n47380 = n47379 ^ n47279;
  assign n47381 = ~n47282 & ~n47380;
  assign n47382 = n47381 ^ n47281;
  assign n47383 = n47382 ^ n47275;
  assign n47384 = n47277 & ~n47383;
  assign n47385 = n47384 ^ n47276;
  assign n47386 = n47385 ^ n47270;
  assign n47387 = ~n47273 & ~n47386;
  assign n47388 = n47387 ^ n47272;
  assign n47389 = n47388 ^ n47265;
  assign n47390 = n47268 & ~n47389;
  assign n47391 = n47390 ^ n47267;
  assign n47393 = n47392 ^ n47391;
  assign n47394 = n46072 ^ n45299;
  assign n47395 = n47394 ^ n46699;
  assign n47396 = n47395 ^ n47392;
  assign n47397 = ~n47393 & ~n47396;
  assign n47398 = n47397 ^ n47395;
  assign n47209 = n47069 ^ n47024;
  assign n47210 = n47209 ^ n47021;
  assign n47399 = n47398 ^ n47210;
  assign n47400 = n46255 ^ n45396;
  assign n47401 = n47400 ^ n46310;
  assign n47402 = n47401 ^ n47210;
  assign n47403 = n47399 & ~n47402;
  assign n47404 = n47403 ^ n47401;
  assign n47405 = n47404 ^ n47261;
  assign n47406 = n47264 & n47405;
  assign n47407 = n47406 ^ n47263;
  assign n47408 = n47407 ^ n47256;
  assign n47409 = ~n47259 & n47408;
  assign n47410 = n47409 ^ n47258;
  assign n47411 = n47410 ^ n47252;
  assign n47412 = ~n47255 & n47411;
  assign n47413 = n47412 ^ n47254;
  assign n47251 = n47086 ^ n47083;
  assign n47414 = n47413 ^ n47251;
  assign n47415 = n46300 ^ n45651;
  assign n47416 = n47415 ^ n46286;
  assign n47417 = n47416 ^ n47251;
  assign n47418 = n47414 & n47417;
  assign n47419 = n47418 ^ n47416;
  assign n47249 = n47094 ^ n47091;
  assign n47247 = n46294 ^ n45676;
  assign n47248 = n47247 ^ n46277;
  assign n47250 = n47249 ^ n47248;
  assign n47499 = n47419 ^ n47250;
  assign n47500 = n47499 ^ n44811;
  assign n47501 = n47416 ^ n47414;
  assign n47502 = n47501 ^ n44814;
  assign n47503 = n47410 ^ n47255;
  assign n47504 = n47503 ^ n44746;
  assign n47505 = n47407 ^ n47259;
  assign n47506 = n47505 ^ n44752;
  assign n47507 = n47404 ^ n47264;
  assign n47508 = n47507 ^ n44757;
  assign n47509 = n47401 ^ n47399;
  assign n47510 = n47509 ^ n44762;
  assign n47511 = n47395 ^ n47393;
  assign n47512 = n47511 ^ n44765;
  assign n47513 = n47388 ^ n47268;
  assign n47514 = n47513 ^ n44771;
  assign n47515 = n47385 ^ n47273;
  assign n47516 = n47515 ^ n44844;
  assign n47542 = n47379 ^ n47282;
  assign n47537 = n47376 ^ n47286;
  assign n47532 = n47373 ^ n47355;
  assign n47517 = n47370 ^ n47357;
  assign n47518 = n47517 ^ n47358;
  assign n47519 = n47518 ^ n44635;
  assign n47520 = n47367 ^ n47363;
  assign n47521 = n47520 ^ n47361;
  assign n47522 = n47521 ^ n44623;
  assign n47198 = n47194 ^ n47192;
  assign n47199 = n44581 & n47198;
  assign n47200 = n47199 ^ n44607;
  assign n47197 = n47196 ^ n47188;
  assign n47523 = n47199 ^ n47197;
  assign n47524 = n47200 & ~n47523;
  assign n47525 = n47524 ^ n44607;
  assign n47526 = n47525 ^ n47521;
  assign n47527 = ~n47522 & n47526;
  assign n47528 = n47527 ^ n44623;
  assign n47529 = n47528 ^ n47518;
  assign n47530 = n47519 & ~n47529;
  assign n47531 = n47530 ^ n44635;
  assign n47533 = n47532 ^ n47531;
  assign n47534 = n47532 ^ n44731;
  assign n47535 = n47533 & ~n47534;
  assign n47536 = n47535 ^ n44731;
  assign n47538 = n47537 ^ n47536;
  assign n47539 = n47537 ^ n44825;
  assign n47540 = n47538 & n47539;
  assign n47541 = n47540 ^ n44825;
  assign n47543 = n47542 ^ n47541;
  assign n47544 = n47542 ^ n44781;
  assign n47545 = n47543 & ~n47544;
  assign n47546 = n47545 ^ n44781;
  assign n47547 = n47546 ^ n44776;
  assign n47548 = n47382 ^ n47277;
  assign n47549 = n47548 ^ n47546;
  assign n47550 = n47547 & n47549;
  assign n47551 = n47550 ^ n44776;
  assign n47552 = n47551 ^ n47515;
  assign n47553 = n47516 & ~n47552;
  assign n47554 = n47553 ^ n44844;
  assign n47555 = n47554 ^ n47513;
  assign n47556 = n47514 & ~n47555;
  assign n47557 = n47556 ^ n44771;
  assign n47558 = n47557 ^ n47511;
  assign n47559 = ~n47512 & n47558;
  assign n47560 = n47559 ^ n44765;
  assign n47561 = n47560 ^ n47509;
  assign n47562 = ~n47510 & ~n47561;
  assign n47563 = n47562 ^ n44762;
  assign n47564 = n47563 ^ n47507;
  assign n47565 = n47508 & ~n47564;
  assign n47566 = n47565 ^ n44757;
  assign n47567 = n47566 ^ n47505;
  assign n47568 = n47506 & ~n47567;
  assign n47569 = n47568 ^ n44752;
  assign n47570 = n47569 ^ n47503;
  assign n47571 = ~n47504 & ~n47570;
  assign n47572 = n47571 ^ n44746;
  assign n47573 = n47572 ^ n47501;
  assign n47574 = n47502 & ~n47573;
  assign n47575 = n47574 ^ n44814;
  assign n47576 = n47575 ^ n47499;
  assign n47577 = n47500 & ~n47576;
  assign n47578 = n47577 ^ n44811;
  assign n47424 = n46272 ^ n45756;
  assign n47425 = n47424 ^ n46289;
  assign n47420 = n47419 ^ n47249;
  assign n47421 = ~n47250 & n47420;
  assign n47422 = n47421 ^ n47248;
  assign n47245 = n47097 ^ n47004;
  assign n47246 = n47245 ^ n47001;
  assign n47423 = n47422 ^ n47246;
  assign n47497 = n47425 ^ n47423;
  assign n47498 = n47497 ^ n44807;
  assign n47679 = n47578 ^ n47498;
  assign n47646 = n47575 ^ n47500;
  assign n47647 = n47572 ^ n47502;
  assign n47648 = n47563 ^ n47508;
  assign n47649 = n47560 ^ n47510;
  assign n47650 = n47557 ^ n47512;
  assign n47651 = n47551 ^ n47516;
  assign n47652 = n47548 ^ n44776;
  assign n47653 = n47652 ^ n47546;
  assign n47654 = n47543 ^ n44781;
  assign n47655 = n47533 ^ n44731;
  assign n47201 = n47200 ^ n47197;
  assign n47656 = n47525 ^ n47522;
  assign n47657 = ~n47201 & n47656;
  assign n47658 = n47528 ^ n44635;
  assign n47659 = n47658 ^ n47518;
  assign n47660 = ~n47657 & n47659;
  assign n47661 = n47655 & ~n47660;
  assign n47662 = n47538 ^ n44825;
  assign n47663 = ~n47661 & n47662;
  assign n47664 = ~n47654 & ~n47663;
  assign n47665 = ~n47653 & n47664;
  assign n47666 = n47651 & n47665;
  assign n47667 = n47554 ^ n44771;
  assign n47668 = n47667 ^ n47513;
  assign n47669 = ~n47666 & ~n47668;
  assign n47670 = n47650 & n47669;
  assign n47671 = n47649 & n47670;
  assign n47672 = n47648 & n47671;
  assign n47673 = n47566 ^ n47506;
  assign n47674 = n47672 & n47673;
  assign n47675 = n47569 ^ n47504;
  assign n47676 = ~n47674 & n47675;
  assign n47677 = n47647 & n47676;
  assign n47678 = ~n47646 & ~n47677;
  assign n47863 = n47679 ^ n47678;
  assign n47855 = n47677 ^ n47646;
  assign n47743 = n45506 ^ n37989;
  assign n47744 = n47743 ^ n42229;
  assign n47745 = n47744 ^ n36473;
  assign n47742 = n47676 ^ n47647;
  assign n47746 = n47745 ^ n47742;
  assign n47747 = n47675 ^ n47674;
  assign n47751 = n47750 ^ n47747;
  assign n47753 = n45511 ^ n37978;
  assign n47754 = n47753 ^ n2111;
  assign n47755 = n47754 ^ n35953;
  assign n47752 = n47673 ^ n47672;
  assign n47756 = n47755 ^ n47752;
  assign n47838 = n47671 ^ n47648;
  assign n47760 = n47669 ^ n47650;
  assign n47757 = n45520 ^ n37944;
  assign n47758 = n47757 ^ n42140;
  assign n47759 = n47758 ^ n1957;
  assign n47761 = n47760 ^ n47759;
  assign n47763 = n45525 ^ n1803;
  assign n47764 = n47763 ^ n42204;
  assign n47765 = n47764 ^ n35963;
  assign n47762 = n47668 ^ n47666;
  assign n47766 = n47765 ^ n47762;
  assign n47768 = n45530 ^ n37949;
  assign n47769 = n47768 ^ n42146;
  assign n47770 = n47769 ^ n35969;
  assign n47767 = n47665 ^ n47651;
  assign n47771 = n47770 ^ n47767;
  assign n47772 = n47664 ^ n47653;
  assign n47776 = n47775 ^ n47772;
  assign n47780 = n47663 ^ n47654;
  assign n47777 = n45575 ^ n37359;
  assign n47778 = n47777 ^ n42156;
  assign n47779 = n47778 ^ n35979;
  assign n47781 = n47780 ^ n47779;
  assign n47783 = n45541 ^ n37364;
  assign n47784 = n47783 ^ n42161;
  assign n47785 = n47784 ^ n35984;
  assign n47782 = n47662 ^ n47661;
  assign n47786 = n47785 ^ n47782;
  assign n47807 = n47660 ^ n47655;
  assign n47788 = n45559 ^ n37373;
  assign n47789 = n47788 ^ n42165;
  assign n47790 = n47789 ^ n35993;
  assign n47787 = n47659 ^ n47657;
  assign n47791 = n47790 ^ n47787;
  assign n47796 = n45552 ^ n37379;
  assign n47797 = n47796 ^ n42171;
  assign n47798 = n47797 ^ n35999;
  assign n47203 = n47198 ^ n44581;
  assign n47204 = n45895 ^ n38048;
  assign n47205 = n47204 ^ n42523;
  assign n47206 = n47205 ^ n2602;
  assign n47207 = n47203 & n47206;
  assign n2580 = n2579 ^ n2543;
  assign n2611 = n2610 ^ n2580;
  assign n2621 = n2620 ^ n2611;
  assign n47792 = n47207 ^ n2621;
  assign n47793 = n47207 ^ n47201;
  assign n47794 = n47792 & n47793;
  assign n47795 = n47794 ^ n2621;
  assign n47799 = n47798 ^ n47795;
  assign n47800 = n47656 ^ n47201;
  assign n47801 = n47800 ^ n47795;
  assign n47802 = n47799 & ~n47801;
  assign n47803 = n47802 ^ n47798;
  assign n47804 = n47803 ^ n47787;
  assign n47805 = ~n47791 & n47804;
  assign n47806 = n47805 ^ n47790;
  assign n47808 = n47807 ^ n47806;
  assign n47809 = n45546 ^ n37369;
  assign n47810 = n47809 ^ n42184;
  assign n47811 = n47810 ^ n35988;
  assign n47812 = n47811 ^ n47807;
  assign n47813 = ~n47808 & n47812;
  assign n47814 = n47813 ^ n47811;
  assign n47815 = n47814 ^ n47782;
  assign n47816 = ~n47786 & n47815;
  assign n47817 = n47816 ^ n47785;
  assign n47818 = n47817 ^ n47780;
  assign n47819 = ~n47781 & n47818;
  assign n47820 = n47819 ^ n47779;
  assign n47821 = n47820 ^ n47772;
  assign n47822 = n47776 & ~n47821;
  assign n47823 = n47822 ^ n47775;
  assign n47824 = n47823 ^ n47767;
  assign n47825 = ~n47771 & n47824;
  assign n47826 = n47825 ^ n47770;
  assign n47827 = n47826 ^ n47762;
  assign n47828 = n47766 & ~n47827;
  assign n47829 = n47828 ^ n47765;
  assign n47830 = n47829 ^ n47760;
  assign n47831 = n47761 & ~n47830;
  assign n47832 = n47831 ^ n47759;
  assign n1932 = n1931 ^ n1892;
  assign n1966 = n1965 ^ n1932;
  assign n1976 = n1975 ^ n1966;
  assign n47833 = n47832 ^ n1976;
  assign n47834 = n47670 ^ n47649;
  assign n47835 = n47834 ^ n47832;
  assign n47836 = n47833 & ~n47835;
  assign n47837 = n47836 ^ n1976;
  assign n47839 = n47838 ^ n47837;
  assign n47840 = n45515 ^ n37940;
  assign n47841 = n47840 ^ n42133;
  assign n47842 = n47841 ^ n2103;
  assign n47843 = n47842 ^ n47838;
  assign n47844 = ~n47839 & n47843;
  assign n47845 = n47844 ^ n47842;
  assign n47846 = n47845 ^ n47752;
  assign n47847 = n47756 & ~n47846;
  assign n47848 = n47847 ^ n47755;
  assign n47849 = n47848 ^ n47747;
  assign n47850 = n47751 & ~n47849;
  assign n47851 = n47850 ^ n47750;
  assign n47852 = n47851 ^ n47742;
  assign n47853 = ~n47746 & n47852;
  assign n47854 = n47853 ^ n47745;
  assign n47856 = n47855 ^ n47854;
  assign n47857 = n45615 ^ n37929;
  assign n47858 = n47857 ^ n42124;
  assign n47859 = n47858 ^ n36468;
  assign n47860 = n47859 ^ n47855;
  assign n47861 = ~n47856 & n47860;
  assign n47862 = n47861 ^ n47859;
  assign n47864 = n47863 ^ n47862;
  assign n48199 = n47867 ^ n47864;
  assign n47450 = n47123 ^ n46974;
  assign n47451 = n47450 ^ n46971;
  assign n48895 = n48199 ^ n47451;
  assign n48896 = n48895 ^ n46732;
  assign n48498 = n46142 ^ n2047;
  assign n48499 = n48498 ^ n42719;
  assign n48500 = n48499 ^ n36685;
  assign n48062 = n46310 ^ n45977;
  assign n48063 = n48062 ^ n47252;
  assign n48061 = n47811 ^ n47808;
  assign n48064 = n48063 ^ n48061;
  assign n48013 = n47803 ^ n47790;
  assign n48014 = n48013 ^ n47787;
  assign n48011 = n46699 ^ n45689;
  assign n48012 = n48011 ^ n47256;
  assign n48015 = n48014 ^ n48012;
  assign n48003 = n47800 ^ n47798;
  assign n48004 = n48003 ^ n47795;
  assign n47211 = n47210 ^ n45700;
  assign n47212 = n47211 ^ n46314;
  assign n47202 = n47201 ^ n2621;
  assign n47208 = n47207 ^ n47202;
  assign n47213 = n47212 ^ n47208;
  assign n47993 = n47206 ^ n47203;
  assign n47961 = n47265 ^ n45706;
  assign n47962 = n47961 ^ n46323;
  assign n47637 = n45732 ^ n44791;
  assign n47638 = n47637 ^ n46619;
  assign n47623 = n45911 ^ n45249;
  assign n47624 = n47623 ^ n46634;
  assign n47622 = n47138 ^ n46950;
  assign n47625 = n47624 ^ n47622;
  assign n47476 = n47135 ^ n46955;
  assign n47468 = n47132 ^ n46959;
  assign n47469 = n47468 ^ n46956;
  assign n47461 = n47129 ^ n46965;
  assign n47219 = n47218 ^ n45921;
  assign n47220 = n47219 ^ n45209;
  assign n47216 = n47126 ^ n46970;
  assign n47221 = n47220 ^ n47216;
  assign n47224 = n47180 ^ n46583;
  assign n47225 = n47224 ^ n45686;
  assign n47222 = n47120 ^ n46979;
  assign n47223 = n47222 ^ n46976;
  assign n47226 = n47225 ^ n47223;
  assign n47229 = n46878 ^ n45738;
  assign n47230 = n47229 ^ n45685;
  assign n47228 = n47114 ^ n47111;
  assign n47231 = n47230 ^ n47228;
  assign n47234 = n46865 ^ n46274;
  assign n47235 = n47234 ^ n45742;
  assign n47232 = n47106 ^ n46989;
  assign n47233 = n47232 ^ n46986;
  assign n47236 = n47235 ^ n47233;
  assign n47238 = n46732 ^ n46279;
  assign n47239 = n47238 ^ n45746;
  assign n47237 = n47103 ^ n46995;
  assign n47240 = n47239 ^ n47237;
  assign n47242 = n46283 ^ n45750;
  assign n47243 = n47242 ^ n46270;
  assign n47241 = n47100 ^ n47000;
  assign n47244 = n47243 ^ n47241;
  assign n47426 = n47425 ^ n47246;
  assign n47427 = ~n47423 & n47426;
  assign n47428 = n47427 ^ n47425;
  assign n47429 = n47428 ^ n47241;
  assign n47430 = n47244 & n47429;
  assign n47431 = n47430 ^ n47243;
  assign n47432 = n47431 ^ n47239;
  assign n47433 = ~n47240 & n47432;
  assign n47434 = n47433 ^ n47237;
  assign n47435 = n47434 ^ n47233;
  assign n47436 = n47236 & ~n47435;
  assign n47437 = n47436 ^ n47235;
  assign n47438 = n47437 ^ n47228;
  assign n47439 = ~n47231 & n47438;
  assign n47440 = n47439 ^ n47230;
  assign n47227 = n47117 ^ n46985;
  assign n47441 = n47440 ^ n47227;
  assign n47442 = n46481 ^ n45779;
  assign n47443 = n47442 ^ n47150;
  assign n47444 = n47443 ^ n47227;
  assign n47445 = ~n47441 & n47444;
  assign n47446 = n47445 ^ n47443;
  assign n47447 = n47446 ^ n47223;
  assign n47448 = ~n47226 & ~n47447;
  assign n47449 = n47448 ^ n47225;
  assign n47452 = n47451 ^ n47449;
  assign n47453 = n47299 ^ n45902;
  assign n47454 = n47453 ^ n46605;
  assign n47455 = n47454 ^ n47451;
  assign n47456 = n47452 & n47455;
  assign n47457 = n47456 ^ n47454;
  assign n47458 = n47457 ^ n47216;
  assign n47459 = ~n47221 & ~n47458;
  assign n47460 = n47459 ^ n47220;
  assign n47462 = n47461 ^ n47460;
  assign n47463 = n45924 ^ n45212;
  assign n47464 = n47463 ^ n47345;
  assign n47465 = n47464 ^ n47461;
  assign n47466 = ~n47462 & ~n47465;
  assign n47467 = n47466 ^ n47464;
  assign n47470 = n47469 ^ n47467;
  assign n47471 = n45913 ^ n45216;
  assign n47472 = n47471 ^ n46625;
  assign n47473 = n47472 ^ n47469;
  assign n47474 = ~n47470 & ~n47473;
  assign n47475 = n47474 ^ n47472;
  assign n47477 = n47476 ^ n47475;
  assign n47214 = n45931 ^ n45201;
  assign n47215 = n47214 ^ n46630;
  assign n47619 = n47476 ^ n47215;
  assign n47620 = ~n47477 & ~n47619;
  assign n47621 = n47620 ^ n47215;
  assign n47633 = n47622 ^ n47621;
  assign n47634 = n47625 & ~n47633;
  assign n47635 = n47634 ^ n47624;
  assign n47631 = n47141 ^ n46944;
  assign n47632 = n47631 ^ n46941;
  assign n47636 = n47635 ^ n47632;
  assign n47639 = n47638 ^ n47636;
  assign n47640 = n47639 ^ n43753;
  assign n47626 = n47625 ^ n47621;
  assign n47478 = n47477 ^ n47215;
  assign n47479 = n47478 ^ n44485;
  assign n47480 = n47472 ^ n47470;
  assign n47481 = n47480 ^ n44490;
  assign n47482 = n47464 ^ n47462;
  assign n47483 = n47482 ^ n44501;
  assign n47484 = n47457 ^ n47221;
  assign n47485 = n47484 ^ n44498;
  assign n47486 = n47454 ^ n47452;
  assign n47487 = n47486 ^ n45240;
  assign n47599 = n47446 ^ n47226;
  assign n47594 = n47443 ^ n47441;
  assign n47488 = n47437 ^ n47231;
  assign n47489 = n47488 ^ n44910;
  assign n47490 = n47434 ^ n47235;
  assign n47491 = n47490 ^ n47233;
  assign n47492 = n47491 ^ n44903;
  assign n47493 = n47431 ^ n47240;
  assign n47494 = n47493 ^ n44896;
  assign n47495 = n47428 ^ n47244;
  assign n47496 = n47495 ^ n44803;
  assign n47579 = n47578 ^ n47497;
  assign n47580 = n47498 & n47579;
  assign n47581 = n47580 ^ n44807;
  assign n47582 = n47581 ^ n47495;
  assign n47583 = n47496 & ~n47582;
  assign n47584 = n47583 ^ n44803;
  assign n47585 = n47584 ^ n47493;
  assign n47586 = ~n47494 & ~n47585;
  assign n47587 = n47586 ^ n44896;
  assign n47588 = n47587 ^ n47491;
  assign n47589 = ~n47492 & ~n47588;
  assign n47590 = n47589 ^ n44903;
  assign n47591 = n47590 ^ n47488;
  assign n47592 = n47489 & ~n47591;
  assign n47593 = n47592 ^ n44910;
  assign n47595 = n47594 ^ n47593;
  assign n47596 = n47594 ^ n45005;
  assign n47597 = n47595 & n47596;
  assign n47598 = n47597 ^ n45005;
  assign n47600 = n47599 ^ n47598;
  assign n47601 = n47599 ^ n45191;
  assign n47602 = n47600 & ~n47601;
  assign n47603 = n47602 ^ n45191;
  assign n47604 = n47603 ^ n47486;
  assign n47605 = n47487 & n47604;
  assign n47606 = n47605 ^ n45240;
  assign n47607 = n47606 ^ n47484;
  assign n47608 = n47485 & ~n47607;
  assign n47609 = n47608 ^ n44498;
  assign n47610 = n47609 ^ n47482;
  assign n47611 = ~n47483 & n47610;
  assign n47612 = n47611 ^ n44501;
  assign n47613 = n47612 ^ n47480;
  assign n47614 = n47481 & ~n47613;
  assign n47615 = n47614 ^ n44490;
  assign n47616 = n47615 ^ n47478;
  assign n47617 = ~n47479 & n47616;
  assign n47618 = n47617 ^ n44485;
  assign n47627 = n47626 ^ n47618;
  assign n47628 = n47626 ^ n44532;
  assign n47629 = n47627 & ~n47628;
  assign n47630 = n47629 ^ n44532;
  assign n47641 = n47640 ^ n47630;
  assign n47642 = n47612 ^ n44490;
  assign n47643 = n47642 ^ n47480;
  assign n47644 = n47584 ^ n44896;
  assign n47645 = n47644 ^ n47493;
  assign n47680 = ~n47678 & n47679;
  assign n47681 = n47581 ^ n47496;
  assign n47682 = ~n47680 & n47681;
  assign n47683 = ~n47645 & n47682;
  assign n47684 = n47587 ^ n47492;
  assign n47685 = n47683 & n47684;
  assign n47686 = n47590 ^ n47489;
  assign n47687 = ~n47685 & ~n47686;
  assign n47688 = n47595 ^ n45005;
  assign n47689 = n47687 & ~n47688;
  assign n47690 = n47600 ^ n45191;
  assign n47691 = ~n47689 & n47690;
  assign n47692 = n47603 ^ n45240;
  assign n47693 = n47692 ^ n47486;
  assign n47694 = n47691 & ~n47693;
  assign n47695 = n47606 ^ n44498;
  assign n47696 = n47695 ^ n47484;
  assign n47697 = ~n47694 & ~n47696;
  assign n47698 = n47609 ^ n44501;
  assign n47699 = n47698 ^ n47482;
  assign n47700 = ~n47697 & ~n47699;
  assign n47701 = ~n47643 & ~n47700;
  assign n47702 = n47615 ^ n44485;
  assign n47703 = n47702 ^ n47478;
  assign n47704 = ~n47701 & ~n47703;
  assign n47705 = n47627 ^ n44532;
  assign n47706 = n47704 & ~n47705;
  assign n47957 = ~n47641 & ~n47706;
  assign n47952 = n47144 ^ n46939;
  assign n47953 = n47952 ^ n46936;
  assign n47949 = n46617 ^ n44787;
  assign n47950 = n47949 ^ n45730;
  assign n47946 = n47638 ^ n47632;
  assign n47947 = ~n47636 & n47946;
  assign n47948 = n47947 ^ n47638;
  assign n47951 = n47950 ^ n47948;
  assign n47954 = n47953 ^ n47951;
  assign n47955 = n47954 ^ n44543;
  assign n47943 = n47639 ^ n47630;
  assign n47944 = n47640 & n47943;
  assign n47945 = n47944 ^ n43753;
  assign n47956 = n47955 ^ n47945;
  assign n47958 = n47957 ^ n47956;
  assign n47940 = n45737 ^ n2460;
  assign n47941 = n47940 ^ n42477;
  assign n47942 = n47941 ^ n36404;
  assign n47959 = n47958 ^ n47942;
  assign n47708 = n45840 ^ n37874;
  assign n47709 = n47708 ^ n42427;
  assign n47710 = n47709 ^ n36408;
  assign n47707 = n47706 ^ n47641;
  assign n47711 = n47710 ^ n47707;
  assign n47929 = n47705 ^ n47704;
  assign n47713 = n45850 ^ n1397;
  assign n47714 = n47713 ^ n42460;
  assign n47715 = n47714 ^ n36419;
  assign n47712 = n47703 ^ n47701;
  assign n47716 = n47715 ^ n47712;
  assign n47918 = n47700 ^ n47643;
  assign n47720 = n47699 ^ n47697;
  assign n47721 = n47720 ^ n47719;
  assign n47723 = n45866 ^ n37888;
  assign n47724 = n47723 ^ n42437;
  assign n47725 = n47724 ^ n977;
  assign n47722 = n47696 ^ n47694;
  assign n47726 = n47725 ^ n47722;
  assign n47728 = n45668 ^ n37892;
  assign n47729 = n47728 ^ n869;
  assign n47730 = n47729 ^ n36436;
  assign n47727 = n47693 ^ n47691;
  assign n47731 = n47730 ^ n47727;
  assign n47901 = n47690 ^ n47689;
  assign n47733 = n45481 ^ n752;
  assign n47734 = n47733 ^ n42104;
  assign n47735 = n47734 ^ n36443;
  assign n47732 = n47688 ^ n47687;
  assign n47736 = n47735 ^ n47732;
  assign n47738 = n45637 ^ n37905;
  assign n47739 = n47738 ^ n42109;
  assign n47740 = n47739 ^ n36448;
  assign n47737 = n47686 ^ n47685;
  assign n47741 = n47740 ^ n47737;
  assign n47887 = n47684 ^ n47683;
  assign n47879 = n47682 ^ n47645;
  assign n47871 = n47681 ^ n47680;
  assign n47868 = n47867 ^ n47863;
  assign n47869 = ~n47864 & n47868;
  assign n47870 = n47869 ^ n47867;
  assign n47872 = n47871 ^ n47870;
  assign n47873 = n45495 ^ n37920;
  assign n47874 = n47873 ^ n42118;
  assign n47875 = n47874 ^ n36463;
  assign n47876 = n47875 ^ n47871;
  assign n47877 = n47872 & ~n47876;
  assign n47878 = n47877 ^ n47875;
  assign n47880 = n47879 ^ n47878;
  assign n47881 = n45491 ^ n37915;
  assign n47882 = n47881 ^ n42251;
  assign n47883 = n47882 ^ n36458;
  assign n47884 = n47883 ^ n47879;
  assign n47885 = n47880 & ~n47884;
  assign n47886 = n47885 ^ n47883;
  assign n47888 = n47887 ^ n47886;
  assign n47889 = n45486 ^ n37910;
  assign n47890 = n47889 ^ n42114;
  assign n47891 = n47890 ^ n36453;
  assign n47892 = n47891 ^ n47887;
  assign n47893 = ~n47888 & n47892;
  assign n47894 = n47893 ^ n47891;
  assign n47895 = n47894 ^ n47737;
  assign n47896 = ~n47741 & n47895;
  assign n47897 = n47896 ^ n47740;
  assign n47898 = n47897 ^ n47732;
  assign n47899 = n47736 & ~n47898;
  assign n47900 = n47899 ^ n47735;
  assign n47902 = n47901 ^ n47900;
  assign n47903 = n45662 ^ n37898;
  assign n47904 = n47903 ^ n42099;
  assign n47905 = n47904 ^ n861;
  assign n47906 = n47905 ^ n47901;
  assign n47907 = n47902 & ~n47906;
  assign n47908 = n47907 ^ n47905;
  assign n47909 = n47908 ^ n47727;
  assign n47910 = ~n47731 & n47909;
  assign n47911 = n47910 ^ n47730;
  assign n47912 = n47911 ^ n47722;
  assign n47913 = ~n47726 & n47912;
  assign n47914 = n47913 ^ n47725;
  assign n47915 = n47914 ^ n47720;
  assign n47916 = n47721 & ~n47915;
  assign n47917 = n47916 ^ n47719;
  assign n47919 = n47918 ^ n47917;
  assign n47920 = n45856 ^ n1382;
  assign n47921 = n47920 ^ n42432;
  assign n47922 = n47921 ^ n36424;
  assign n47923 = n47922 ^ n47918;
  assign n47924 = n47919 & ~n47923;
  assign n47925 = n47924 ^ n47922;
  assign n47926 = n47925 ^ n47712;
  assign n47927 = n47716 & ~n47926;
  assign n47928 = n47927 ^ n47715;
  assign n47930 = n47929 ^ n47928;
  assign n47931 = n45845 ^ n37878;
  assign n47932 = n47931 ^ n42468;
  assign n47933 = n47932 ^ n36414;
  assign n47934 = n47933 ^ n47929;
  assign n47935 = n47930 & ~n47934;
  assign n47936 = n47935 ^ n47933;
  assign n47937 = n47936 ^ n47707;
  assign n47938 = ~n47711 & n47937;
  assign n47939 = n47938 ^ n47710;
  assign n47960 = n47959 ^ n47939;
  assign n47963 = n47962 ^ n47960;
  assign n47965 = n46328 ^ n45710;
  assign n47966 = n47965 ^ n47270;
  assign n47964 = n47936 ^ n47711;
  assign n47967 = n47966 ^ n47964;
  assign n47970 = n47933 ^ n47930;
  assign n47968 = n47276 ^ n45714;
  assign n47969 = n47968 ^ n46672;
  assign n47971 = n47970 ^ n47969;
  assign n47974 = n47922 ^ n47919;
  assign n47975 = n46658 ^ n45723;
  assign n47976 = n47975 ^ n47283;
  assign n47977 = ~n47974 & n47976;
  assign n47972 = n46665 ^ n45718;
  assign n47973 = n47972 ^ n47279;
  assign n47978 = n47977 ^ n47973;
  assign n47979 = n47925 ^ n47715;
  assign n47980 = n47979 ^ n47712;
  assign n47981 = n47980 ^ n47973;
  assign n47982 = n47978 & ~n47981;
  assign n47983 = n47982 ^ n47977;
  assign n47984 = n47983 ^ n47969;
  assign n47985 = ~n47971 & ~n47984;
  assign n47986 = n47985 ^ n47970;
  assign n47987 = n47986 ^ n47964;
  assign n47988 = n47967 & ~n47987;
  assign n47989 = n47988 ^ n47966;
  assign n47990 = n47989 ^ n47960;
  assign n47991 = n47963 & ~n47990;
  assign n47992 = n47991 ^ n47962;
  assign n47994 = n47993 ^ n47992;
  assign n47995 = n46318 ^ n45704;
  assign n47996 = n47995 ^ n47392;
  assign n47997 = n47996 ^ n47993;
  assign n47998 = n47994 & n47997;
  assign n47999 = n47998 ^ n47996;
  assign n48000 = n47999 ^ n47208;
  assign n48001 = ~n47213 & n48000;
  assign n48002 = n48001 ^ n47212;
  assign n48005 = n48004 ^ n48002;
  assign n48006 = n47263 ^ n46691;
  assign n48007 = n48006 ^ n45696;
  assign n48008 = n48007 ^ n48004;
  assign n48009 = ~n48005 & n48008;
  assign n48010 = n48009 ^ n48007;
  assign n48058 = n48014 ^ n48010;
  assign n48059 = ~n48015 & n48058;
  assign n48060 = n48059 ^ n48012;
  assign n48065 = n48064 ^ n48060;
  assign n48016 = n48015 ^ n48010;
  assign n48017 = n48016 ^ n44750;
  assign n48050 = n48007 ^ n48005;
  assign n48045 = n47999 ^ n47213;
  assign n48040 = n47996 ^ n47994;
  assign n48035 = n47989 ^ n47963;
  assign n48018 = n47986 ^ n47967;
  assign n48019 = n48018 ^ n45274;
  assign n48020 = n47976 ^ n47974;
  assign n48021 = n44785 & ~n48020;
  assign n48022 = n48021 ^ n44783;
  assign n48023 = n47980 ^ n47978;
  assign n48024 = n48023 ^ n48021;
  assign n48025 = ~n48022 & ~n48024;
  assign n48026 = n48025 ^ n44783;
  assign n48027 = n48026 ^ n44778;
  assign n48028 = n47983 ^ n47971;
  assign n48029 = n48028 ^ n48026;
  assign n48030 = n48027 & ~n48029;
  assign n48031 = n48030 ^ n44778;
  assign n48032 = n48031 ^ n48018;
  assign n48033 = n48019 & ~n48032;
  assign n48034 = n48033 ^ n45274;
  assign n48036 = n48035 ^ n48034;
  assign n48037 = n48035 ^ n44773;
  assign n48038 = ~n48036 & ~n48037;
  assign n48039 = n48038 ^ n44773;
  assign n48041 = n48040 ^ n48039;
  assign n48042 = n48040 ^ n44768;
  assign n48043 = n48041 & n48042;
  assign n48044 = n48043 ^ n44768;
  assign n48046 = n48045 ^ n48044;
  assign n48047 = n48045 ^ n44760;
  assign n48048 = ~n48046 & n48047;
  assign n48049 = n48048 ^ n44760;
  assign n48051 = n48050 ^ n48049;
  assign n48052 = n48050 ^ n44755;
  assign n48053 = n48051 & n48052;
  assign n48054 = n48053 ^ n44755;
  assign n48055 = n48054 ^ n48016;
  assign n48056 = n48017 & n48055;
  assign n48057 = n48056 ^ n44750;
  assign n48066 = n48065 ^ n48057;
  assign n48067 = n48066 ^ n44745;
  assign n48068 = n48051 ^ n44755;
  assign n48069 = n48041 ^ n44768;
  assign n48070 = n48036 ^ n44773;
  assign n48071 = n48031 ^ n45274;
  assign n48072 = n48071 ^ n48018;
  assign n48073 = n48023 ^ n48022;
  assign n48074 = n48028 ^ n48027;
  assign n48075 = n48073 & n48074;
  assign n48076 = ~n48072 & ~n48075;
  assign n48077 = ~n48070 & ~n48076;
  assign n48078 = n48069 & ~n48077;
  assign n48079 = n48046 ^ n44760;
  assign n48080 = ~n48078 & n48079;
  assign n48081 = n48068 & n48080;
  assign n48082 = n48054 ^ n48017;
  assign n48083 = n48081 & ~n48082;
  assign n48160 = n48067 & ~n48083;
  assign n48169 = n47814 ^ n47785;
  assign n48170 = n48169 ^ n47782;
  assign n48167 = n46303 ^ n46072;
  assign n48168 = n48167 ^ n47251;
  assign n48171 = n48170 ^ n48168;
  assign n48164 = n48063 ^ n48060;
  assign n48165 = n48064 & ~n48164;
  assign n48166 = n48165 ^ n48061;
  assign n48172 = n48171 ^ n48166;
  assign n48173 = n48172 ^ n45299;
  assign n48161 = n48065 ^ n44745;
  assign n48162 = n48066 & ~n48161;
  assign n48163 = n48162 ^ n44745;
  assign n48174 = n48173 ^ n48163;
  assign n48407 = n48160 & n48174;
  assign n48327 = n48172 ^ n48163;
  assign n48328 = ~n48173 & ~n48327;
  assign n48329 = n48328 ^ n45299;
  assign n48242 = n47249 ^ n46298;
  assign n48243 = n48242 ^ n46255;
  assign n48239 = n47817 ^ n47779;
  assign n48240 = n48239 ^ n47780;
  assign n48236 = n48170 ^ n48166;
  assign n48237 = ~n48171 & n48236;
  assign n48238 = n48237 ^ n48168;
  assign n48241 = n48240 ^ n48238;
  assign n48325 = n48243 ^ n48241;
  assign n48326 = n48325 ^ n45396;
  assign n48406 = n48329 ^ n48326;
  assign n48497 = n48407 ^ n48406;
  assign n48501 = n48500 ^ n48497;
  assign n48176 = n46146 ^ n38244;
  assign n48177 = n48176 ^ n42793;
  assign n48178 = n48177 ^ n36690;
  assign n48175 = n48174 ^ n48160;
  assign n48179 = n48178 ^ n48175;
  assign n48085 = n46151 ^ n38310;
  assign n48086 = n48085 ^ n42723;
  assign n48087 = n48086 ^ n36753;
  assign n48084 = n48083 ^ n48067;
  assign n48088 = n48087 ^ n48084;
  assign n48090 = n46156 ^ n38249;
  assign n48091 = n48090 ^ n42782;
  assign n48092 = n48091 ^ n36694;
  assign n48089 = n48082 ^ n48081;
  assign n48093 = n48092 ^ n48089;
  assign n48095 = n46162 ^ n38254;
  assign n48096 = n48095 ^ n42728;
  assign n48097 = n48096 ^ n1637;
  assign n48094 = n48080 ^ n48068;
  assign n48098 = n48097 ^ n48094;
  assign n48100 = n46166 ^ n38259;
  assign n48101 = n48100 ^ n42771;
  assign n48102 = n48101 ^ n36701;
  assign n48099 = n48079 ^ n48078;
  assign n48103 = n48102 ^ n48099;
  assign n48105 = n46201 ^ n38263;
  assign n48106 = n48105 ^ n42734;
  assign n48107 = n48106 ^ n36706;
  assign n48104 = n48077 ^ n48069;
  assign n48108 = n48107 ^ n48104;
  assign n48110 = n46193 ^ n38290;
  assign n48111 = n48110 ^ n42739;
  assign n48112 = n48111 ^ n36733;
  assign n48109 = n48076 ^ n48070;
  assign n48113 = n48112 ^ n48109;
  assign n48115 = n46172 ^ n38268;
  assign n48116 = n48115 ^ n42743;
  assign n48117 = n48116 ^ n36711;
  assign n48114 = n48075 ^ n48072;
  assign n48118 = n48117 ^ n48114;
  assign n48131 = n46181 ^ n38277;
  assign n48132 = n48131 ^ n42753;
  assign n48133 = n48132 ^ n36720;
  assign n48122 = n46613 ^ n38827;
  assign n48123 = n48122 ^ n43204;
  assign n48124 = n48123 ^ n37292;
  assign n48125 = n48020 ^ n44785;
  assign n48126 = n48124 & ~n48125;
  assign n48119 = n46176 ^ n38272;
  assign n48120 = n48119 ^ n42749;
  assign n48121 = n48120 ^ n36715;
  assign n48127 = n48126 ^ n48121;
  assign n48128 = n48126 ^ n48073;
  assign n48129 = n48127 & ~n48128;
  assign n48130 = n48129 ^ n48121;
  assign n48134 = n48133 ^ n48130;
  assign n48135 = n48074 ^ n48073;
  assign n48136 = n48135 ^ n48130;
  assign n48137 = n48134 & n48136;
  assign n48138 = n48137 ^ n48133;
  assign n48139 = n48138 ^ n48114;
  assign n48140 = n48118 & ~n48139;
  assign n48141 = n48140 ^ n48117;
  assign n48142 = n48141 ^ n48109;
  assign n48143 = ~n48113 & n48142;
  assign n48144 = n48143 ^ n48112;
  assign n48145 = n48144 ^ n48104;
  assign n48146 = ~n48108 & n48145;
  assign n48147 = n48146 ^ n48107;
  assign n48148 = n48147 ^ n48099;
  assign n48149 = n48103 & ~n48148;
  assign n48150 = n48149 ^ n48102;
  assign n48151 = n48150 ^ n48094;
  assign n48152 = ~n48098 & n48151;
  assign n48153 = n48152 ^ n48097;
  assign n48154 = n48153 ^ n48089;
  assign n48155 = n48093 & ~n48154;
  assign n48156 = n48155 ^ n48092;
  assign n48157 = n48156 ^ n48084;
  assign n48158 = ~n48088 & n48157;
  assign n48159 = n48158 ^ n48087;
  assign n48502 = n48175 ^ n48159;
  assign n48503 = n48179 & ~n48502;
  assign n48504 = n48503 ^ n48178;
  assign n48505 = n48504 ^ n48497;
  assign n48506 = ~n48501 & n48505;
  assign n48507 = n48506 ^ n48500;
  assign n48493 = n46137 ^ n2065;
  assign n48494 = n48493 ^ n42714;
  assign n48495 = n48494 ^ n2237;
  assign n48892 = n48507 ^ n48495;
  assign n48244 = n48243 ^ n48240;
  assign n48245 = n48241 & ~n48244;
  assign n48246 = n48245 ^ n48243;
  assign n48234 = n47820 ^ n47776;
  assign n48232 = n46365 ^ n46291;
  assign n48233 = n48232 ^ n47246;
  assign n48235 = n48234 ^ n48233;
  assign n48333 = n48246 ^ n48235;
  assign n48330 = n48329 ^ n48325;
  assign n48331 = ~n48326 & n48330;
  assign n48332 = n48331 ^ n45396;
  assign n48334 = n48333 ^ n48332;
  assign n48409 = n48334 ^ n45441;
  assign n48408 = ~n48406 & n48407;
  assign n48492 = n48409 ^ n48408;
  assign n48893 = n48892 ^ n48492;
  assign n48816 = n48504 ^ n48501;
  assign n48203 = n47859 ^ n47856;
  assign n48814 = n48203 ^ n47223;
  assign n48815 = n48814 ^ n46270;
  assign n48817 = n48816 ^ n48815;
  assign n48207 = n47851 ^ n47746;
  assign n48818 = n48207 ^ n46272;
  assign n48819 = n48818 ^ n47227;
  assign n48180 = n48179 ^ n48159;
  assign n48820 = n48819 ^ n48180;
  assign n48823 = n48153 ^ n48093;
  assign n48821 = n47233 ^ n46286;
  assign n48210 = n47845 ^ n47756;
  assign n48822 = n48821 ^ n48210;
  assign n48824 = n48823 ^ n48822;
  assign n48181 = n47842 ^ n47839;
  assign n48825 = n48181 ^ n47237;
  assign n48826 = n48825 ^ n46291;
  assign n48766 = n48150 ^ n48098;
  assign n48827 = n48826 ^ n48766;
  assign n48221 = n47829 ^ n47761;
  assign n48830 = n48221 ^ n47246;
  assign n48831 = n48830 ^ n46303;
  assign n48829 = n48144 ^ n48108;
  assign n48832 = n48831 ^ n48829;
  assign n48851 = n48138 ^ n48117;
  assign n48852 = n48851 ^ n48114;
  assign n48835 = n48135 ^ n48134;
  assign n48833 = n47252 ^ n46691;
  assign n48834 = n48833 ^ n48234;
  assign n48836 = n48835 ^ n48834;
  assign n48839 = n48121 ^ n48073;
  assign n48840 = n48839 ^ n48126;
  assign n48837 = n48240 ^ n46314;
  assign n48838 = n48837 ^ n47256;
  assign n48841 = n48840 ^ n48838;
  assign n48750 = n48125 ^ n48124;
  assign n48687 = n46331 ^ n45730;
  assign n48688 = n48687 ^ n47352;
  assign n48685 = n47914 ^ n47719;
  assign n48686 = n48685 ^ n47720;
  assign n48689 = n48688 ^ n48686;
  assign n48648 = n46647 ^ n45732;
  assign n48649 = n48648 ^ n47358;
  assign n48647 = n47911 ^ n47726;
  assign n48650 = n48649 ^ n48647;
  assign n48391 = n47897 ^ n47735;
  assign n48392 = n48391 ^ n47732;
  assign n48389 = n47192 ^ n45913;
  assign n48390 = n48389 ^ n46634;
  assign n48393 = n48392 ^ n48390;
  assign n48298 = n47894 ^ n47741;
  assign n48296 = n46630 ^ n45924;
  assign n48297 = n48296 ^ n47953;
  assign n48299 = n48298 ^ n48297;
  assign n48188 = n47632 ^ n45921;
  assign n48189 = n48188 ^ n46625;
  assign n48187 = n47891 ^ n47888;
  assign n48190 = n48189 ^ n48187;
  assign n48193 = n47883 ^ n47880;
  assign n48191 = n47622 ^ n47345;
  assign n48192 = n48191 ^ n46605;
  assign n48194 = n48193 ^ n48192;
  assign n48197 = n47875 ^ n47872;
  assign n48195 = n47476 ^ n47218;
  assign n48196 = n48195 ^ n46583;
  assign n48198 = n48197 ^ n48196;
  assign n48200 = n47469 ^ n46481;
  assign n48201 = n48200 ^ n47299;
  assign n48202 = n48201 ^ n48199;
  assign n48204 = n47180 ^ n45685;
  assign n48205 = n48204 ^ n47461;
  assign n48206 = n48205 ^ n48203;
  assign n48268 = n47848 ^ n47751;
  assign n48208 = n46865 ^ n46283;
  assign n48209 = n48208 ^ n47223;
  assign n48211 = n48210 ^ n48209;
  assign n48212 = n47227 ^ n46732;
  assign n48213 = n48212 ^ n46289;
  assign n48214 = n48213 ^ n48181;
  assign n48217 = n47834 ^ n47833;
  assign n48215 = n47228 ^ n46294;
  assign n48216 = n48215 ^ n46270;
  assign n48218 = n48217 ^ n48216;
  assign n48219 = n47233 ^ n46300;
  assign n48220 = n48219 ^ n46272;
  assign n48222 = n48221 ^ n48220;
  assign n48225 = n47826 ^ n47765;
  assign n48226 = n48225 ^ n47762;
  assign n48223 = n47237 ^ n46277;
  assign n48224 = n48223 ^ n46306;
  assign n48227 = n48226 ^ n48224;
  assign n48229 = n47241 ^ n46357;
  assign n48230 = n48229 ^ n46286;
  assign n48228 = n47823 ^ n47771;
  assign n48231 = n48230 ^ n48228;
  assign n48247 = n48246 ^ n48233;
  assign n48248 = ~n48235 & n48247;
  assign n48249 = n48248 ^ n48234;
  assign n48250 = n48249 ^ n48228;
  assign n48251 = ~n48231 & n48250;
  assign n48252 = n48251 ^ n48230;
  assign n48253 = n48252 ^ n48226;
  assign n48254 = n48227 & ~n48253;
  assign n48255 = n48254 ^ n48224;
  assign n48256 = n48255 ^ n48221;
  assign n48257 = n48222 & ~n48256;
  assign n48258 = n48257 ^ n48220;
  assign n48259 = n48258 ^ n48217;
  assign n48260 = ~n48218 & ~n48259;
  assign n48261 = n48260 ^ n48216;
  assign n48262 = n48261 ^ n48181;
  assign n48263 = ~n48214 & n48262;
  assign n48264 = n48263 ^ n48213;
  assign n48265 = n48264 ^ n48210;
  assign n48266 = ~n48211 & n48265;
  assign n48267 = n48266 ^ n48209;
  assign n48269 = n48268 ^ n48267;
  assign n48270 = n46878 ^ n46279;
  assign n48271 = n48270 ^ n47451;
  assign n48272 = n48271 ^ n48268;
  assign n48273 = n48269 & n48272;
  assign n48274 = n48273 ^ n48271;
  assign n48275 = n48274 ^ n48207;
  assign n48276 = n47216 ^ n47150;
  assign n48277 = n48276 ^ n46274;
  assign n48278 = n48277 ^ n48207;
  assign n48279 = n48275 & n48278;
  assign n48280 = n48279 ^ n48277;
  assign n48281 = n48280 ^ n48203;
  assign n48282 = n48206 & n48281;
  assign n48283 = n48282 ^ n48205;
  assign n48284 = n48283 ^ n48199;
  assign n48285 = n48202 & ~n48284;
  assign n48286 = n48285 ^ n48201;
  assign n48287 = n48286 ^ n48197;
  assign n48288 = n48198 & n48287;
  assign n48289 = n48288 ^ n48196;
  assign n48290 = n48289 ^ n48193;
  assign n48291 = ~n48194 & ~n48290;
  assign n48292 = n48291 ^ n48192;
  assign n48293 = n48292 ^ n48187;
  assign n48294 = n48190 & ~n48293;
  assign n48295 = n48294 ^ n48189;
  assign n48386 = n48298 ^ n48295;
  assign n48387 = n48299 & n48386;
  assign n48388 = n48387 ^ n48297;
  assign n48567 = n48392 ^ n48388;
  assign n48568 = ~n48393 & n48567;
  assign n48569 = n48568 ^ n48390;
  assign n48566 = n47905 ^ n47902;
  assign n48570 = n48569 ^ n48566;
  assign n48564 = n46619 ^ n45931;
  assign n48565 = n48564 ^ n47188;
  assign n48614 = n48566 ^ n48565;
  assign n48615 = ~n48570 & n48614;
  assign n48616 = n48615 ^ n48565;
  assign n48613 = n47908 ^ n47731;
  assign n48617 = n48616 ^ n48613;
  assign n48611 = n47361 ^ n45911;
  assign n48612 = n48611 ^ n46617;
  assign n48644 = n48613 ^ n48612;
  assign n48645 = ~n48617 & ~n48644;
  assign n48646 = n48645 ^ n48612;
  assign n48682 = n48647 ^ n48646;
  assign n48683 = n48650 & n48682;
  assign n48684 = n48683 ^ n48649;
  assign n48690 = n48689 ^ n48684;
  assign n48691 = n48690 ^ n44787;
  assign n48618 = n48617 ^ n48612;
  assign n48619 = n48618 ^ n45249;
  assign n48571 = n48570 ^ n48565;
  assign n48394 = n48393 ^ n48388;
  assign n48395 = n48394 ^ n45216;
  assign n48300 = n48299 ^ n48295;
  assign n48301 = n48300 ^ n45212;
  assign n48302 = n48292 ^ n48189;
  assign n48303 = n48302 ^ n48187;
  assign n48304 = n48303 ^ n45209;
  assign n48375 = n48289 ^ n48194;
  assign n48305 = n48286 ^ n48196;
  assign n48306 = n48305 ^ n48197;
  assign n48307 = n48306 ^ n45686;
  assign n48308 = n48283 ^ n48202;
  assign n48309 = n48308 ^ n45779;
  assign n48310 = n48280 ^ n48206;
  assign n48311 = n48310 ^ n45738;
  assign n48312 = n48277 ^ n48275;
  assign n48313 = n48312 ^ n45742;
  assign n48358 = n48271 ^ n48269;
  assign n48314 = n48264 ^ n48211;
  assign n48315 = n48314 ^ n45750;
  assign n48316 = n48261 ^ n48214;
  assign n48317 = n48316 ^ n45756;
  assign n48318 = n48258 ^ n48218;
  assign n48319 = n48318 ^ n45676;
  assign n48344 = n48255 ^ n48222;
  assign n48320 = n48252 ^ n48224;
  assign n48321 = n48320 ^ n48226;
  assign n48322 = n48321 ^ n45471;
  assign n48323 = n48249 ^ n48231;
  assign n48324 = n48323 ^ n45455;
  assign n48335 = n48333 ^ n45441;
  assign n48336 = n48334 & ~n48335;
  assign n48337 = n48336 ^ n45441;
  assign n48338 = n48337 ^ n48323;
  assign n48339 = n48324 & n48338;
  assign n48340 = n48339 ^ n45455;
  assign n48341 = n48340 ^ n48321;
  assign n48342 = n48322 & n48341;
  assign n48343 = n48342 ^ n45471;
  assign n48345 = n48344 ^ n48343;
  assign n48346 = n48344 ^ n45651;
  assign n48347 = ~n48345 & n48346;
  assign n48348 = n48347 ^ n45651;
  assign n48349 = n48348 ^ n48318;
  assign n48350 = n48319 & n48349;
  assign n48351 = n48350 ^ n45676;
  assign n48352 = n48351 ^ n48316;
  assign n48353 = n48317 & n48352;
  assign n48354 = n48353 ^ n45756;
  assign n48355 = n48354 ^ n48314;
  assign n48356 = n48315 & ~n48355;
  assign n48357 = n48356 ^ n45750;
  assign n48359 = n48358 ^ n48357;
  assign n48360 = n48358 ^ n45746;
  assign n48361 = n48359 & ~n48360;
  assign n48362 = n48361 ^ n45746;
  assign n48363 = n48362 ^ n48312;
  assign n48364 = ~n48313 & ~n48363;
  assign n48365 = n48364 ^ n45742;
  assign n48366 = n48365 ^ n48310;
  assign n48367 = ~n48311 & ~n48366;
  assign n48368 = n48367 ^ n45738;
  assign n48369 = n48368 ^ n48308;
  assign n48370 = ~n48309 & ~n48369;
  assign n48371 = n48370 ^ n45779;
  assign n48372 = n48371 ^ n48306;
  assign n48373 = ~n48307 & n48372;
  assign n48374 = n48373 ^ n45686;
  assign n48376 = n48375 ^ n48374;
  assign n48377 = n48375 ^ n45902;
  assign n48378 = n48376 & n48377;
  assign n48379 = n48378 ^ n45902;
  assign n48380 = n48379 ^ n48303;
  assign n48381 = n48304 & ~n48380;
  assign n48382 = n48381 ^ n45209;
  assign n48383 = n48382 ^ n48300;
  assign n48384 = n48301 & ~n48383;
  assign n48385 = n48384 ^ n45212;
  assign n48561 = n48394 ^ n48385;
  assign n48562 = ~n48395 & ~n48561;
  assign n48563 = n48562 ^ n45216;
  assign n48572 = n48571 ^ n48563;
  assign n48608 = n48571 ^ n45201;
  assign n48609 = ~n48572 & ~n48608;
  assign n48610 = n48609 ^ n45201;
  assign n48653 = n48618 ^ n48610;
  assign n48654 = n48619 & ~n48653;
  assign n48655 = n48654 ^ n45249;
  assign n48678 = n48655 ^ n44791;
  assign n48651 = n48650 ^ n48646;
  assign n48679 = n48655 ^ n48651;
  assign n48680 = ~n48678 & ~n48679;
  assign n48681 = n48680 ^ n44791;
  assign n48692 = n48691 ^ n48681;
  assign n48573 = n48572 ^ n45201;
  assign n48396 = n48395 ^ n48385;
  assign n48397 = n48379 ^ n48304;
  assign n48398 = n48376 ^ n45902;
  assign n48399 = n48368 ^ n48309;
  assign n48400 = n48365 ^ n48311;
  assign n48401 = n48362 ^ n48313;
  assign n48402 = n48354 ^ n45750;
  assign n48403 = n48402 ^ n48314;
  assign n48404 = n48340 ^ n48322;
  assign n48405 = n48337 ^ n48324;
  assign n48410 = n48408 & ~n48409;
  assign n48411 = n48405 & n48410;
  assign n48412 = n48404 & ~n48411;
  assign n48413 = n48345 ^ n45651;
  assign n48414 = n48412 & ~n48413;
  assign n48415 = n48348 ^ n48319;
  assign n48416 = ~n48414 & n48415;
  assign n48417 = n48351 ^ n48317;
  assign n48418 = ~n48416 & n48417;
  assign n48419 = n48403 & ~n48418;
  assign n48420 = n48359 ^ n45746;
  assign n48421 = n48419 & ~n48420;
  assign n48422 = ~n48401 & n48421;
  assign n48423 = ~n48400 & ~n48422;
  assign n48424 = n48399 & n48423;
  assign n48425 = n48371 ^ n48307;
  assign n48426 = ~n48424 & n48425;
  assign n48427 = ~n48398 & n48426;
  assign n48428 = ~n48397 & ~n48427;
  assign n48429 = n48382 ^ n48301;
  assign n48430 = ~n48428 & n48429;
  assign n48574 = n48396 & ~n48430;
  assign n48607 = n48573 & ~n48574;
  assign n48620 = n48619 ^ n48610;
  assign n48643 = n48607 & n48620;
  assign n48652 = n48651 ^ n44791;
  assign n48656 = n48655 ^ n48652;
  assign n48676 = ~n48643 & n48656;
  assign n48673 = n46594 ^ n38477;
  assign n48674 = n48673 ^ n43160;
  assign n48675 = n48674 ^ n37252;
  assign n48677 = n48676 ^ n48675;
  assign n48693 = n48692 ^ n48677;
  assign n48657 = n48656 ^ n48643;
  assign n48640 = n46491 ^ n38716;
  assign n48641 = n48640 ^ n43044;
  assign n48642 = n48641 ^ n37102;
  assign n48658 = n48657 ^ n48642;
  assign n48621 = n48620 ^ n48607;
  assign n48576 = n46501 ^ n38721;
  assign n48577 = n48576 ^ n1253;
  assign n48578 = n48577 ^ n37107;
  assign n48575 = n48574 ^ n48573;
  assign n48579 = n48578 ^ n48575;
  assign n48431 = n48430 ^ n48396;
  assign n48184 = n46506 ^ n38725;
  assign n48185 = n48184 ^ n43053;
  assign n48186 = n48185 ^ n1245;
  assign n48432 = n48431 ^ n48186;
  assign n48433 = n48429 ^ n48428;
  assign n1065 = n1064 ^ n1022;
  assign n1099 = n1098 ^ n1065;
  assign n1109 = n1108 ^ n1099;
  assign n48434 = n48433 ^ n1109;
  assign n48436 = n46513 ^ n38731;
  assign n48437 = n48436 ^ n43121;
  assign n48438 = n48437 ^ n1090;
  assign n48435 = n48427 ^ n48397;
  assign n48439 = n48438 ^ n48435;
  assign n48441 = n46518 ^ n933;
  assign n48442 = n48441 ^ n43061;
  assign n48443 = n48442 ^ n37118;
  assign n48440 = n48426 ^ n48398;
  assign n48444 = n48443 ^ n48440;
  assign n48446 = n46522 ^ n38738;
  assign n48447 = n48446 ^ n43110;
  assign n48448 = n48447 ^ n37123;
  assign n48445 = n48425 ^ n48424;
  assign n48449 = n48448 ^ n48445;
  assign n48453 = n48423 ^ n48399;
  assign n48450 = n46528 ^ n38743;
  assign n48451 = n48450 ^ n43066;
  assign n48452 = n48451 ^ n37127;
  assign n48454 = n48453 ^ n48452;
  assign n48458 = n48422 ^ n48400;
  assign n48455 = n46545 ^ n38747;
  assign n48456 = n48455 ^ n43070;
  assign n48457 = n48456 ^ n37132;
  assign n48459 = n48458 ^ n48457;
  assign n48463 = n48421 ^ n48401;
  assign n48460 = n46532 ^ n38752;
  assign n48461 = n48460 ^ n43075;
  assign n48462 = n48461 ^ n37137;
  assign n48464 = n48463 ^ n48462;
  assign n48466 = n46269 ^ n38778;
  assign n48467 = n48466 ^ n43081;
  assign n48468 = n48467 ^ n37142;
  assign n48465 = n48420 ^ n48419;
  assign n48469 = n48468 ^ n48465;
  assign n48526 = n48418 ^ n48403;
  assign n48471 = n46242 ^ n38767;
  assign n48472 = n48471 ^ n42833;
  assign n48473 = n48472 ^ n37186;
  assign n48470 = n48417 ^ n48416;
  assign n48474 = n48473 ^ n48470;
  assign n48475 = n48415 ^ n48414;
  assign n48479 = n48478 ^ n48475;
  assign n48481 = n46124 ^ n38351;
  assign n48482 = n48481 ^ n42705;
  assign n48483 = n48482 ^ n37175;
  assign n48480 = n48413 ^ n48412;
  assign n48484 = n48483 ^ n48480;
  assign n48486 = n46130 ^ n38235;
  assign n48487 = n48486 ^ n2263;
  assign n48488 = n48487 ^ n37157;
  assign n48485 = n48411 ^ n48404;
  assign n48489 = n48488 ^ n48485;
  assign n48490 = n48410 ^ n48405;
  assign n2218 = n2208 ^ n2148;
  assign n2246 = n2245 ^ n2218;
  assign n2253 = n2252 ^ n2246;
  assign n48491 = n48490 ^ n2253;
  assign n48496 = n48495 ^ n48492;
  assign n48508 = n48507 ^ n48492;
  assign n48509 = ~n48496 & n48508;
  assign n48510 = n48509 ^ n48495;
  assign n48511 = n48510 ^ n48490;
  assign n48512 = n48491 & ~n48511;
  assign n48513 = n48512 ^ n2253;
  assign n48514 = n48513 ^ n48485;
  assign n48515 = n48489 & ~n48514;
  assign n48516 = n48515 ^ n48488;
  assign n48517 = n48516 ^ n48480;
  assign n48518 = n48484 & ~n48517;
  assign n48519 = n48518 ^ n48483;
  assign n48520 = n48519 ^ n48475;
  assign n48521 = ~n48479 & n48520;
  assign n48522 = n48521 ^ n48478;
  assign n48523 = n48522 ^ n48470;
  assign n48524 = n48474 & ~n48523;
  assign n48525 = n48524 ^ n48473;
  assign n48527 = n48526 ^ n48525;
  assign n48528 = n46115 ^ n38758;
  assign n48529 = n48528 ^ n43086;
  assign n48530 = n48529 ^ n37148;
  assign n48531 = n48530 ^ n48526;
  assign n48532 = n48527 & ~n48531;
  assign n48533 = n48532 ^ n48530;
  assign n48534 = n48533 ^ n48468;
  assign n48535 = ~n48469 & ~n48534;
  assign n48536 = n48535 ^ n48465;
  assign n48537 = n48536 ^ n48463;
  assign n48538 = ~n48464 & ~n48537;
  assign n48539 = n48538 ^ n48462;
  assign n48540 = n48539 ^ n48458;
  assign n48541 = ~n48459 & n48540;
  assign n48542 = n48541 ^ n48457;
  assign n48543 = n48542 ^ n48452;
  assign n48544 = ~n48454 & ~n48543;
  assign n48545 = n48544 ^ n48453;
  assign n48546 = n48545 ^ n48445;
  assign n48547 = ~n48449 & ~n48546;
  assign n48548 = n48547 ^ n48448;
  assign n48549 = n48548 ^ n48440;
  assign n48550 = ~n48444 & n48549;
  assign n48551 = n48550 ^ n48443;
  assign n48552 = n48551 ^ n48435;
  assign n48553 = ~n48439 & n48552;
  assign n48554 = n48553 ^ n48438;
  assign n48555 = n48554 ^ n48433;
  assign n48556 = ~n48434 & n48555;
  assign n48557 = n48556 ^ n1109;
  assign n48558 = n48557 ^ n48186;
  assign n48559 = n48432 & ~n48558;
  assign n48560 = n48559 ^ n48431;
  assign n48604 = n48578 ^ n48560;
  assign n48605 = ~n48579 & ~n48604;
  assign n48606 = n48605 ^ n48575;
  assign n48622 = n48621 ^ n48606;
  assign n48601 = n46495 ^ n38815;
  assign n48602 = n48601 ^ n43048;
  assign n48603 = n48602 ^ n2303;
  assign n48637 = n48621 ^ n48603;
  assign n48638 = n48622 & n48637;
  assign n48639 = n48638 ^ n48603;
  assign n48670 = n48642 ^ n48639;
  assign n48671 = n48658 & ~n48670;
  assign n48672 = n48671 ^ n48657;
  assign n48694 = n48693 ^ n48672;
  assign n48668 = n48061 ^ n46323;
  assign n48669 = n48668 ^ n47210;
  assign n48695 = n48694 ^ n48669;
  assign n48659 = n48658 ^ n48639;
  assign n48635 = n48014 ^ n47392;
  assign n48636 = n48635 ^ n46328;
  assign n48660 = n48659 ^ n48636;
  assign n48623 = n48622 ^ n48603;
  assign n48585 = n47270 ^ n47208;
  assign n48586 = n48585 ^ n46665;
  assign n48581 = n47993 ^ n47276;
  assign n48582 = n48581 ^ n46658;
  assign n48583 = n48557 ^ n48432;
  assign n48584 = ~n48582 & n48583;
  assign n48587 = n48586 ^ n48584;
  assign n48580 = n48579 ^ n48560;
  assign n48598 = n48584 ^ n48580;
  assign n48599 = n48587 & n48598;
  assign n48600 = n48599 ^ n48586;
  assign n48624 = n48623 ^ n48600;
  assign n48596 = n47265 ^ n46672;
  assign n48597 = n48596 ^ n48004;
  assign n48632 = n48623 ^ n48597;
  assign n48633 = n48624 & n48632;
  assign n48634 = n48633 ^ n48597;
  assign n48665 = n48636 ^ n48634;
  assign n48666 = ~n48660 & ~n48665;
  assign n48667 = n48666 ^ n48659;
  assign n48747 = n48669 ^ n48667;
  assign n48748 = ~n48695 & ~n48747;
  assign n48749 = n48748 ^ n48694;
  assign n48751 = n48750 ^ n48749;
  assign n48745 = n48170 ^ n47263;
  assign n48746 = n48745 ^ n46318;
  assign n48842 = n48750 ^ n48746;
  assign n48843 = ~n48751 & ~n48842;
  assign n48844 = n48843 ^ n48746;
  assign n48845 = n48844 ^ n48840;
  assign n48846 = n48841 & ~n48845;
  assign n48847 = n48846 ^ n48838;
  assign n48848 = n48847 ^ n48835;
  assign n48849 = n48836 & n48848;
  assign n48850 = n48849 ^ n48834;
  assign n48853 = n48852 ^ n48850;
  assign n48854 = n48228 ^ n47251;
  assign n48855 = n48854 ^ n46699;
  assign n48856 = n48855 ^ n48852;
  assign n48857 = n48853 & n48856;
  assign n48858 = n48857 ^ n48855;
  assign n48773 = n48141 ^ n48113;
  assign n48859 = n48858 ^ n48773;
  assign n48860 = n47249 ^ n46310;
  assign n48861 = n48860 ^ n48226;
  assign n48862 = n48861 ^ n48773;
  assign n48863 = n48859 & ~n48862;
  assign n48864 = n48863 ^ n48861;
  assign n48865 = n48864 ^ n48829;
  assign n48866 = n48832 & n48865;
  assign n48867 = n48866 ^ n48831;
  assign n48828 = n48147 ^ n48103;
  assign n48868 = n48867 ^ n48828;
  assign n48869 = n47241 ^ n46298;
  assign n48870 = n48869 ^ n48217;
  assign n48871 = n48870 ^ n48828;
  assign n48872 = n48868 & ~n48871;
  assign n48873 = n48872 ^ n48870;
  assign n48874 = n48873 ^ n48826;
  assign n48875 = ~n48827 & n48874;
  assign n48876 = n48875 ^ n48766;
  assign n48877 = n48876 ^ n48823;
  assign n48878 = n48824 & n48877;
  assign n48879 = n48878 ^ n48822;
  assign n48760 = n48156 ^ n48088;
  assign n48880 = n48879 ^ n48760;
  assign n48881 = n48268 ^ n46277;
  assign n48882 = n48881 ^ n47228;
  assign n48883 = n48882 ^ n48760;
  assign n48884 = n48880 & n48883;
  assign n48885 = n48884 ^ n48882;
  assign n48886 = n48885 ^ n48180;
  assign n48887 = n48820 & n48886;
  assign n48888 = n48887 ^ n48819;
  assign n48889 = n48888 ^ n48816;
  assign n48890 = ~n48817 & n48889;
  assign n48891 = n48890 ^ n48815;
  assign n48894 = n48893 ^ n48891;
  assign n48958 = n48896 ^ n48894;
  assign n48959 = n48958 ^ n46289;
  assign n48960 = n48888 ^ n48817;
  assign n48961 = n48960 ^ n46294;
  assign n48962 = n48885 ^ n48819;
  assign n48963 = n48962 ^ n48180;
  assign n48964 = n48963 ^ n46300;
  assign n49008 = n48882 ^ n48880;
  assign n48965 = n48876 ^ n48824;
  assign n48966 = n48965 ^ n46357;
  assign n49000 = n48873 ^ n48827;
  assign n48967 = n48870 ^ n48868;
  assign n48968 = n48967 ^ n46255;
  assign n48969 = n48864 ^ n48832;
  assign n48970 = n48969 ^ n46072;
  assign n48989 = n48861 ^ n48859;
  assign n48971 = n48855 ^ n48853;
  assign n48972 = n48971 ^ n45689;
  assign n48973 = n48847 ^ n48836;
  assign n48974 = n48973 ^ n45696;
  assign n48975 = n48844 ^ n48841;
  assign n48976 = n48975 ^ n45700;
  assign n48752 = n48751 ^ n48746;
  assign n48753 = n48752 ^ n45704;
  assign n48661 = n48660 ^ n48634;
  assign n48662 = n48661 ^ n45710;
  assign n48625 = n48624 ^ n48597;
  assign n48626 = n48625 ^ n45714;
  assign n48589 = n48583 ^ n48582;
  assign n48590 = n45723 & ~n48589;
  assign n48591 = n48590 ^ n45718;
  assign n48588 = n48587 ^ n48580;
  assign n48593 = n48590 ^ n48588;
  assign n48594 = n48591 & n48593;
  assign n48595 = n48594 ^ n45718;
  assign n48629 = n48625 ^ n48595;
  assign n48630 = n48626 & ~n48629;
  assign n48631 = n48630 ^ n45714;
  assign n48697 = n48661 ^ n48631;
  assign n48698 = n48662 & ~n48697;
  assign n48699 = n48698 ^ n45710;
  assign n48696 = n48695 ^ n48667;
  assign n48700 = n48699 ^ n48696;
  assign n48742 = n48699 ^ n45706;
  assign n48743 = n48700 & ~n48742;
  assign n48744 = n48743 ^ n45706;
  assign n48977 = n48752 ^ n48744;
  assign n48978 = ~n48753 & n48977;
  assign n48979 = n48978 ^ n45704;
  assign n48980 = n48979 ^ n48975;
  assign n48981 = n48976 & n48980;
  assign n48982 = n48981 ^ n45700;
  assign n48983 = n48982 ^ n48973;
  assign n48984 = n48974 & ~n48983;
  assign n48985 = n48984 ^ n45696;
  assign n48986 = n48985 ^ n48971;
  assign n48987 = n48972 & n48986;
  assign n48988 = n48987 ^ n45689;
  assign n48990 = n48989 ^ n48988;
  assign n48991 = n48989 ^ n45977;
  assign n48992 = ~n48990 & n48991;
  assign n48993 = n48992 ^ n45977;
  assign n48994 = n48993 ^ n48969;
  assign n48995 = ~n48970 & n48994;
  assign n48996 = n48995 ^ n46072;
  assign n48997 = n48996 ^ n48967;
  assign n48998 = ~n48968 & n48997;
  assign n48999 = n48998 ^ n46255;
  assign n49001 = n49000 ^ n48999;
  assign n49002 = n48999 ^ n46365;
  assign n49003 = n49001 & ~n49002;
  assign n49004 = n49003 ^ n46365;
  assign n49005 = n49004 ^ n48965;
  assign n49006 = ~n48966 & n49005;
  assign n49007 = n49006 ^ n46357;
  assign n49009 = n49008 ^ n49007;
  assign n49010 = n49008 ^ n46306;
  assign n49011 = ~n49009 & n49010;
  assign n49012 = n49011 ^ n46306;
  assign n49013 = n49012 ^ n48963;
  assign n49014 = n48964 & n49013;
  assign n49015 = n49014 ^ n46300;
  assign n49016 = n49015 ^ n48960;
  assign n49017 = ~n48961 & ~n49016;
  assign n49018 = n49017 ^ n46294;
  assign n49019 = n49018 ^ n48958;
  assign n49020 = n48959 & ~n49019;
  assign n49021 = n49020 ^ n46289;
  assign n49074 = n49021 ^ n46283;
  assign n48897 = n48896 ^ n48893;
  assign n48898 = n48894 & n48897;
  assign n48899 = n48898 ^ n48896;
  assign n48810 = n48197 ^ n46865;
  assign n48811 = n48810 ^ n47216;
  assign n48955 = n48899 ^ n48811;
  assign n48812 = n48510 ^ n48491;
  assign n48956 = n48955 ^ n48812;
  assign n49075 = n49074 ^ n48956;
  assign n49076 = n49018 ^ n48959;
  assign n49077 = n49009 ^ n46306;
  assign n49078 = n49004 ^ n48966;
  assign n49079 = n49000 ^ n46365;
  assign n49080 = n49079 ^ n48999;
  assign n49081 = n48996 ^ n48968;
  assign n49082 = n48985 ^ n48972;
  assign n49083 = n48982 ^ n48974;
  assign n48754 = n48753 ^ n48744;
  assign n48592 = n48591 ^ n48588;
  assign n48627 = n48626 ^ n48595;
  assign n48628 = n48592 & ~n48627;
  assign n48663 = n48662 ^ n48631;
  assign n48664 = ~n48628 & n48663;
  assign n48701 = n48700 ^ n45706;
  assign n48755 = ~n48664 & ~n48701;
  assign n49084 = n48754 & ~n48755;
  assign n49085 = n48979 ^ n48976;
  assign n49086 = ~n49084 & n49085;
  assign n49087 = ~n49083 & n49086;
  assign n49088 = ~n49082 & n49087;
  assign n49089 = n48990 ^ n45977;
  assign n49090 = ~n49088 & ~n49089;
  assign n49091 = n48993 ^ n48970;
  assign n49092 = n49090 & n49091;
  assign n49093 = n49081 & n49092;
  assign n49094 = ~n49080 & n49093;
  assign n49095 = ~n49078 & n49094;
  assign n49096 = ~n49077 & ~n49095;
  assign n49097 = n49012 ^ n48964;
  assign n49098 = n49096 & ~n49097;
  assign n49099 = n49015 ^ n46294;
  assign n49100 = n49099 ^ n48960;
  assign n49101 = ~n49098 & n49100;
  assign n49102 = ~n49076 & ~n49101;
  assign n49103 = ~n49075 & ~n49102;
  assign n48957 = n48956 ^ n46283;
  assign n49022 = n49021 ^ n48956;
  assign n49023 = ~n48957 & n49022;
  assign n49024 = n49023 ^ n46283;
  assign n48813 = n48812 ^ n48811;
  assign n48900 = n48899 ^ n48812;
  assign n48901 = n48813 & n48900;
  assign n48902 = n48901 ^ n48811;
  assign n48808 = n48513 ^ n48489;
  assign n48806 = n48193 ^ n46878;
  assign n48807 = n48806 ^ n47461;
  assign n48809 = n48808 ^ n48807;
  assign n48953 = n48902 ^ n48809;
  assign n48954 = n48953 ^ n46279;
  assign n49073 = n49024 ^ n48954;
  assign n49187 = n49103 ^ n49073;
  assign n49191 = n49190 ^ n49187;
  assign n49193 = n46984 ^ n39157;
  assign n49194 = n49193 ^ n43674;
  assign n49195 = n49194 ^ n37920;
  assign n49192 = n49102 ^ n49075;
  assign n49196 = n49195 ^ n49192;
  assign n49198 = n47114 ^ n39163;
  assign n49199 = n49198 ^ n43666;
  assign n49200 = n49199 ^ n37925;
  assign n49197 = n49101 ^ n49076;
  assign n49201 = n49200 ^ n49197;
  assign n49203 = n46989 ^ n39168;
  assign n49204 = n49203 ^ n43544;
  assign n49205 = n49204 ^ n37929;
  assign n49202 = n49100 ^ n49098;
  assign n49206 = n49205 ^ n49202;
  assign n49208 = n46994 ^ n39279;
  assign n49209 = n49208 ^ n43549;
  assign n49210 = n49209 ^ n37989;
  assign n49207 = n49097 ^ n49096;
  assign n49211 = n49210 ^ n49207;
  assign n49213 = n46999 ^ n39173;
  assign n49214 = n49213 ^ n43554;
  assign n49215 = n49214 ^ n37935;
  assign n49212 = n49095 ^ n49077;
  assign n49216 = n49215 ^ n49212;
  assign n49218 = n47004 ^ n39178;
  assign n49219 = n49218 ^ n43559;
  assign n49220 = n49219 ^ n37978;
  assign n49217 = n49094 ^ n49078;
  assign n49221 = n49220 ^ n49217;
  assign n49223 = n47094 ^ n39183;
  assign n49224 = n49223 ^ n43564;
  assign n49225 = n49224 ^ n37940;
  assign n49222 = n49093 ^ n49080;
  assign n49226 = n49225 ^ n49222;
  assign n49230 = n49092 ^ n49081;
  assign n49227 = n47086 ^ n39188;
  assign n49228 = n49227 ^ n43643;
  assign n49229 = n49228 ^ n1931;
  assign n49231 = n49230 ^ n49229;
  assign n49268 = n49091 ^ n49090;
  assign n49260 = n49089 ^ n49088;
  assign n49235 = n49087 ^ n49082;
  assign n49232 = n47018 ^ n1685;
  assign n49233 = n49232 ^ n43627;
  assign n49234 = n49233 ^ n37949;
  assign n49236 = n49235 ^ n49234;
  assign n49238 = n47024 ^ n39199;
  assign n49239 = n49238 ^ n43574;
  assign n49240 = n49239 ^ n37399;
  assign n49237 = n49086 ^ n49083;
  assign n49241 = n49240 ^ n49237;
  assign n49242 = n49085 ^ n49084;
  assign n49246 = n49245 ^ n49242;
  assign n48756 = n48755 ^ n48754;
  assign n48738 = n47063 ^ n39210;
  assign n48739 = n48738 ^ n43579;
  assign n48740 = n48739 ^ n37364;
  assign n49247 = n48756 ^ n48740;
  assign n48703 = n47055 ^ n39236;
  assign n48704 = n48703 ^ n43584;
  assign n48705 = n48704 ^ n37369;
  assign n48702 = n48701 ^ n48664;
  assign n48706 = n48705 ^ n48702;
  assign n48727 = n48663 ^ n48628;
  assign n48719 = n47033 ^ n39218;
  assign n48720 = n48719 ^ n43598;
  assign n48721 = n48720 ^ n37379;
  assign n48712 = n47036 ^ n39221;
  assign n48713 = n48712 ^ n43593;
  assign n48714 = n48713 ^ n2579;
  assign n48707 = n48589 ^ n45723;
  assign n48708 = n47342 ^ n39440;
  assign n48709 = n48708 ^ n2468;
  assign n48710 = n48709 ^ n38048;
  assign n48711 = ~n48707 & n48710;
  assign n48715 = n48714 ^ n48711;
  assign n48716 = n48711 ^ n48592;
  assign n48717 = n48715 & ~n48716;
  assign n48718 = n48717 ^ n48714;
  assign n48722 = n48721 ^ n48718;
  assign n48723 = n48627 ^ n48592;
  assign n48724 = n48723 ^ n48718;
  assign n48725 = n48722 & ~n48724;
  assign n48726 = n48725 ^ n48721;
  assign n48728 = n48727 ^ n48726;
  assign n48729 = n47047 ^ n39214;
  assign n48730 = n48729 ^ n43589;
  assign n48731 = n48730 ^ n37373;
  assign n48732 = n48731 ^ n48727;
  assign n48733 = n48728 & ~n48732;
  assign n48734 = n48733 ^ n48731;
  assign n48735 = n48734 ^ n48702;
  assign n48736 = ~n48706 & n48735;
  assign n48737 = n48736 ^ n48705;
  assign n49248 = n48756 ^ n48737;
  assign n49249 = ~n49247 & n49248;
  assign n49250 = n49249 ^ n48740;
  assign n49251 = n49250 ^ n49242;
  assign n49252 = n49246 & ~n49251;
  assign n49253 = n49252 ^ n49245;
  assign n49254 = n49253 ^ n49237;
  assign n49255 = n49241 & ~n49254;
  assign n49256 = n49255 ^ n49240;
  assign n49257 = n49256 ^ n49235;
  assign n49258 = n49236 & ~n49257;
  assign n49259 = n49258 ^ n49234;
  assign n49261 = n49260 ^ n49259;
  assign n49262 = n47013 ^ n39256;
  assign n49263 = n49262 ^ n43568;
  assign n49264 = n49263 ^ n1803;
  assign n49265 = n49264 ^ n49260;
  assign n49266 = ~n49261 & n49265;
  assign n49267 = n49266 ^ n49264;
  assign n49269 = n49268 ^ n49267;
  assign n49270 = n47008 ^ n39193;
  assign n49271 = n49270 ^ n1811;
  assign n49272 = n49271 ^ n37944;
  assign n49273 = n49272 ^ n49268;
  assign n49274 = ~n49269 & n49273;
  assign n49275 = n49274 ^ n49272;
  assign n49276 = n49275 ^ n49230;
  assign n49277 = n49231 & ~n49276;
  assign n49278 = n49277 ^ n49229;
  assign n49279 = n49278 ^ n49222;
  assign n49280 = ~n49226 & n49279;
  assign n49281 = n49280 ^ n49225;
  assign n49282 = n49281 ^ n49217;
  assign n49283 = ~n49221 & n49282;
  assign n49284 = n49283 ^ n49220;
  assign n49285 = n49284 ^ n49212;
  assign n49286 = ~n49216 & n49285;
  assign n49287 = n49286 ^ n49215;
  assign n49288 = n49287 ^ n49207;
  assign n49289 = n49211 & ~n49288;
  assign n49290 = n49289 ^ n49210;
  assign n49291 = n49290 ^ n49202;
  assign n49292 = ~n49206 & n49291;
  assign n49293 = n49292 ^ n49205;
  assign n49294 = n49293 ^ n49197;
  assign n49295 = ~n49201 & n49294;
  assign n49296 = n49295 ^ n49200;
  assign n49297 = n49296 ^ n49192;
  assign n49298 = n49196 & ~n49297;
  assign n49299 = n49298 ^ n49195;
  assign n49300 = n49299 ^ n49187;
  assign n49301 = n49191 & ~n49300;
  assign n49302 = n49301 ^ n49190;
  assign n49025 = n49024 ^ n48953;
  assign n49026 = n48954 & ~n49025;
  assign n49027 = n49026 ^ n46279;
  assign n48903 = n48902 ^ n48808;
  assign n48904 = n48809 & ~n48903;
  assign n48905 = n48904 ^ n48807;
  assign n48803 = n48516 ^ n48483;
  assign n48804 = n48803 ^ n48480;
  assign n48801 = n47469 ^ n47150;
  assign n48802 = n48801 ^ n48187;
  assign n48805 = n48804 ^ n48802;
  assign n48951 = n48905 ^ n48805;
  assign n48952 = n48951 ^ n46274;
  assign n49105 = n49027 ^ n48952;
  assign n49104 = n49073 & n49103;
  assign n49185 = n49105 ^ n49104;
  assign n49182 = n46974 ^ n39153;
  assign n49183 = n49182 ^ n43533;
  assign n49184 = n49183 ^ n37910;
  assign n49186 = n49185 ^ n49184;
  assign n49751 = n49302 ^ n49186;
  assign n49675 = n48686 ^ n47953;
  assign n49065 = n48548 ^ n48444;
  assign n49676 = n49675 ^ n49065;
  assign n49673 = n49299 ^ n49190;
  assign n49674 = n49673 ^ n49187;
  assign n49677 = n49676 ^ n49674;
  assign n49678 = n48647 ^ n47632;
  assign n48938 = n48545 ^ n48449;
  assign n49679 = n49678 ^ n48938;
  assign n49630 = n49296 ^ n49196;
  assign n49680 = n49679 ^ n49630;
  assign n49683 = n49293 ^ n49201;
  assign n48776 = n48542 ^ n48454;
  assign n49681 = n48776 ^ n48613;
  assign n49682 = n49681 ^ n47622;
  assign n49684 = n49683 ^ n49682;
  assign n48777 = n48539 ^ n48457;
  assign n48778 = n48777 ^ n48458;
  assign n49686 = n48778 ^ n48566;
  assign n49687 = n49686 ^ n47476;
  assign n49685 = n49290 ^ n49206;
  assign n49688 = n49687 ^ n49685;
  assign n48779 = n48536 ^ n48462;
  assign n48780 = n48779 ^ n48463;
  assign n49690 = n48780 ^ n47469;
  assign n49691 = n49690 ^ n48392;
  assign n49689 = n49287 ^ n49211;
  assign n49692 = n49691 ^ n49689;
  assign n49693 = n48298 ^ n47461;
  assign n48784 = n48533 ^ n48469;
  assign n49694 = n49693 ^ n48784;
  assign n49636 = n49284 ^ n49215;
  assign n49637 = n49636 ^ n49212;
  assign n49695 = n49694 ^ n49637;
  assign n49698 = n49281 ^ n49220;
  assign n49699 = n49698 ^ n49217;
  assign n48788 = n48530 ^ n48527;
  assign n49696 = n48788 ^ n47216;
  assign n49697 = n49696 ^ n48187;
  assign n49700 = n49699 ^ n49697;
  assign n49701 = n48193 ^ n47451;
  assign n48794 = n48522 ^ n48474;
  assign n49702 = n49701 ^ n48794;
  assign n49644 = n49278 ^ n49225;
  assign n49645 = n49644 ^ n49222;
  assign n49703 = n49702 ^ n49645;
  assign n48798 = n48519 ^ n48478;
  assign n48799 = n48798 ^ n48475;
  assign n49705 = n48799 ^ n47223;
  assign n49706 = n49705 ^ n48197;
  assign n49704 = n49275 ^ n49231;
  assign n49707 = n49706 ^ n49704;
  assign n49708 = n48804 ^ n47227;
  assign n49709 = n49708 ^ n48199;
  assign n49649 = n49272 ^ n49269;
  assign n49710 = n49709 ^ n49649;
  assign n49712 = n48203 ^ n47228;
  assign n49713 = n49712 ^ n48808;
  assign n49711 = n49264 ^ n49261;
  assign n49714 = n49713 ^ n49711;
  assign n49619 = n49256 ^ n49236;
  assign n49484 = n49253 ^ n49240;
  assign n49485 = n49484 ^ n49237;
  assign n49482 = n48893 ^ n48268;
  assign n49483 = n49482 ^ n47237;
  assign n49486 = n49485 ^ n49483;
  assign n49419 = n49250 ^ n49246;
  assign n49417 = n48816 ^ n47241;
  assign n49418 = n49417 ^ n48210;
  assign n49420 = n49419 ^ n49418;
  assign n48741 = n48740 ^ n48737;
  assign n48757 = n48756 ^ n48741;
  assign n48182 = n48181 ^ n48180;
  assign n48183 = n48182 ^ n47246;
  assign n48758 = n48757 ^ n48183;
  assign n48761 = n48217 ^ n47249;
  assign n48762 = n48761 ^ n48760;
  assign n48759 = n48734 ^ n48706;
  assign n48763 = n48762 ^ n48759;
  assign n49404 = n48731 ^ n48728;
  assign n48767 = n48766 ^ n48226;
  assign n48768 = n48767 ^ n47252;
  assign n48764 = n48723 ^ n48721;
  assign n48765 = n48764 ^ n48718;
  assign n48769 = n48768 ^ n48765;
  assign n49063 = n47970 ^ n47352;
  assign n49064 = n49063 ^ n46617;
  assign n49066 = n49065 ^ n49064;
  assign n48936 = n47358 ^ n46619;
  assign n48937 = n48936 ^ n47980;
  assign n48939 = n48938 ^ n48937;
  assign n48781 = n47192 ^ n46625;
  assign n48782 = n48781 ^ n48647;
  assign n48783 = n48782 ^ n48780;
  assign n48785 = n47953 ^ n47345;
  assign n48786 = n48785 ^ n48613;
  assign n48787 = n48786 ^ n48784;
  assign n48789 = n47632 ^ n47218;
  assign n48790 = n48789 ^ n48566;
  assign n48791 = n48790 ^ n48788;
  assign n48792 = n47622 ^ n47299;
  assign n48793 = n48792 ^ n48392;
  assign n48795 = n48794 ^ n48793;
  assign n48796 = n47476 ^ n47180;
  assign n48797 = n48796 ^ n48298;
  assign n48800 = n48799 ^ n48797;
  assign n48906 = n48905 ^ n48804;
  assign n48907 = ~n48805 & ~n48906;
  assign n48908 = n48907 ^ n48802;
  assign n48909 = n48908 ^ n48797;
  assign n48910 = n48800 & ~n48909;
  assign n48911 = n48910 ^ n48799;
  assign n48912 = n48911 ^ n48794;
  assign n48913 = n48795 & n48912;
  assign n48914 = n48913 ^ n48793;
  assign n48915 = n48914 ^ n48788;
  assign n48916 = ~n48791 & n48915;
  assign n48917 = n48916 ^ n48790;
  assign n48918 = n48917 ^ n48784;
  assign n48919 = ~n48787 & n48918;
  assign n48920 = n48919 ^ n48786;
  assign n48921 = n48920 ^ n48782;
  assign n48922 = ~n48783 & n48921;
  assign n48923 = n48922 ^ n48780;
  assign n48924 = n48923 ^ n48778;
  assign n48925 = n47188 ^ n46630;
  assign n48926 = n48925 ^ n48686;
  assign n48927 = n48926 ^ n48778;
  assign n48928 = n48924 & ~n48927;
  assign n48929 = n48928 ^ n48926;
  assign n48930 = n48929 ^ n48776;
  assign n48931 = n47974 ^ n47361;
  assign n48932 = n48931 ^ n46634;
  assign n48933 = n48932 ^ n48776;
  assign n48934 = n48930 & ~n48933;
  assign n48935 = n48934 ^ n48932;
  assign n49060 = n48937 ^ n48935;
  assign n49061 = n48939 & ~n49060;
  assign n49062 = n49061 ^ n48938;
  assign n49067 = n49066 ^ n49062;
  assign n48941 = n48932 ^ n48930;
  assign n48942 = n48941 ^ n45913;
  assign n48943 = n48926 ^ n48924;
  assign n48944 = n48943 ^ n45924;
  assign n49040 = n48917 ^ n48787;
  assign n48945 = n48914 ^ n48791;
  assign n48946 = n48945 ^ n46583;
  assign n48947 = n48911 ^ n48795;
  assign n48948 = n48947 ^ n46481;
  assign n48949 = n48908 ^ n48800;
  assign n48950 = n48949 ^ n45685;
  assign n49028 = n49027 ^ n48951;
  assign n49029 = ~n48952 & n49028;
  assign n49030 = n49029 ^ n46274;
  assign n49031 = n49030 ^ n48949;
  assign n49032 = ~n48950 & n49031;
  assign n49033 = n49032 ^ n45685;
  assign n49034 = n49033 ^ n48947;
  assign n49035 = ~n48948 & n49034;
  assign n49036 = n49035 ^ n46481;
  assign n49037 = n49036 ^ n48945;
  assign n49038 = n48946 & n49037;
  assign n49039 = n49038 ^ n46583;
  assign n49041 = n49040 ^ n49039;
  assign n49042 = n49040 ^ n46605;
  assign n49043 = ~n49041 & ~n49042;
  assign n49044 = n49043 ^ n46605;
  assign n49045 = n49044 ^ n45921;
  assign n49046 = n48920 ^ n48783;
  assign n49047 = n49046 ^ n49044;
  assign n49048 = n49045 & n49047;
  assign n49049 = n49048 ^ n45921;
  assign n49050 = n49049 ^ n48943;
  assign n49051 = ~n48944 & n49050;
  assign n49052 = n49051 ^ n45924;
  assign n49053 = n49052 ^ n48941;
  assign n49054 = ~n48942 & n49053;
  assign n49055 = n49054 ^ n45913;
  assign n48940 = n48939 ^ n48935;
  assign n49056 = n49055 ^ n48940;
  assign n49057 = n49055 ^ n45931;
  assign n49058 = ~n49056 & n49057;
  assign n49059 = n49058 ^ n45931;
  assign n49068 = n49067 ^ n49059;
  assign n49069 = n49068 ^ n45911;
  assign n49070 = n48940 ^ n45931;
  assign n49071 = n49070 ^ n49055;
  assign n49072 = n49052 ^ n48942;
  assign n49106 = n49104 & ~n49105;
  assign n49107 = n49030 ^ n48950;
  assign n49108 = ~n49106 & n49107;
  assign n49109 = n49033 ^ n46481;
  assign n49110 = n49109 ^ n48947;
  assign n49111 = n49108 & n49110;
  assign n49112 = n49036 ^ n46583;
  assign n49113 = n49112 ^ n48945;
  assign n49114 = ~n49111 & n49113;
  assign n49115 = n49041 ^ n46605;
  assign n49116 = n49114 & n49115;
  assign n49117 = n49046 ^ n49045;
  assign n49118 = ~n49116 & n49117;
  assign n49119 = n49049 ^ n48944;
  assign n49120 = ~n49118 & ~n49119;
  assign n49121 = n49072 & ~n49120;
  assign n49122 = n49071 & ~n49121;
  assign n49123 = ~n49069 & n49122;
  assign n49131 = n49065 ^ n49062;
  assign n49132 = n49066 & n49131;
  assign n49133 = n49132 ^ n49064;
  assign n49128 = n47964 ^ n46647;
  assign n49129 = n49128 ^ n47283;
  assign n49127 = n48551 ^ n48439;
  assign n49130 = n49129 ^ n49127;
  assign n49134 = n49133 ^ n49130;
  assign n49135 = n49134 ^ n45732;
  assign n49124 = n49067 ^ n45911;
  assign n49125 = ~n49068 & ~n49124;
  assign n49126 = n49125 ^ n45911;
  assign n49136 = n49135 ^ n49126;
  assign n49355 = ~n49123 & ~n49136;
  assign n49352 = n47289 ^ n39542;
  assign n49353 = n49352 ^ n43877;
  assign n49354 = n49353 ^ n2460;
  assign n49356 = n49355 ^ n49354;
  assign n49348 = n47279 ^ n46331;
  assign n49349 = n49348 ^ n47960;
  assign n49345 = n48554 ^ n1109;
  assign n49346 = n49345 ^ n48433;
  assign n49342 = n49133 ^ n49129;
  assign n49343 = ~n49130 & n49342;
  assign n49344 = n49343 ^ n49133;
  assign n49347 = n49346 ^ n49344;
  assign n49350 = n49349 ^ n49347;
  assign n49338 = n49134 ^ n49126;
  assign n49339 = ~n49135 & ~n49338;
  assign n49340 = n49339 ^ n45732;
  assign n49341 = n49340 ^ n45730;
  assign n49351 = n49350 ^ n49341;
  assign n49357 = n49356 ^ n49351;
  assign n49138 = n47322 ^ n2345;
  assign n49139 = n49138 ^ n43849;
  assign n49140 = n49139 ^ n37874;
  assign n49137 = n49136 ^ n49123;
  assign n49141 = n49140 ^ n49137;
  assign n49145 = n49122 ^ n49069;
  assign n49142 = n47169 ^ n39549;
  assign n49143 = n49142 ^ n1408;
  assign n49144 = n49143 ^ n37878;
  assign n49146 = n49145 ^ n49144;
  assign n49327 = n49121 ^ n49071;
  assign n49150 = n49120 ^ n49072;
  assign n49147 = n46939 ^ n1198;
  assign n49148 = n49147 ^ n43725;
  assign n49149 = n49148 ^ n1382;
  assign n49151 = n49150 ^ n49149;
  assign n49153 = n46944 ^ n1180;
  assign n49154 = n49153 ^ n43509;
  assign n49155 = n49154 ^ n38027;
  assign n49152 = n49119 ^ n49118;
  assign n49156 = n49155 ^ n49152;
  assign n49157 = n49117 ^ n49116;
  assign n49161 = n49160 ^ n49157;
  assign n49163 = n46954 ^ n39138;
  assign n49164 = n49163 ^ n43519;
  assign n49165 = n49164 ^ n37892;
  assign n49162 = n49115 ^ n49114;
  assign n49166 = n49165 ^ n49162;
  assign n49168 = n46959 ^ n39142;
  assign n49169 = n49168 ^ n43694;
  assign n49170 = n49169 ^ n37898;
  assign n49167 = n49113 ^ n49111;
  assign n49171 = n49170 ^ n49167;
  assign n49173 = n46964 ^ n39148;
  assign n49174 = n49173 ^ n43524;
  assign n49175 = n49174 ^ n752;
  assign n49172 = n49110 ^ n49108;
  assign n49176 = n49175 ^ n49172;
  assign n49178 = n46969 ^ n39307;
  assign n49179 = n49178 ^ n43529;
  assign n49180 = n49179 ^ n37905;
  assign n49177 = n49107 ^ n49106;
  assign n49181 = n49180 ^ n49177;
  assign n49303 = n49302 ^ n49184;
  assign n49304 = ~n49186 & ~n49303;
  assign n49305 = n49304 ^ n49185;
  assign n49306 = n49305 ^ n49177;
  assign n49307 = n49181 & n49306;
  assign n49308 = n49307 ^ n49180;
  assign n49309 = n49308 ^ n49172;
  assign n49310 = ~n49176 & n49309;
  assign n49311 = n49310 ^ n49175;
  assign n49312 = n49311 ^ n49167;
  assign n49313 = ~n49171 & n49312;
  assign n49314 = n49313 ^ n49170;
  assign n49315 = n49314 ^ n49162;
  assign n49316 = n49166 & ~n49315;
  assign n49317 = n49316 ^ n49165;
  assign n49318 = n49317 ^ n49157;
  assign n49319 = n49161 & ~n49318;
  assign n49320 = n49319 ^ n49160;
  assign n49321 = n49320 ^ n49152;
  assign n49322 = n49156 & ~n49321;
  assign n49323 = n49322 ^ n49155;
  assign n49324 = n49323 ^ n49150;
  assign n49325 = n49151 & ~n49324;
  assign n49326 = n49325 ^ n49149;
  assign n49328 = n49327 ^ n49326;
  assign n1363 = n1353 ^ n1290;
  assign n1391 = n1390 ^ n1363;
  assign n1398 = n1397 ^ n1391;
  assign n49329 = n49327 ^ n1398;
  assign n49330 = n49328 & ~n49329;
  assign n49331 = n49330 ^ n1398;
  assign n49332 = n49331 ^ n49145;
  assign n49333 = ~n49146 & n49332;
  assign n49334 = n49333 ^ n49144;
  assign n49335 = n49334 ^ n49137;
  assign n49336 = ~n49141 & n49335;
  assign n49337 = n49336 ^ n49140;
  assign n49358 = n49357 ^ n49337;
  assign n48774 = n48773 ^ n48240;
  assign n48775 = n48774 ^ n47210;
  assign n49359 = n49358 ^ n48775;
  assign n49362 = n49334 ^ n49141;
  assign n49360 = n48170 ^ n47392;
  assign n49361 = n49360 ^ n48852;
  assign n49363 = n49362 ^ n49361;
  assign n49376 = n48835 ^ n48061;
  assign n49377 = n49376 ^ n47265;
  assign n49366 = n49323 ^ n49149;
  assign n49367 = n49366 ^ n49150;
  assign n49368 = n48004 ^ n47276;
  assign n49369 = n49368 ^ n48750;
  assign n49370 = n49367 & ~n49369;
  assign n49364 = n48840 ^ n48014;
  assign n49365 = n49364 ^ n47270;
  assign n49371 = n49370 ^ n49365;
  assign n49372 = n49328 ^ n1398;
  assign n49373 = n49372 ^ n49365;
  assign n49374 = ~n49371 & ~n49373;
  assign n49375 = n49374 ^ n49370;
  assign n49378 = n49377 ^ n49375;
  assign n49379 = n49331 ^ n49146;
  assign n49380 = n49379 ^ n49375;
  assign n49381 = n49378 & n49380;
  assign n49382 = n49381 ^ n49377;
  assign n49383 = n49382 ^ n49362;
  assign n49384 = ~n49363 & n49383;
  assign n49385 = n49384 ^ n49361;
  assign n49386 = n49385 ^ n48775;
  assign n49387 = ~n49359 & n49386;
  assign n49388 = n49387 ^ n49358;
  assign n48772 = n48710 ^ n48707;
  assign n49389 = n49388 ^ n48772;
  assign n49390 = n48234 ^ n47263;
  assign n49391 = n49390 ^ n48829;
  assign n49392 = n49391 ^ n48772;
  assign n49393 = n49389 & ~n49392;
  assign n49394 = n49393 ^ n49391;
  assign n48770 = n48714 ^ n48592;
  assign n48771 = n48770 ^ n48711;
  assign n49395 = n49394 ^ n48771;
  assign n49396 = n48228 ^ n47256;
  assign n49397 = n49396 ^ n48828;
  assign n49398 = n49397 ^ n48771;
  assign n49399 = ~n49395 & ~n49398;
  assign n49400 = n49399 ^ n49397;
  assign n49401 = n49400 ^ n48765;
  assign n49402 = ~n48769 & n49401;
  assign n49403 = n49402 ^ n48768;
  assign n49405 = n49404 ^ n49403;
  assign n49406 = n48221 ^ n47251;
  assign n49407 = n49406 ^ n48823;
  assign n49408 = n49407 ^ n49404;
  assign n49409 = ~n49405 & ~n49408;
  assign n49410 = n49409 ^ n49407;
  assign n49411 = n49410 ^ n48759;
  assign n49412 = ~n48763 & n49411;
  assign n49413 = n49412 ^ n48762;
  assign n49414 = n49413 ^ n48757;
  assign n49415 = ~n48758 & n49414;
  assign n49416 = n49415 ^ n48183;
  assign n49479 = n49418 ^ n49416;
  assign n49480 = n49420 & ~n49479;
  assign n49481 = n49480 ^ n49419;
  assign n49616 = n49485 ^ n49481;
  assign n49617 = n49486 & ~n49616;
  assign n49618 = n49617 ^ n49483;
  assign n49620 = n49619 ^ n49618;
  assign n49614 = n48812 ^ n47233;
  assign n49615 = n49614 ^ n48207;
  assign n49715 = n49619 ^ n49615;
  assign n49716 = ~n49620 & n49715;
  assign n49717 = n49716 ^ n49615;
  assign n49718 = n49717 ^ n49711;
  assign n49719 = n49714 & ~n49718;
  assign n49720 = n49719 ^ n49713;
  assign n49721 = n49720 ^ n49649;
  assign n49722 = ~n49710 & ~n49721;
  assign n49723 = n49722 ^ n49709;
  assign n49724 = n49723 ^ n49704;
  assign n49725 = ~n49707 & n49724;
  assign n49726 = n49725 ^ n49706;
  assign n49727 = n49726 ^ n49702;
  assign n49728 = ~n49703 & n49727;
  assign n49729 = n49728 ^ n49645;
  assign n49730 = n49729 ^ n49699;
  assign n49731 = ~n49700 & ~n49730;
  assign n49732 = n49731 ^ n49697;
  assign n49733 = n49732 ^ n49637;
  assign n49734 = ~n49695 & n49733;
  assign n49735 = n49734 ^ n49694;
  assign n49736 = n49735 ^ n49689;
  assign n49737 = ~n49692 & ~n49736;
  assign n49738 = n49737 ^ n49691;
  assign n49739 = n49738 ^ n49685;
  assign n49740 = ~n49688 & ~n49739;
  assign n49741 = n49740 ^ n49687;
  assign n49742 = n49741 ^ n49683;
  assign n49743 = n49684 & n49742;
  assign n49744 = n49743 ^ n49682;
  assign n49745 = n49744 ^ n49630;
  assign n49746 = n49680 & n49745;
  assign n49747 = n49746 ^ n49679;
  assign n49748 = n49747 ^ n49676;
  assign n49749 = ~n49677 & n49748;
  assign n49750 = n49749 ^ n49674;
  assign n49752 = n49751 ^ n49750;
  assign n49671 = n47974 ^ n47192;
  assign n49672 = n49671 ^ n49127;
  assign n49824 = n49751 ^ n49672;
  assign n49825 = n49752 & n49824;
  assign n49826 = n49825 ^ n49672;
  assign n49822 = n49305 ^ n49180;
  assign n49823 = n49822 ^ n49177;
  assign n49827 = n49826 ^ n49823;
  assign n49820 = n49346 ^ n47188;
  assign n49821 = n49820 ^ n47980;
  assign n49828 = n49827 ^ n49821;
  assign n49829 = n49828 ^ n46630;
  assign n49753 = n49752 ^ n49672;
  assign n49754 = n49753 ^ n46625;
  assign n49812 = n49747 ^ n49677;
  assign n49755 = n49744 ^ n49680;
  assign n49756 = n49755 ^ n47218;
  assign n49757 = n49741 ^ n49682;
  assign n49758 = n49757 ^ n49683;
  assign n49759 = n49758 ^ n47299;
  assign n49760 = n49738 ^ n49687;
  assign n49761 = n49760 ^ n49685;
  assign n49762 = n49761 ^ n47180;
  assign n49763 = n49735 ^ n49691;
  assign n49764 = n49763 ^ n49689;
  assign n49765 = n49764 ^ n47150;
  assign n49766 = n49732 ^ n49695;
  assign n49767 = n49766 ^ n46878;
  assign n49768 = n49729 ^ n49700;
  assign n49769 = n49768 ^ n46865;
  assign n49770 = n49726 ^ n49703;
  assign n49771 = n49770 ^ n46732;
  assign n49772 = n49723 ^ n49707;
  assign n49773 = n49772 ^ n46270;
  assign n49774 = n49720 ^ n49709;
  assign n49775 = n49774 ^ n49649;
  assign n49776 = n49775 ^ n46272;
  assign n49777 = n49717 ^ n49714;
  assign n49778 = n49777 ^ n46277;
  assign n49621 = n49620 ^ n49615;
  assign n49622 = n49621 ^ n46286;
  assign n49487 = n49486 ^ n49481;
  assign n49488 = n49487 ^ n46291;
  assign n49421 = n49420 ^ n49416;
  assign n49422 = n49421 ^ n46298;
  assign n49423 = n49413 ^ n48758;
  assign n49424 = n49423 ^ n46303;
  assign n49425 = n49410 ^ n48763;
  assign n49426 = n49425 ^ n46310;
  assign n49465 = n49407 ^ n49405;
  assign n49460 = n49400 ^ n48769;
  assign n49427 = n49397 ^ n49395;
  assign n49428 = n49427 ^ n46314;
  assign n49429 = n49391 ^ n49389;
  assign n49430 = n49429 ^ n46318;
  assign n49431 = n49385 ^ n49359;
  assign n49432 = n49431 ^ n46323;
  assign n49433 = n49382 ^ n49361;
  assign n49434 = n49433 ^ n49362;
  assign n49435 = n49434 ^ n46328;
  assign n49436 = n49369 ^ n49367;
  assign n49437 = ~n46658 & ~n49436;
  assign n49438 = n49437 ^ n46665;
  assign n49439 = n49372 ^ n49371;
  assign n49440 = n49439 ^ n49437;
  assign n49441 = ~n49438 & ~n49440;
  assign n49442 = n49441 ^ n46665;
  assign n49443 = n49442 ^ n46672;
  assign n49444 = n49379 ^ n49378;
  assign n49445 = n49444 ^ n49442;
  assign n49446 = ~n49443 & ~n49445;
  assign n49447 = n49446 ^ n46672;
  assign n49448 = n49447 ^ n49434;
  assign n49449 = n49435 & n49448;
  assign n49450 = n49449 ^ n46328;
  assign n49451 = n49450 ^ n49431;
  assign n49452 = n49432 & ~n49451;
  assign n49453 = n49452 ^ n46323;
  assign n49454 = n49453 ^ n49429;
  assign n49455 = ~n49430 & ~n49454;
  assign n49456 = n49455 ^ n46318;
  assign n49457 = n49456 ^ n49427;
  assign n49458 = n49428 & n49457;
  assign n49459 = n49458 ^ n46314;
  assign n49461 = n49460 ^ n49459;
  assign n49462 = n49460 ^ n46691;
  assign n49463 = n49461 & ~n49462;
  assign n49464 = n49463 ^ n46691;
  assign n49466 = n49465 ^ n49464;
  assign n49467 = n49465 ^ n46699;
  assign n49468 = n49466 & ~n49467;
  assign n49469 = n49468 ^ n46699;
  assign n49470 = n49469 ^ n49425;
  assign n49471 = n49426 & ~n49470;
  assign n49472 = n49471 ^ n46310;
  assign n49473 = n49472 ^ n49423;
  assign n49474 = n49424 & ~n49473;
  assign n49475 = n49474 ^ n46303;
  assign n49476 = n49475 ^ n49421;
  assign n49477 = n49422 & n49476;
  assign n49478 = n49477 ^ n46298;
  assign n49611 = n49487 ^ n49478;
  assign n49612 = ~n49488 & ~n49611;
  assign n49613 = n49612 ^ n46291;
  assign n49779 = n49621 ^ n49613;
  assign n49780 = ~n49622 & n49779;
  assign n49781 = n49780 ^ n46286;
  assign n49782 = n49781 ^ n49777;
  assign n49783 = ~n49778 & n49782;
  assign n49784 = n49783 ^ n46277;
  assign n49785 = n49784 ^ n49775;
  assign n49786 = ~n49776 & ~n49785;
  assign n49787 = n49786 ^ n46272;
  assign n49788 = n49787 ^ n49772;
  assign n49789 = ~n49773 & ~n49788;
  assign n49790 = n49789 ^ n46270;
  assign n49791 = n49790 ^ n49770;
  assign n49792 = n49771 & n49791;
  assign n49793 = n49792 ^ n46732;
  assign n49794 = n49793 ^ n49768;
  assign n49795 = n49769 & ~n49794;
  assign n49796 = n49795 ^ n46865;
  assign n49797 = n49796 ^ n49766;
  assign n49798 = n49767 & n49797;
  assign n49799 = n49798 ^ n46878;
  assign n49800 = n49799 ^ n49764;
  assign n49801 = ~n49765 & ~n49800;
  assign n49802 = n49801 ^ n47150;
  assign n49803 = n49802 ^ n49761;
  assign n49804 = n49762 & ~n49803;
  assign n49805 = n49804 ^ n47180;
  assign n49806 = n49805 ^ n49758;
  assign n49807 = ~n49759 & ~n49806;
  assign n49808 = n49807 ^ n47299;
  assign n49809 = n49808 ^ n49755;
  assign n49810 = ~n49756 & ~n49809;
  assign n49811 = n49810 ^ n47218;
  assign n49813 = n49812 ^ n49811;
  assign n49814 = n49812 ^ n47345;
  assign n49815 = n49813 & n49814;
  assign n49816 = n49815 ^ n47345;
  assign n49817 = n49816 ^ n49753;
  assign n49818 = ~n49754 & n49817;
  assign n49819 = n49818 ^ n46625;
  assign n49830 = n49829 ^ n49819;
  assign n49831 = n49813 ^ n47345;
  assign n49832 = n49802 ^ n47180;
  assign n49833 = n49832 ^ n49761;
  assign n49834 = n49799 ^ n49765;
  assign n49835 = n49796 ^ n49767;
  assign n49489 = n49488 ^ n49478;
  assign n49490 = n49466 ^ n46699;
  assign n49491 = n49461 ^ n46691;
  assign n49492 = n49456 ^ n46314;
  assign n49493 = n49492 ^ n49427;
  assign n49494 = n49453 ^ n49430;
  assign n49495 = n49447 ^ n49435;
  assign n49496 = n49439 ^ n49438;
  assign n49497 = n49444 ^ n49443;
  assign n49498 = n49496 & ~n49497;
  assign n49499 = n49495 & ~n49498;
  assign n49500 = n49450 ^ n49432;
  assign n49501 = ~n49499 & n49500;
  assign n49502 = n49494 & ~n49501;
  assign n49503 = ~n49493 & ~n49502;
  assign n49504 = ~n49491 & n49503;
  assign n49505 = ~n49490 & n49504;
  assign n49506 = n49469 ^ n49426;
  assign n49507 = ~n49505 & ~n49506;
  assign n49508 = n49472 ^ n49424;
  assign n49509 = n49507 & ~n49508;
  assign n49510 = n49475 ^ n46298;
  assign n49511 = n49510 ^ n49421;
  assign n49512 = n49509 & ~n49511;
  assign n49610 = ~n49489 & n49512;
  assign n49623 = n49622 ^ n49613;
  assign n49836 = n49610 & n49623;
  assign n49837 = n49781 ^ n46277;
  assign n49838 = n49837 ^ n49777;
  assign n49839 = ~n49836 & ~n49838;
  assign n49840 = n49784 ^ n49776;
  assign n49841 = n49839 & ~n49840;
  assign n49842 = n49787 ^ n49773;
  assign n49843 = ~n49841 & ~n49842;
  assign n49844 = n49790 ^ n49771;
  assign n49845 = ~n49843 & n49844;
  assign n49846 = n49793 ^ n49769;
  assign n49847 = ~n49845 & n49846;
  assign n49848 = n49835 & n49847;
  assign n49849 = n49834 & n49848;
  assign n49850 = ~n49833 & ~n49849;
  assign n49851 = n49805 ^ n49759;
  assign n49852 = n49850 & n49851;
  assign n49853 = n49808 ^ n49756;
  assign n49854 = ~n49852 & n49853;
  assign n49855 = n49831 & n49854;
  assign n49856 = n49816 ^ n46625;
  assign n49857 = n49856 ^ n49753;
  assign n49858 = ~n49855 & ~n49857;
  assign n49979 = n49830 & ~n49858;
  assign n49974 = n48583 ^ n47361;
  assign n49975 = n49974 ^ n47970;
  assign n49973 = n49308 ^ n49176;
  assign n49976 = n49975 ^ n49973;
  assign n49970 = n49823 ^ n49821;
  assign n49971 = ~n49827 & ~n49970;
  assign n49972 = n49971 ^ n49821;
  assign n49977 = n49976 ^ n49972;
  assign n49966 = n49828 ^ n49819;
  assign n49967 = ~n49829 & n49966;
  assign n49968 = n49967 ^ n46630;
  assign n49969 = n49968 ^ n46634;
  assign n49978 = n49977 ^ n49969;
  assign n49980 = n49979 ^ n49978;
  assign n49860 = n47725 ^ n40271;
  assign n49861 = n49860 ^ n44448;
  assign n49862 = n49861 ^ n1064;
  assign n49859 = n49858 ^ n49830;
  assign n49863 = n49862 ^ n49859;
  assign n49865 = n47730 ^ n40250;
  assign n49866 = n49865 ^ n941;
  assign n49867 = n49866 ^ n38731;
  assign n49864 = n49857 ^ n49855;
  assign n49868 = n49867 ^ n49864;
  assign n49872 = n49854 ^ n49831;
  assign n49869 = n47905 ^ n40260;
  assign n49870 = n49869 ^ n44266;
  assign n49871 = n49870 ^ n933;
  assign n49873 = n49872 ^ n49871;
  assign n49875 = n47735 ^ n809;
  assign n49876 = n49875 ^ n44271;
  assign n49877 = n49876 ^ n38738;
  assign n49874 = n49853 ^ n49852;
  assign n49878 = n49877 ^ n49874;
  assign n49880 = n47740 ^ n39843;
  assign n49881 = n49880 ^ n44276;
  assign n49882 = n49881 ^ n38743;
  assign n49879 = n49851 ^ n49850;
  assign n49883 = n49882 ^ n49879;
  assign n49885 = n47891 ^ n39999;
  assign n49886 = n49885 ^ n44280;
  assign n49887 = n49886 ^ n38747;
  assign n49884 = n49849 ^ n49833;
  assign n49888 = n49887 ^ n49884;
  assign n49890 = n47883 ^ n39848;
  assign n49891 = n49890 ^ n44425;
  assign n49892 = n49891 ^ n38752;
  assign n49889 = n49848 ^ n49834;
  assign n49893 = n49892 ^ n49889;
  assign n49897 = n49847 ^ n49835;
  assign n49894 = n47875 ^ n39988;
  assign n49895 = n49894 ^ n44285;
  assign n49896 = n49895 ^ n38778;
  assign n49898 = n49897 ^ n49896;
  assign n49900 = n47867 ^ n39853;
  assign n49901 = n49900 ^ n44291;
  assign n49902 = n49901 ^ n38758;
  assign n49899 = n49846 ^ n49845;
  assign n49903 = n49902 ^ n49899;
  assign n49905 = n47859 ^ n39857;
  assign n49906 = n49905 ^ n44296;
  assign n49907 = n49906 ^ n38767;
  assign n49904 = n49844 ^ n49843;
  assign n49908 = n49907 ^ n49904;
  assign n49910 = n47745 ^ n39863;
  assign n49911 = n49910 ^ n44301;
  assign n49912 = n49911 ^ n38374;
  assign n49909 = n49842 ^ n49841;
  assign n49913 = n49912 ^ n49909;
  assign n49914 = n49840 ^ n49839;
  assign n49918 = n49917 ^ n49914;
  assign n49922 = n49838 ^ n49836;
  assign n49625 = n47842 ^ n39965;
  assign n49626 = n49625 ^ n44313;
  assign n49627 = n49626 ^ n2208;
  assign n49624 = n49623 ^ n49610;
  assign n49628 = n49627 ^ n49624;
  assign n49513 = n49512 ^ n49489;
  assign n2022 = n2021 ^ n1976;
  assign n2056 = n2055 ^ n2022;
  assign n2066 = n2065 ^ n2056;
  assign n49514 = n49513 ^ n2066;
  assign n49516 = n47759 ^ n39879;
  assign n49517 = n49516 ^ n44320;
  assign n49518 = n49517 ^ n2047;
  assign n49515 = n49511 ^ n49509;
  assign n49519 = n49518 ^ n49515;
  assign n49596 = n47765 ^ n1881;
  assign n49597 = n49596 ^ n44390;
  assign n49598 = n49597 ^ n38244;
  assign n49521 = n47770 ^ n39886;
  assign n49522 = n49521 ^ n44382;
  assign n49523 = n49522 ^ n38310;
  assign n49520 = n49506 ^ n49505;
  assign n49524 = n49523 ^ n49520;
  assign n49525 = n49504 ^ n49490;
  assign n49529 = n49528 ^ n49525;
  assign n49531 = n47779 ^ n39897;
  assign n49532 = n49531 ^ n44325;
  assign n49533 = n49532 ^ n38254;
  assign n49530 = n49503 ^ n49491;
  assign n49534 = n49533 ^ n49530;
  assign n49536 = n47785 ^ n39902;
  assign n49537 = n49536 ^ n44363;
  assign n49538 = n49537 ^ n38259;
  assign n49535 = n49502 ^ n49493;
  assign n49539 = n49538 ^ n49535;
  assign n49576 = n49501 ^ n49494;
  assign n49541 = n47790 ^ n39933;
  assign n49542 = n49541 ^ n44335;
  assign n49543 = n49542 ^ n38290;
  assign n49540 = n49500 ^ n49499;
  assign n49544 = n49543 ^ n49540;
  assign n49565 = n49498 ^ n49495;
  assign n49557 = n49497 ^ n49496;
  assign n49550 = n47206 ^ n39915;
  assign n49551 = n49550 ^ n43752;
  assign n49552 = n49551 ^ n38272;
  assign n49545 = n47942 ^ n2532;
  assign n49546 = n49545 ^ n44520;
  assign n49547 = n49546 ^ n38827;
  assign n49548 = n49436 ^ n46658;
  assign n49549 = n49547 & n49548;
  assign n49553 = n49552 ^ n49549;
  assign n49554 = n49549 ^ n49496;
  assign n49555 = n49553 & ~n49554;
  assign n49556 = n49555 ^ n49552;
  assign n49558 = n49557 ^ n49556;
  assign n49559 = n39920 ^ n2621;
  assign n49560 = n49559 ^ n44345;
  assign n49561 = n49560 ^ n38277;
  assign n49562 = n49561 ^ n49556;
  assign n49563 = ~n49558 & n49562;
  assign n49564 = n49563 ^ n49561;
  assign n49566 = n49565 ^ n49564;
  assign n49567 = n47798 ^ n39911;
  assign n49568 = n49567 ^ n44340;
  assign n49569 = n49568 ^ n38268;
  assign n49570 = n49569 ^ n49564;
  assign n49571 = n49566 & n49570;
  assign n49572 = n49571 ^ n49569;
  assign n49573 = n49572 ^ n49540;
  assign n49574 = n49544 & ~n49573;
  assign n49575 = n49574 ^ n49543;
  assign n49577 = n49576 ^ n49575;
  assign n49578 = n47811 ^ n39907;
  assign n49579 = n49578 ^ n44330;
  assign n49580 = n49579 ^ n38263;
  assign n49581 = n49580 ^ n49576;
  assign n49582 = n49577 & ~n49581;
  assign n49583 = n49582 ^ n49580;
  assign n49584 = n49583 ^ n49535;
  assign n49585 = ~n49539 & n49584;
  assign n49586 = n49585 ^ n49538;
  assign n49587 = n49586 ^ n49530;
  assign n49588 = n49534 & ~n49587;
  assign n49589 = n49588 ^ n49533;
  assign n49590 = n49589 ^ n49525;
  assign n49591 = n49529 & ~n49590;
  assign n49592 = n49591 ^ n49528;
  assign n49593 = n49592 ^ n49520;
  assign n49594 = n49524 & ~n49593;
  assign n49595 = n49594 ^ n49523;
  assign n49599 = n49598 ^ n49595;
  assign n49600 = n49508 ^ n49507;
  assign n49601 = n49600 ^ n49595;
  assign n49602 = n49599 & n49601;
  assign n49603 = n49602 ^ n49598;
  assign n49604 = n49603 ^ n49515;
  assign n49605 = ~n49519 & n49604;
  assign n49606 = n49605 ^ n49518;
  assign n49607 = n49606 ^ n49513;
  assign n49608 = ~n49514 & n49607;
  assign n49609 = n49608 ^ n2066;
  assign n49919 = n49624 ^ n49609;
  assign n49920 = n49628 & ~n49919;
  assign n49921 = n49920 ^ n49627;
  assign n49923 = n49922 ^ n49921;
  assign n49924 = n47755 ^ n39873;
  assign n49925 = n49924 ^ n2216;
  assign n49926 = n49925 ^ n38235;
  assign n49927 = n49926 ^ n49922;
  assign n49928 = n49923 & ~n49927;
  assign n49929 = n49928 ^ n49926;
  assign n49930 = n49929 ^ n49914;
  assign n49931 = n49918 & ~n49930;
  assign n49932 = n49931 ^ n49917;
  assign n49933 = n49932 ^ n49909;
  assign n49934 = n49913 & ~n49933;
  assign n49935 = n49934 ^ n49912;
  assign n49936 = n49935 ^ n49904;
  assign n49937 = n49908 & ~n49936;
  assign n49938 = n49937 ^ n49907;
  assign n49939 = n49938 ^ n49899;
  assign n49940 = ~n49903 & n49939;
  assign n49941 = n49940 ^ n49902;
  assign n49942 = n49941 ^ n49897;
  assign n49943 = n49898 & ~n49942;
  assign n49944 = n49943 ^ n49896;
  assign n49945 = n49944 ^ n49889;
  assign n49946 = n49893 & ~n49945;
  assign n49947 = n49946 ^ n49892;
  assign n49948 = n49947 ^ n49884;
  assign n49949 = ~n49888 & n49948;
  assign n49950 = n49949 ^ n49887;
  assign n49951 = n49950 ^ n49879;
  assign n49952 = ~n49883 & n49951;
  assign n49953 = n49952 ^ n49882;
  assign n49954 = n49953 ^ n49874;
  assign n49955 = ~n49878 & n49954;
  assign n49956 = n49955 ^ n49877;
  assign n49957 = n49956 ^ n49871;
  assign n49958 = n49873 & ~n49957;
  assign n49959 = n49958 ^ n49872;
  assign n49960 = n49959 ^ n49864;
  assign n49961 = ~n49868 & n49960;
  assign n49962 = n49961 ^ n49867;
  assign n49963 = n49962 ^ n49859;
  assign n49964 = ~n49863 & n49963;
  assign n49965 = n49964 ^ n49862;
  assign n49981 = n49980 ^ n49965;
  assign n49668 = n47719 ^ n40245;
  assign n49669 = n49668 ^ n44260;
  assign n49670 = n49669 ^ n38725;
  assign n49982 = n49981 ^ n49670;
  assign n51795 = n49982 ^ n49367;
  assign n50405 = n48448 ^ n40995;
  assign n50406 = n50405 ^ n45061;
  assign n50407 = n50406 ^ n39138;
  assign n50380 = n49941 ^ n49898;
  assign n50378 = n49346 ^ n48686;
  assign n50025 = n49314 ^ n49166;
  assign n50379 = n50378 ^ n50025;
  assign n50381 = n50380 ^ n50379;
  assign n50366 = n49938 ^ n49903;
  assign n50351 = n49065 ^ n48613;
  assign n50352 = n50351 ^ n49973;
  assign n50350 = n49935 ^ n49908;
  assign n50353 = n50352 ^ n50350;
  assign n50337 = n49823 ^ n48938;
  assign n50338 = n50337 ^ n48566;
  assign n50335 = n49932 ^ n49912;
  assign n50336 = n50335 ^ n49909;
  assign n50339 = n50338 ^ n50336;
  assign n50323 = n49929 ^ n49918;
  assign n50267 = n48778 ^ n48298;
  assign n50268 = n50267 ^ n49674;
  assign n50266 = n49926 ^ n49923;
  assign n50269 = n50268 ^ n50266;
  assign n49631 = n49630 ^ n48780;
  assign n49632 = n49631 ^ n48187;
  assign n49629 = n49628 ^ n49609;
  assign n50262 = n49632 ^ n49629;
  assign n50159 = n49606 ^ n2066;
  assign n50160 = n50159 ^ n49513;
  assign n49638 = n49637 ^ n48799;
  assign n49639 = n49638 ^ n48203;
  assign n49635 = n49592 ^ n49524;
  assign n49640 = n49639 ^ n49635;
  assign n49643 = n48808 ^ n48268;
  assign n49646 = n49645 ^ n49643;
  assign n49642 = n49586 ^ n49534;
  assign n49647 = n49646 ^ n49642;
  assign n50128 = n49583 ^ n49539;
  assign n49650 = n49649 ^ n48181;
  assign n49651 = n49650 ^ n48893;
  assign n49648 = n49580 ^ n49577;
  assign n49652 = n49651 ^ n49648;
  assign n50118 = n49572 ^ n49544;
  assign n49654 = n48221 ^ n48180;
  assign n49655 = n49654 ^ n49619;
  assign n49653 = n49569 ^ n49566;
  assign n49656 = n49655 ^ n49653;
  assign n50108 = n49561 ^ n49558;
  assign n49659 = n49552 ^ n49496;
  assign n49660 = n49659 ^ n49549;
  assign n49657 = n48823 ^ n48228;
  assign n49658 = n49657 ^ n49419;
  assign n49661 = n49660 ^ n49658;
  assign n49664 = n49548 ^ n49547;
  assign n49662 = n48757 ^ n48234;
  assign n49663 = n49662 ^ n48766;
  assign n49665 = n49664 ^ n49663;
  assign n50029 = n48623 ^ n47352;
  assign n50030 = n50029 ^ n47960;
  assign n50060 = n50030 ^ n50025;
  assign n50003 = n49311 ^ n49171;
  assign n50000 = n49973 ^ n49972;
  assign n50001 = ~n49976 & n50000;
  assign n50002 = n50001 ^ n49975;
  assign n50004 = n50003 ^ n50002;
  assign n49998 = n47964 ^ n47358;
  assign n49999 = n49998 ^ n48580;
  assign n50026 = n50003 ^ n49999;
  assign n50027 = n50004 & ~n50026;
  assign n50028 = n50027 ^ n49999;
  assign n50061 = n50028 ^ n50025;
  assign n50062 = n50060 & ~n50061;
  assign n50063 = n50062 ^ n50030;
  assign n50057 = n47993 ^ n47283;
  assign n50058 = n50057 ^ n48659;
  assign n50056 = n49317 ^ n49161;
  assign n50059 = n50058 ^ n50056;
  assign n50064 = n50063 ^ n50059;
  assign n50065 = n50064 ^ n46647;
  assign n50031 = n50030 ^ n50028;
  assign n50032 = n50031 ^ n50025;
  assign n50033 = n50032 ^ n46617;
  assign n50005 = n50004 ^ n49999;
  assign n50006 = n50005 ^ n46619;
  assign n49994 = n49977 ^ n46634;
  assign n49995 = n49977 ^ n49968;
  assign n49996 = ~n49994 & ~n49995;
  assign n49997 = n49996 ^ n46634;
  assign n50022 = n50005 ^ n49997;
  assign n50023 = ~n50006 & n50022;
  assign n50024 = n50023 ^ n46619;
  assign n50053 = n50032 ^ n50024;
  assign n50054 = n50033 & ~n50053;
  assign n50055 = n50054 ^ n46617;
  assign n50066 = n50065 ^ n50055;
  assign n49993 = ~n49978 & ~n49979;
  assign n50007 = n50006 ^ n49997;
  assign n50021 = ~n49993 & ~n50007;
  assign n50034 = n50033 ^ n50024;
  assign n50067 = n50021 & n50034;
  assign n50091 = ~n50066 & ~n50067;
  assign n50086 = n47710 ^ n40231;
  assign n50087 = n50086 ^ n44484;
  assign n50088 = n50087 ^ n38477;
  assign n50084 = n49348 ^ n47208;
  assign n50083 = n49320 ^ n49156;
  assign n50085 = n50084 ^ n50083;
  assign n50089 = n50088 ^ n50085;
  assign n50080 = n50064 ^ n50055;
  assign n50081 = n50065 & n50080;
  assign n50082 = n50081 ^ n46647;
  assign n50090 = n50089 ^ n50082;
  assign n50092 = n50091 ^ n50090;
  assign n50093 = n50092 ^ n48694;
  assign n50077 = n50063 ^ n50056;
  assign n50078 = ~n50059 & ~n50077;
  assign n50079 = n50078 ^ n50058;
  assign n50094 = n50093 ^ n50079;
  assign n50068 = n50067 ^ n50066;
  assign n50050 = n47933 ^ n40235;
  assign n50051 = n50050 ^ n43760;
  assign n50052 = n50051 ^ n38716;
  assign n50069 = n50068 ^ n50052;
  assign n50035 = n50034 ^ n50021;
  assign n50017 = n47715 ^ n40241;
  assign n50018 = n50017 ^ n44251;
  assign n50019 = n50018 ^ n38815;
  assign n50046 = n50035 ^ n50019;
  assign n50008 = n50007 ^ n49993;
  assign n49990 = n49980 ^ n49670;
  assign n49991 = n49981 & ~n49990;
  assign n49992 = n49991 ^ n49670;
  assign n50009 = n50008 ^ n49992;
  assign n49987 = n47922 ^ n40282;
  assign n49988 = n49987 ^ n44255;
  assign n49989 = n49988 ^ n38721;
  assign n50014 = n50008 ^ n49989;
  assign n50015 = ~n50009 & n50014;
  assign n50016 = n50015 ^ n49989;
  assign n50047 = n50035 ^ n50016;
  assign n50048 = n50046 & ~n50047;
  assign n50049 = n50048 ^ n50019;
  assign n50074 = n50052 ^ n50049;
  assign n50075 = ~n50069 & ~n50074;
  assign n50076 = n50075 ^ n50068;
  assign n50095 = n50094 ^ n50076;
  assign n50043 = n49404 ^ n48829;
  assign n50044 = n50043 ^ n48170;
  assign n50020 = n50019 ^ n50016;
  assign n50036 = n50035 ^ n50020;
  assign n49983 = n48772 ^ n48004;
  assign n49984 = n49983 ^ n48835;
  assign n49985 = ~n49982 & n49984;
  assign n49666 = n48852 ^ n48771;
  assign n49667 = n49666 ^ n48014;
  assign n49986 = n49985 ^ n49667;
  assign n50010 = n50009 ^ n49989;
  assign n50011 = n50010 ^ n49667;
  assign n50012 = ~n49986 & n50011;
  assign n50013 = n50012 ^ n49985;
  assign n50037 = n50036 ^ n50013;
  assign n50038 = n48773 ^ n48765;
  assign n50039 = n50038 ^ n48061;
  assign n50040 = n50039 ^ n50036;
  assign n50041 = ~n50037 & ~n50040;
  assign n50042 = n50041 ^ n50039;
  assign n50045 = n50044 ^ n50042;
  assign n50070 = n50069 ^ n50049;
  assign n50071 = n50070 ^ n50042;
  assign n50072 = n50045 & ~n50071;
  assign n50073 = n50072 ^ n50044;
  assign n50096 = n50095 ^ n50073;
  assign n50097 = n48759 ^ n48240;
  assign n50098 = n50097 ^ n48828;
  assign n50099 = n50098 ^ n50095;
  assign n50100 = n50096 & n50099;
  assign n50101 = n50100 ^ n50098;
  assign n50102 = n50101 ^ n49664;
  assign n50103 = n49665 & ~n50102;
  assign n50104 = n50103 ^ n49663;
  assign n50105 = n50104 ^ n49660;
  assign n50106 = ~n49661 & ~n50105;
  assign n50107 = n50106 ^ n49658;
  assign n50109 = n50108 ^ n50107;
  assign n50110 = n49485 ^ n48226;
  assign n50111 = n50110 ^ n48760;
  assign n50112 = n50111 ^ n50108;
  assign n50113 = n50109 & ~n50112;
  assign n50114 = n50113 ^ n50111;
  assign n50115 = n50114 ^ n49653;
  assign n50116 = ~n49656 & ~n50115;
  assign n50117 = n50116 ^ n49655;
  assign n50119 = n50118 ^ n50117;
  assign n50120 = n49711 ^ n48217;
  assign n50121 = n50120 ^ n48816;
  assign n50122 = n50121 ^ n50118;
  assign n50123 = ~n50119 & ~n50122;
  assign n50124 = n50123 ^ n50121;
  assign n50125 = n50124 ^ n49648;
  assign n50126 = n49652 & ~n50125;
  assign n50127 = n50126 ^ n49651;
  assign n50129 = n50128 ^ n50127;
  assign n50130 = n48812 ^ n48210;
  assign n50131 = n50130 ^ n49704;
  assign n50132 = n50131 ^ n50128;
  assign n50133 = ~n50129 & ~n50132;
  assign n50134 = n50133 ^ n50131;
  assign n50135 = n50134 ^ n49642;
  assign n50136 = ~n49647 & ~n50135;
  assign n50137 = n50136 ^ n49646;
  assign n49641 = n49589 ^ n49529;
  assign n50138 = n50137 ^ n49641;
  assign n50139 = n48804 ^ n48207;
  assign n50140 = n50139 ^ n49699;
  assign n50141 = n50140 ^ n49641;
  assign n50142 = n50138 & n50141;
  assign n50143 = n50142 ^ n50140;
  assign n50144 = n50143 ^ n49635;
  assign n50145 = n49640 & ~n50144;
  assign n50146 = n50145 ^ n49639;
  assign n49634 = n49600 ^ n49599;
  assign n50147 = n50146 ^ n49634;
  assign n50148 = n49689 ^ n48199;
  assign n50149 = n50148 ^ n48794;
  assign n50150 = n50149 ^ n49634;
  assign n50151 = n50147 & ~n50150;
  assign n50152 = n50151 ^ n50149;
  assign n49633 = n49603 ^ n49519;
  assign n50153 = n50152 ^ n49633;
  assign n50154 = n48788 ^ n48197;
  assign n50155 = n50154 ^ n49685;
  assign n50156 = n50155 ^ n49633;
  assign n50157 = n50153 & n50156;
  assign n50158 = n50157 ^ n50155;
  assign n50161 = n50160 ^ n50158;
  assign n50162 = n48784 ^ n48193;
  assign n50163 = n50162 ^ n49683;
  assign n50164 = n50163 ^ n50160;
  assign n50165 = ~n50161 & n50164;
  assign n50166 = n50165 ^ n50163;
  assign n50263 = n50166 ^ n49629;
  assign n50264 = n50262 & n50263;
  assign n50265 = n50264 ^ n49632;
  assign n50320 = n50266 ^ n50265;
  assign n50321 = ~n50269 & n50320;
  assign n50322 = n50321 ^ n50268;
  assign n50324 = n50323 ^ n50322;
  assign n50318 = n49751 ^ n48776;
  assign n50319 = n50318 ^ n48392;
  assign n50332 = n50323 ^ n50319;
  assign n50333 = ~n50324 & n50332;
  assign n50334 = n50333 ^ n50319;
  assign n50347 = n50336 ^ n50334;
  assign n50348 = n50339 & ~n50347;
  assign n50349 = n50348 ^ n50338;
  assign n50363 = n50350 ^ n50349;
  assign n50364 = ~n50353 & ~n50363;
  assign n50365 = n50364 ^ n50352;
  assign n50367 = n50366 ^ n50365;
  assign n50361 = n50003 ^ n49127;
  assign n50362 = n50361 ^ n48647;
  assign n50375 = n50366 ^ n50362;
  assign n50376 = ~n50367 & n50375;
  assign n50377 = n50376 ^ n50362;
  assign n50382 = n50381 ^ n50377;
  assign n50383 = n50382 ^ n47953;
  assign n50368 = n50367 ^ n50362;
  assign n50369 = n50368 ^ n47632;
  assign n50354 = n50353 ^ n50349;
  assign n50355 = n50354 ^ n47622;
  assign n50340 = n50339 ^ n50334;
  assign n50341 = n50340 ^ n47476;
  assign n50325 = n50324 ^ n50319;
  assign n50326 = n50325 ^ n47469;
  assign n50270 = n50269 ^ n50265;
  assign n50271 = n50270 ^ n47461;
  assign n50167 = n50166 ^ n49632;
  assign n50168 = n50167 ^ n49629;
  assign n50169 = n50168 ^ n47216;
  assign n50170 = n50163 ^ n50161;
  assign n50171 = n50170 ^ n47451;
  assign n50172 = n50155 ^ n50153;
  assign n50173 = n50172 ^ n47223;
  assign n50174 = n50149 ^ n50147;
  assign n50175 = n50174 ^ n47227;
  assign n50244 = n50143 ^ n49639;
  assign n50245 = n50244 ^ n49635;
  assign n50239 = n50140 ^ n50138;
  assign n50176 = n50134 ^ n49646;
  assign n50177 = n50176 ^ n49642;
  assign n50178 = n50177 ^ n47237;
  assign n50179 = n50131 ^ n50129;
  assign n50180 = n50179 ^ n47241;
  assign n50181 = n50124 ^ n49652;
  assign n50182 = n50181 ^ n47246;
  assign n50183 = n50121 ^ n50119;
  assign n50184 = n50183 ^ n47249;
  assign n50185 = n50114 ^ n49656;
  assign n50186 = n50185 ^ n47251;
  assign n50187 = n50111 ^ n50109;
  assign n50188 = n50187 ^ n47252;
  assign n50189 = n50104 ^ n49661;
  assign n50190 = n50189 ^ n47256;
  assign n50191 = n50101 ^ n49665;
  assign n50192 = n50191 ^ n47263;
  assign n50205 = n50070 ^ n50045;
  assign n50193 = n50039 ^ n50037;
  assign n50194 = n50193 ^ n47265;
  assign n50195 = n49984 ^ n49982;
  assign n50196 = n47276 & ~n50195;
  assign n50197 = n50196 ^ n47270;
  assign n50198 = n50010 ^ n49986;
  assign n50199 = n50198 ^ n50196;
  assign n50200 = n50197 & n50199;
  assign n50201 = n50200 ^ n47270;
  assign n50202 = n50201 ^ n50193;
  assign n50203 = n50194 & n50202;
  assign n50204 = n50203 ^ n47265;
  assign n50206 = n50205 ^ n50204;
  assign n50207 = n50205 ^ n47392;
  assign n50208 = ~n50206 & n50207;
  assign n50209 = n50208 ^ n47392;
  assign n50210 = n50209 ^ n47210;
  assign n50211 = n50098 ^ n50096;
  assign n50212 = n50211 ^ n50209;
  assign n50213 = n50210 & ~n50212;
  assign n50214 = n50213 ^ n47210;
  assign n50215 = n50214 ^ n50191;
  assign n50216 = ~n50192 & n50215;
  assign n50217 = n50216 ^ n47263;
  assign n50218 = n50217 ^ n50189;
  assign n50219 = ~n50190 & ~n50218;
  assign n50220 = n50219 ^ n47256;
  assign n50221 = n50220 ^ n50187;
  assign n50222 = n50188 & ~n50221;
  assign n50223 = n50222 ^ n47252;
  assign n50224 = n50223 ^ n50185;
  assign n50225 = n50186 & ~n50224;
  assign n50226 = n50225 ^ n47251;
  assign n50227 = n50226 ^ n50183;
  assign n50228 = n50184 & n50227;
  assign n50229 = n50228 ^ n47249;
  assign n50230 = n50229 ^ n50181;
  assign n50231 = ~n50182 & ~n50230;
  assign n50232 = n50231 ^ n47246;
  assign n50233 = n50232 ^ n50179;
  assign n50234 = ~n50180 & ~n50233;
  assign n50235 = n50234 ^ n47241;
  assign n50236 = n50235 ^ n50177;
  assign n50237 = n50178 & ~n50236;
  assign n50238 = n50237 ^ n47237;
  assign n50240 = n50239 ^ n50238;
  assign n50241 = n50239 ^ n47233;
  assign n50242 = ~n50240 & n50241;
  assign n50243 = n50242 ^ n47233;
  assign n50246 = n50245 ^ n50243;
  assign n50247 = n50245 ^ n47228;
  assign n50248 = n50246 & n50247;
  assign n50249 = n50248 ^ n47228;
  assign n50250 = n50249 ^ n50174;
  assign n50251 = n50175 & n50250;
  assign n50252 = n50251 ^ n47227;
  assign n50253 = n50252 ^ n50172;
  assign n50254 = ~n50173 & n50253;
  assign n50255 = n50254 ^ n47223;
  assign n50256 = n50255 ^ n50170;
  assign n50257 = n50171 & ~n50256;
  assign n50258 = n50257 ^ n47451;
  assign n50259 = n50258 ^ n50168;
  assign n50260 = n50169 & ~n50259;
  assign n50261 = n50260 ^ n47216;
  assign n50315 = n50270 ^ n50261;
  assign n50316 = ~n50271 & ~n50315;
  assign n50317 = n50316 ^ n47461;
  assign n50329 = n50325 ^ n50317;
  assign n50330 = ~n50326 & ~n50329;
  assign n50331 = n50330 ^ n47469;
  assign n50344 = n50340 ^ n50331;
  assign n50345 = n50341 & n50344;
  assign n50346 = n50345 ^ n47476;
  assign n50358 = n50354 ^ n50346;
  assign n50359 = n50355 & n50358;
  assign n50360 = n50359 ^ n47622;
  assign n50372 = n50368 ^ n50360;
  assign n50373 = n50369 & ~n50372;
  assign n50374 = n50373 ^ n47632;
  assign n50384 = n50383 ^ n50374;
  assign n50272 = n50271 ^ n50261;
  assign n50273 = n50235 ^ n50178;
  assign n50274 = n50232 ^ n47241;
  assign n50275 = n50274 ^ n50179;
  assign n50276 = n50229 ^ n50182;
  assign n50277 = n50220 ^ n47252;
  assign n50278 = n50277 ^ n50187;
  assign n50279 = n50198 ^ n50197;
  assign n50280 = n50201 ^ n50194;
  assign n50281 = n50279 & ~n50280;
  assign n50282 = n50206 ^ n47392;
  assign n50283 = ~n50281 & ~n50282;
  assign n50284 = n50211 ^ n47210;
  assign n50285 = n50284 ^ n50209;
  assign n50286 = ~n50283 & n50285;
  assign n50287 = n50214 ^ n50192;
  assign n50288 = ~n50286 & n50287;
  assign n50289 = n50217 ^ n50190;
  assign n50290 = ~n50288 & ~n50289;
  assign n50291 = ~n50278 & n50290;
  assign n50292 = n50223 ^ n50186;
  assign n50293 = n50291 & ~n50292;
  assign n50294 = n50226 ^ n47249;
  assign n50295 = n50294 ^ n50183;
  assign n50296 = ~n50293 & n50295;
  assign n50297 = n50276 & n50296;
  assign n50298 = ~n50275 & n50297;
  assign n50299 = ~n50273 & n50298;
  assign n50300 = n50240 ^ n47233;
  assign n50301 = n50299 & ~n50300;
  assign n50302 = n50246 ^ n47228;
  assign n50303 = ~n50301 & n50302;
  assign n50304 = n50249 ^ n47227;
  assign n50305 = n50304 ^ n50174;
  assign n50306 = n50303 & ~n50305;
  assign n50307 = n50252 ^ n50173;
  assign n50308 = ~n50306 & n50307;
  assign n50309 = n50255 ^ n47451;
  assign n50310 = n50309 ^ n50170;
  assign n50311 = ~n50308 & n50310;
  assign n50312 = n50258 ^ n50169;
  assign n50313 = ~n50311 & ~n50312;
  assign n50314 = n50272 & n50313;
  assign n50327 = n50326 ^ n50317;
  assign n50328 = n50314 & ~n50327;
  assign n50342 = n50341 ^ n50331;
  assign n50343 = ~n50328 & n50342;
  assign n50356 = n50355 ^ n50346;
  assign n50357 = n50343 & ~n50356;
  assign n50370 = n50369 ^ n50360;
  assign n50371 = ~n50357 & ~n50370;
  assign n50404 = n50384 ^ n50371;
  assign n50408 = n50407 ^ n50404;
  assign n50410 = n48452 ^ n41000;
  assign n50411 = n50410 ^ n45150;
  assign n50412 = n50411 ^ n39142;
  assign n50409 = n50370 ^ n50357;
  assign n50413 = n50412 ^ n50409;
  assign n50586 = n50356 ^ n50343;
  assign n50415 = n48462 ^ n41030;
  assign n50416 = n50415 ^ n45071;
  assign n50417 = n50416 ^ n39307;
  assign n50414 = n50342 ^ n50328;
  assign n50418 = n50417 ^ n50414;
  assign n50420 = n48468 ^ n41009;
  assign n50421 = n50420 ^ n45136;
  assign n50422 = n50421 ^ n39153;
  assign n50419 = n50327 ^ n50314;
  assign n50423 = n50422 ^ n50419;
  assign n50572 = n50313 ^ n50272;
  assign n50425 = n48473 ^ n40654;
  assign n50426 = n50425 ^ n45120;
  assign n50427 = n50426 ^ n39157;
  assign n50424 = n50312 ^ n50311;
  assign n50428 = n50427 ^ n50424;
  assign n50561 = n50310 ^ n50308;
  assign n50430 = n48483 ^ n40517;
  assign n50431 = n50430 ^ n45081;
  assign n50432 = n50431 ^ n39168;
  assign n50429 = n50307 ^ n50306;
  assign n50433 = n50432 ^ n50429;
  assign n50435 = n48488 ^ n40625;
  assign n50436 = n50435 ^ n45086;
  assign n50437 = n50436 ^ n39279;
  assign n50434 = n50305 ^ n50303;
  assign n50438 = n50437 ^ n50434;
  assign n50440 = n40522 ^ n2253;
  assign n50441 = n50440 ^ n45091;
  assign n50442 = n50441 ^ n39173;
  assign n50439 = n50302 ^ n50301;
  assign n50443 = n50442 ^ n50439;
  assign n50445 = n48495 ^ n2158;
  assign n50446 = n50445 ^ n45096;
  assign n50447 = n50446 ^ n39178;
  assign n50444 = n50300 ^ n50299;
  assign n50448 = n50447 ^ n50444;
  assign n50450 = n48500 ^ n2140;
  assign n50451 = n50450 ^ n44743;
  assign n50452 = n50451 ^ n39183;
  assign n50449 = n50298 ^ n50273;
  assign n50453 = n50452 ^ n50449;
  assign n50538 = n50297 ^ n50275;
  assign n50455 = n48087 ^ n40534;
  assign n50456 = n50455 ^ n44719;
  assign n50457 = n50456 ^ n39193;
  assign n50454 = n50296 ^ n50276;
  assign n50458 = n50457 ^ n50454;
  assign n50527 = n50295 ^ n50293;
  assign n50460 = n48097 ^ n40538;
  assign n50461 = n50460 ^ n44708;
  assign n50462 = n50461 ^ n1685;
  assign n50459 = n50292 ^ n50291;
  assign n50463 = n50462 ^ n50459;
  assign n50516 = n48102 ^ n40544;
  assign n50517 = n50516 ^ n44654;
  assign n50518 = n50517 ^ n39199;
  assign n50465 = n48107 ^ n40548;
  assign n50466 = n50465 ^ n44697;
  assign n50467 = n50466 ^ n39204;
  assign n50464 = n50289 ^ n50288;
  assign n50468 = n50467 ^ n50464;
  assign n50505 = n48112 ^ n40553;
  assign n50506 = n50505 ^ n44660;
  assign n50507 = n50506 ^ n39210;
  assign n50497 = n48117 ^ n40580;
  assign n50498 = n50497 ^ n44665;
  assign n50499 = n50498 ^ n39236;
  assign n50470 = n48133 ^ n40558;
  assign n50471 = n50470 ^ n44669;
  assign n50472 = n50471 ^ n39214;
  assign n50469 = n50282 ^ n50281;
  assign n50473 = n50472 ^ n50469;
  assign n50475 = n48121 ^ n40562;
  assign n50476 = n50475 ^ n44679;
  assign n50477 = n50476 ^ n39218;
  assign n50474 = n50280 ^ n50279;
  assign n50478 = n50477 ^ n50474;
  assign n50482 = n48675 ^ n40771;
  assign n50483 = n50482 ^ n45247;
  assign n50484 = n50483 ^ n39440;
  assign n50485 = n50195 ^ n47276;
  assign n50486 = n50484 & ~n50485;
  assign n50479 = n48124 ^ n40565;
  assign n50480 = n50479 ^ n44674;
  assign n50481 = n50480 ^ n39221;
  assign n50487 = n50486 ^ n50481;
  assign n50488 = n50486 ^ n50279;
  assign n50489 = n50487 & ~n50488;
  assign n50490 = n50489 ^ n50481;
  assign n50491 = n50490 ^ n50474;
  assign n50492 = n50478 & ~n50491;
  assign n50493 = n50492 ^ n50477;
  assign n50494 = n50493 ^ n50469;
  assign n50495 = n50473 & ~n50494;
  assign n50496 = n50495 ^ n50472;
  assign n50500 = n50499 ^ n50496;
  assign n50501 = n50285 ^ n50283;
  assign n50502 = n50501 ^ n50496;
  assign n50503 = n50500 & ~n50502;
  assign n50504 = n50503 ^ n50499;
  assign n50508 = n50507 ^ n50504;
  assign n50509 = n50287 ^ n50286;
  assign n50510 = n50509 ^ n50504;
  assign n50511 = n50508 & n50510;
  assign n50512 = n50511 ^ n50507;
  assign n50513 = n50512 ^ n50464;
  assign n50514 = ~n50468 & n50513;
  assign n50515 = n50514 ^ n50467;
  assign n50519 = n50518 ^ n50515;
  assign n50520 = n50290 ^ n50278;
  assign n50521 = n50520 ^ n50515;
  assign n50522 = n50519 & ~n50521;
  assign n50523 = n50522 ^ n50518;
  assign n50524 = n50523 ^ n50459;
  assign n50525 = n50463 & ~n50524;
  assign n50526 = n50525 ^ n50462;
  assign n50528 = n50527 ^ n50526;
  assign n50529 = n48092 ^ n40600;
  assign n50530 = n50529 ^ n44650;
  assign n50531 = n50530 ^ n39256;
  assign n50532 = n50531 ^ n50527;
  assign n50533 = n50528 & ~n50532;
  assign n50534 = n50533 ^ n50531;
  assign n50535 = n50534 ^ n50454;
  assign n50536 = n50458 & ~n50535;
  assign n50537 = n50536 ^ n50457;
  assign n50539 = n50538 ^ n50537;
  assign n50540 = n48178 ^ n40529;
  assign n50541 = n50540 ^ n44645;
  assign n50542 = n50541 ^ n39188;
  assign n50543 = n50542 ^ n50538;
  assign n50544 = n50539 & ~n50543;
  assign n50545 = n50544 ^ n50542;
  assign n50546 = n50545 ^ n50449;
  assign n50547 = ~n50453 & n50546;
  assign n50548 = n50547 ^ n50452;
  assign n50549 = n50548 ^ n50444;
  assign n50550 = ~n50448 & n50549;
  assign n50551 = n50550 ^ n50447;
  assign n50552 = n50551 ^ n50439;
  assign n50553 = n50443 & ~n50552;
  assign n50554 = n50553 ^ n50442;
  assign n50555 = n50554 ^ n50434;
  assign n50556 = n50438 & ~n50555;
  assign n50557 = n50556 ^ n50437;
  assign n50558 = n50557 ^ n50429;
  assign n50559 = ~n50433 & n50558;
  assign n50560 = n50559 ^ n50432;
  assign n50562 = n50561 ^ n50560;
  assign n50566 = n50565 ^ n50561;
  assign n50567 = ~n50562 & n50566;
  assign n50568 = n50567 ^ n50565;
  assign n50569 = n50568 ^ n50424;
  assign n50570 = n50428 & ~n50569;
  assign n50571 = n50570 ^ n50427;
  assign n50573 = n50572 ^ n50571;
  assign n50574 = n48530 ^ n41015;
  assign n50575 = n50574 ^ n45128;
  assign n50576 = n50575 ^ n39296;
  assign n50577 = n50576 ^ n50572;
  assign n50578 = ~n50573 & n50577;
  assign n50579 = n50578 ^ n50576;
  assign n50580 = n50579 ^ n50419;
  assign n50581 = ~n50423 & n50580;
  assign n50582 = n50581 ^ n50422;
  assign n50583 = n50582 ^ n50414;
  assign n50584 = n50418 & ~n50583;
  assign n50585 = n50584 ^ n50417;
  assign n50587 = n50586 ^ n50585;
  assign n50588 = n48457 ^ n41005;
  assign n50589 = n50588 ^ n45066;
  assign n50590 = n50589 ^ n39148;
  assign n50591 = n50590 ^ n50586;
  assign n50592 = ~n50587 & n50591;
  assign n50593 = n50592 ^ n50590;
  assign n50594 = n50593 ^ n50409;
  assign n50595 = n50413 & ~n50594;
  assign n50596 = n50595 ^ n50412;
  assign n50597 = n50596 ^ n50404;
  assign n50598 = ~n50408 & n50597;
  assign n50599 = n50598 ^ n50407;
  assign n50400 = n48443 ^ n1011;
  assign n50401 = n50400 ^ n45161;
  assign n50402 = n50401 ^ n39339;
  assign n50394 = n49944 ^ n49893;
  assign n50392 = n50056 ^ n48583;
  assign n50393 = n50392 ^ n47974;
  assign n50395 = n50394 ^ n50393;
  assign n50389 = n50380 ^ n50377;
  assign n50390 = ~n50381 & n50389;
  assign n50391 = n50390 ^ n50379;
  assign n50396 = n50395 ^ n50391;
  assign n50397 = n50396 ^ n47192;
  assign n50386 = n50382 ^ n50374;
  assign n50387 = n50383 & n50386;
  assign n50388 = n50387 ^ n47953;
  assign n50398 = n50397 ^ n50388;
  assign n50385 = n50371 & ~n50384;
  assign n50399 = n50398 ^ n50385;
  assign n50403 = n50402 ^ n50399;
  assign n51401 = n50599 ^ n50403;
  assign n51796 = n51795 ^ n51401;
  assign n50825 = n50336 ^ n49630;
  assign n50826 = n50825 ^ n48788;
  assign n50824 = n50542 ^ n50539;
  assign n50827 = n50826 ^ n50824;
  assign n50929 = n50534 ^ n50458;
  assign n50829 = n50266 ^ n48799;
  assign n50830 = n50829 ^ n49685;
  assign n50828 = n50531 ^ n50528;
  assign n50831 = n50830 ^ n50828;
  assign n50913 = n50520 ^ n50519;
  assign n50894 = n50501 ^ n50500;
  assign n50886 = n50493 ^ n50472;
  assign n50887 = n50886 ^ n50469;
  assign n50879 = n50490 ^ n50478;
  assign n50834 = n50128 ^ n49619;
  assign n50835 = n50834 ^ n48823;
  assign n50832 = n50481 ^ n50279;
  assign n50833 = n50832 ^ n50486;
  assign n50836 = n50835 ^ n50833;
  assign n50838 = n49648 ^ n48766;
  assign n50839 = n50838 ^ n49485;
  assign n50837 = n50485 ^ n50484;
  assign n50840 = n50839 ^ n50837;
  assign n50862 = n48642 ^ n44797;
  assign n50863 = n50862 ^ n40976;
  assign n50864 = n50863 ^ n39542;
  assign n50755 = n48750 ^ n47993;
  assign n50756 = n50755 ^ n49362;
  assign n50713 = n49956 ^ n49873;
  assign n50671 = n49953 ^ n49878;
  assign n50633 = n49950 ^ n49882;
  assign n50634 = n50633 ^ n49879;
  assign n50612 = n49947 ^ n49888;
  assign n50609 = n50394 ^ n50391;
  assign n50610 = ~n50395 & n50609;
  assign n50611 = n50610 ^ n50393;
  assign n50613 = n50612 ^ n50611;
  assign n50607 = n48580 ^ n47980;
  assign n50608 = n50607 ^ n50083;
  assign n50630 = n50612 ^ n50608;
  assign n50631 = ~n50613 & n50630;
  assign n50632 = n50631 ^ n50608;
  assign n50635 = n50634 ^ n50632;
  assign n50628 = n48623 ^ n47970;
  assign n50629 = n50628 ^ n49367;
  assign n50668 = n50634 ^ n50629;
  assign n50669 = ~n50635 & ~n50668;
  assign n50670 = n50669 ^ n50629;
  assign n50672 = n50671 ^ n50670;
  assign n50666 = n48659 ^ n47964;
  assign n50667 = n50666 ^ n49372;
  assign n50710 = n50671 ^ n50667;
  assign n50711 = n50672 & ~n50710;
  assign n50712 = n50711 ^ n50667;
  assign n50714 = n50713 ^ n50712;
  assign n50708 = n48694 ^ n47960;
  assign n50709 = n50708 ^ n49379;
  assign n50751 = n50713 ^ n50709;
  assign n50752 = ~n50714 & ~n50751;
  assign n50753 = n50752 ^ n50709;
  assign n50750 = n49959 ^ n49868;
  assign n50754 = n50753 ^ n50750;
  assign n50757 = n50756 ^ n50754;
  assign n50758 = n50757 ^ n47283;
  assign n50715 = n50714 ^ n50709;
  assign n50716 = n50715 ^ n47352;
  assign n50673 = n50672 ^ n50667;
  assign n50674 = n50673 ^ n47358;
  assign n50636 = n50635 ^ n50629;
  assign n50637 = n50636 ^ n47361;
  assign n50614 = n50613 ^ n50608;
  assign n50615 = n50614 ^ n47188;
  assign n50604 = n50396 ^ n50388;
  assign n50605 = ~n50397 & ~n50604;
  assign n50606 = n50605 ^ n47192;
  assign n50625 = n50614 ^ n50606;
  assign n50626 = n50615 & ~n50625;
  assign n50627 = n50626 ^ n47188;
  assign n50663 = n50636 ^ n50627;
  assign n50664 = ~n50637 & n50663;
  assign n50665 = n50664 ^ n47361;
  assign n50705 = n50673 ^ n50665;
  assign n50706 = ~n50674 & ~n50705;
  assign n50707 = n50706 ^ n47358;
  assign n50747 = n50715 ^ n50707;
  assign n50748 = ~n50716 & n50747;
  assign n50749 = n50748 ^ n47352;
  assign n50759 = n50758 ^ n50749;
  assign n50717 = n50716 ^ n50707;
  assign n50638 = n50637 ^ n50627;
  assign n50603 = ~n50385 & n50398;
  assign n50616 = n50615 ^ n50606;
  assign n50639 = ~n50603 & ~n50616;
  assign n50662 = ~n50638 & ~n50639;
  assign n50675 = n50674 ^ n50665;
  assign n50718 = ~n50662 & n50675;
  assign n50760 = ~n50717 & n50718;
  assign n50860 = n50759 & ~n50760;
  assign n50857 = n49962 ^ n49863;
  assign n50854 = n48840 ^ n47208;
  assign n50855 = n50854 ^ n49358;
  assign n50851 = n50756 ^ n50750;
  assign n50852 = ~n50754 & ~n50851;
  assign n50853 = n50852 ^ n50756;
  assign n50856 = n50855 ^ n50853;
  assign n50858 = n50857 ^ n50856;
  assign n50847 = n50757 ^ n50749;
  assign n50848 = ~n50758 & ~n50847;
  assign n50849 = n50848 ^ n47283;
  assign n50850 = n50849 ^ n47279;
  assign n50859 = n50858 ^ n50850;
  assign n50861 = n50860 ^ n50859;
  assign n50865 = n50864 ^ n50861;
  assign n50761 = n50760 ^ n50759;
  assign n50720 = n48578 ^ n41064;
  assign n50721 = n50720 ^ n1361;
  assign n50722 = n50721 ^ n39549;
  assign n50719 = n50718 ^ n50717;
  assign n50723 = n50722 ^ n50719;
  assign n50677 = n48186 ^ n40985;
  assign n50678 = n50677 ^ n45175;
  assign n50679 = n50678 ^ n1353;
  assign n50676 = n50675 ^ n50662;
  assign n50680 = n50679 ^ n50676;
  assign n50640 = n50639 ^ n50638;
  assign n1155 = n1154 ^ n1109;
  assign n1189 = n1188 ^ n1155;
  assign n1199 = n1198 ^ n1189;
  assign n50641 = n50640 ^ n1199;
  assign n50617 = n50616 ^ n50603;
  assign n50600 = n50599 ^ n50399;
  assign n50601 = n50403 & ~n50600;
  assign n50602 = n50601 ^ n50402;
  assign n50618 = n50617 ^ n50602;
  assign n50619 = n48438 ^ n41050;
  assign n50620 = n50619 ^ n45056;
  assign n50621 = n50620 ^ n1180;
  assign n50622 = n50621 ^ n50617;
  assign n50623 = ~n50618 & n50622;
  assign n50624 = n50623 ^ n50621;
  assign n50659 = n50640 ^ n50624;
  assign n50660 = ~n50641 & n50659;
  assign n50661 = n50660 ^ n1199;
  assign n50702 = n50676 ^ n50661;
  assign n50703 = ~n50680 & n50702;
  assign n50704 = n50703 ^ n50679;
  assign n50744 = n50719 ^ n50704;
  assign n50745 = ~n50723 & n50744;
  assign n50746 = n50745 ^ n50722;
  assign n50762 = n50761 ^ n50746;
  assign n50741 = n48603 ^ n40981;
  assign n50742 = n50741 ^ n44800;
  assign n50743 = n50742 ^ n2345;
  assign n50844 = n50761 ^ n50743;
  assign n50845 = ~n50762 & n50844;
  assign n50846 = n50845 ^ n50743;
  assign n50866 = n50865 ^ n50846;
  assign n50763 = n50762 ^ n50743;
  assign n50739 = n49653 ^ n48757;
  assign n50740 = n50739 ^ n48829;
  assign n50764 = n50763 ^ n50740;
  assign n50724 = n50723 ^ n50704;
  assign n50681 = n50680 ^ n50661;
  assign n50656 = n49660 ^ n49404;
  assign n50657 = n50656 ^ n48852;
  assign n50698 = n50681 ^ n50657;
  assign n50642 = n50641 ^ n50624;
  assign n50643 = n49664 ^ n48835;
  assign n50644 = n50643 ^ n48765;
  assign n50655 = ~n50642 & ~n50644;
  assign n50699 = n50681 ^ n50655;
  assign n50700 = ~n50698 & ~n50699;
  assign n50701 = n50700 ^ n50655;
  assign n50725 = n50724 ^ n50701;
  assign n50696 = n50108 ^ n48759;
  assign n50697 = n50696 ^ n48773;
  assign n50736 = n50724 ^ n50697;
  assign n50737 = n50725 & ~n50736;
  assign n50738 = n50737 ^ n50697;
  assign n50841 = n50763 ^ n50738;
  assign n50842 = ~n50764 & ~n50841;
  assign n50843 = n50842 ^ n50740;
  assign n50867 = n50866 ^ n50843;
  assign n50868 = n50118 ^ n49419;
  assign n50869 = n50868 ^ n48828;
  assign n50870 = n50869 ^ n50866;
  assign n50871 = n50867 & n50870;
  assign n50872 = n50871 ^ n50869;
  assign n50873 = n50872 ^ n50837;
  assign n50874 = ~n50840 & n50873;
  assign n50875 = n50874 ^ n50839;
  assign n50876 = n50875 ^ n50833;
  assign n50877 = ~n50836 & ~n50876;
  assign n50878 = n50877 ^ n50835;
  assign n50880 = n50879 ^ n50878;
  assign n50881 = n49711 ^ n48760;
  assign n50882 = n50881 ^ n49642;
  assign n50883 = n50882 ^ n50879;
  assign n50884 = n50880 & ~n50883;
  assign n50885 = n50884 ^ n50882;
  assign n50888 = n50887 ^ n50885;
  assign n50889 = n49649 ^ n48180;
  assign n50890 = n50889 ^ n49641;
  assign n50891 = n50890 ^ n50887;
  assign n50892 = n50888 & n50891;
  assign n50893 = n50892 ^ n50890;
  assign n50895 = n50894 ^ n50893;
  assign n50896 = n49704 ^ n48816;
  assign n50897 = n50896 ^ n49635;
  assign n50898 = n50897 ^ n50894;
  assign n50899 = ~n50895 & ~n50898;
  assign n50900 = n50899 ^ n50897;
  assign n50787 = n50509 ^ n50507;
  assign n50788 = n50787 ^ n50504;
  assign n50901 = n50900 ^ n50788;
  assign n50902 = n49634 ^ n48893;
  assign n50903 = n50902 ^ n49645;
  assign n50904 = n50903 ^ n50788;
  assign n50905 = ~n50901 & n50904;
  assign n50906 = n50905 ^ n50903;
  assign n50780 = n50512 ^ n50467;
  assign n50781 = n50780 ^ n50464;
  assign n50907 = n50906 ^ n50781;
  assign n50908 = n49633 ^ n48812;
  assign n50909 = n50908 ^ n49699;
  assign n50910 = n50909 ^ n50781;
  assign n50911 = ~n50907 & ~n50910;
  assign n50912 = n50911 ^ n50909;
  assign n50914 = n50913 ^ n50912;
  assign n50915 = n49637 ^ n48808;
  assign n50916 = n50915 ^ n50160;
  assign n50917 = n50916 ^ n50913;
  assign n50918 = ~n50914 & n50917;
  assign n50919 = n50918 ^ n50916;
  assign n50776 = n50523 ^ n50462;
  assign n50777 = n50776 ^ n50459;
  assign n50920 = n50919 ^ n50777;
  assign n50921 = n49689 ^ n48804;
  assign n50922 = n50921 ^ n49629;
  assign n50923 = n50922 ^ n50777;
  assign n50924 = ~n50920 & n50923;
  assign n50925 = n50924 ^ n50922;
  assign n50926 = n50925 ^ n50828;
  assign n50927 = n50831 & n50926;
  assign n50928 = n50927 ^ n50830;
  assign n50930 = n50929 ^ n50928;
  assign n50931 = n50323 ^ n49683;
  assign n50932 = n50931 ^ n48794;
  assign n50933 = n50932 ^ n50929;
  assign n50934 = n50930 & ~n50933;
  assign n50935 = n50934 ^ n50932;
  assign n50936 = n50935 ^ n50824;
  assign n50937 = n50827 & ~n50936;
  assign n50938 = n50937 ^ n50826;
  assign n50822 = n50545 ^ n50453;
  assign n50820 = n50350 ^ n49674;
  assign n50821 = n50820 ^ n48784;
  assign n50823 = n50822 ^ n50821;
  assign n51017 = n50938 ^ n50823;
  assign n51018 = n51017 ^ n48193;
  assign n51019 = n50935 ^ n50827;
  assign n51020 = n51019 ^ n48197;
  assign n51021 = n50932 ^ n50930;
  assign n51022 = n51021 ^ n48199;
  assign n51023 = n50925 ^ n50831;
  assign n51024 = n51023 ^ n48203;
  assign n51025 = n50922 ^ n50920;
  assign n51026 = n51025 ^ n48207;
  assign n51027 = n50916 ^ n50914;
  assign n51028 = n51027 ^ n48268;
  assign n51029 = n50909 ^ n50907;
  assign n51030 = n51029 ^ n48210;
  assign n51031 = n50903 ^ n50901;
  assign n51032 = n51031 ^ n48181;
  assign n51033 = n50897 ^ n50895;
  assign n51034 = n51033 ^ n48217;
  assign n51035 = n50890 ^ n50888;
  assign n51036 = n51035 ^ n48221;
  assign n51037 = n50882 ^ n50880;
  assign n51038 = n51037 ^ n48226;
  assign n51039 = n50875 ^ n50836;
  assign n51040 = n51039 ^ n48228;
  assign n51041 = n50872 ^ n50840;
  assign n51042 = n51041 ^ n48234;
  assign n51043 = n50869 ^ n50867;
  assign n51044 = n51043 ^ n48240;
  assign n50765 = n50764 ^ n50738;
  assign n50766 = n50765 ^ n48170;
  assign n50726 = n50725 ^ n50697;
  assign n50645 = n50644 ^ n50642;
  assign n50683 = n48004 & n50645;
  assign n50684 = n50683 ^ n48014;
  assign n50658 = n50657 ^ n50655;
  assign n50682 = n50681 ^ n50658;
  assign n50693 = n50683 ^ n50682;
  assign n50694 = ~n50684 & ~n50693;
  assign n50695 = n50694 ^ n48014;
  assign n50727 = n50726 ^ n50695;
  assign n50733 = n50726 ^ n48061;
  assign n50734 = ~n50727 & ~n50733;
  assign n50735 = n50734 ^ n48061;
  assign n51045 = n50765 ^ n50735;
  assign n51046 = n50766 & n51045;
  assign n51047 = n51046 ^ n48170;
  assign n51048 = n51047 ^ n51043;
  assign n51049 = n51044 & ~n51048;
  assign n51050 = n51049 ^ n48240;
  assign n51051 = n51050 ^ n51041;
  assign n51052 = ~n51042 & ~n51051;
  assign n51053 = n51052 ^ n48234;
  assign n51054 = n51053 ^ n51039;
  assign n51055 = n51040 & n51054;
  assign n51056 = n51055 ^ n48228;
  assign n51057 = n51056 ^ n51037;
  assign n51058 = n51038 & n51057;
  assign n51059 = n51058 ^ n48226;
  assign n51060 = n51059 ^ n51035;
  assign n51061 = ~n51036 & n51060;
  assign n51062 = n51061 ^ n48221;
  assign n51063 = n51062 ^ n51033;
  assign n51064 = ~n51034 & n51063;
  assign n51065 = n51064 ^ n48217;
  assign n51066 = n51065 ^ n51031;
  assign n51067 = ~n51032 & n51066;
  assign n51068 = n51067 ^ n48181;
  assign n51069 = n51068 ^ n51029;
  assign n51070 = n51030 & ~n51069;
  assign n51071 = n51070 ^ n48210;
  assign n51072 = n51071 ^ n51027;
  assign n51073 = n51028 & ~n51072;
  assign n51074 = n51073 ^ n48268;
  assign n51075 = n51074 ^ n51025;
  assign n51076 = ~n51026 & ~n51075;
  assign n51077 = n51076 ^ n48207;
  assign n51078 = n51077 ^ n51023;
  assign n51079 = n51024 & n51078;
  assign n51080 = n51079 ^ n48203;
  assign n51081 = n51080 ^ n51021;
  assign n51082 = n51022 & ~n51081;
  assign n51083 = n51082 ^ n48199;
  assign n51084 = n51083 ^ n51019;
  assign n51085 = n51020 & n51084;
  assign n51086 = n51085 ^ n48197;
  assign n51087 = n51086 ^ n51017;
  assign n51088 = n51018 & ~n51087;
  assign n51089 = n51088 ^ n48193;
  assign n50944 = n49751 ^ n48780;
  assign n50945 = n50944 ^ n50366;
  assign n50942 = n50548 ^ n50448;
  assign n50939 = n50938 ^ n50822;
  assign n50940 = n50823 & ~n50939;
  assign n50941 = n50940 ^ n50821;
  assign n50943 = n50942 ^ n50941;
  assign n51015 = n50945 ^ n50943;
  assign n51016 = n51015 ^ n48187;
  assign n51135 = n51089 ^ n51016;
  assign n51136 = n51086 ^ n51018;
  assign n51137 = n51080 ^ n51022;
  assign n51138 = n51077 ^ n51024;
  assign n51139 = n51074 ^ n51026;
  assign n51140 = n51068 ^ n51030;
  assign n51141 = n51065 ^ n51032;
  assign n51142 = n51056 ^ n51038;
  assign n50767 = n50766 ^ n50735;
  assign n50685 = n50684 ^ n50682;
  assign n50728 = n50727 ^ n48061;
  assign n50768 = n50685 & ~n50728;
  assign n51143 = n50767 & ~n50768;
  assign n51144 = n51047 ^ n51044;
  assign n51145 = ~n51143 & n51144;
  assign n51146 = n51050 ^ n51042;
  assign n51147 = ~n51145 & n51146;
  assign n51148 = n51053 ^ n51040;
  assign n51149 = ~n51147 & ~n51148;
  assign n51150 = n51142 & n51149;
  assign n51151 = n51059 ^ n51036;
  assign n51152 = n51150 & n51151;
  assign n51153 = n51062 ^ n51034;
  assign n51154 = ~n51152 & ~n51153;
  assign n51155 = ~n51141 & n51154;
  assign n51156 = n51140 & n51155;
  assign n51157 = n51071 ^ n51028;
  assign n51158 = n51156 & n51157;
  assign n51159 = ~n51139 & n51158;
  assign n51160 = n51138 & ~n51159;
  assign n51161 = ~n51137 & n51160;
  assign n51162 = n51083 ^ n51020;
  assign n51163 = ~n51161 & n51162;
  assign n51164 = n51136 & ~n51163;
  assign n51165 = ~n51135 & ~n51164;
  assign n51090 = n51089 ^ n51015;
  assign n51091 = n51016 & n51090;
  assign n51092 = n51091 ^ n48187;
  assign n50946 = n50945 ^ n50942;
  assign n50947 = ~n50943 & ~n50946;
  assign n50948 = n50947 ^ n50945;
  assign n50817 = n50551 ^ n50442;
  assign n50818 = n50817 ^ n50439;
  assign n50815 = n49823 ^ n48778;
  assign n50816 = n50815 ^ n50380;
  assign n50819 = n50818 ^ n50816;
  assign n51013 = n50948 ^ n50819;
  assign n51014 = n51013 ^ n48298;
  assign n51134 = n51092 ^ n51014;
  assign n51342 = n51165 ^ n51134;
  assign n51220 = n49200 ^ n41414;
  assign n51221 = n51220 ^ n45495;
  assign n51222 = n51221 ^ n39853;
  assign n51219 = n51164 ^ n51135;
  assign n51223 = n51222 ^ n51219;
  assign n51331 = n51163 ^ n51136;
  assign n51225 = n49210 ^ n41418;
  assign n51226 = n51225 ^ n45615;
  assign n51227 = n51226 ^ n39863;
  assign n51224 = n51162 ^ n51161;
  assign n51228 = n51227 ^ n51224;
  assign n51230 = n49215 ^ n41530;
  assign n51231 = n51230 ^ n45506;
  assign n51232 = n51231 ^ n39868;
  assign n51229 = n51160 ^ n51137;
  assign n51233 = n51232 ^ n51229;
  assign n51235 = n49220 ^ n41424;
  assign n51236 = n51235 ^ n45604;
  assign n51237 = n51236 ^ n39873;
  assign n51234 = n51159 ^ n51138;
  assign n51238 = n51237 ^ n51234;
  assign n51240 = n49225 ^ n41519;
  assign n51241 = n51240 ^ n45511;
  assign n51242 = n51241 ^ n39965;
  assign n51239 = n51158 ^ n51139;
  assign n51243 = n51242 ^ n51239;
  assign n51311 = n51157 ^ n51156;
  assign n51245 = n49272 ^ n41429;
  assign n51246 = n51245 ^ n1892;
  assign n51247 = n51246 ^ n39879;
  assign n51244 = n51155 ^ n51140;
  assign n51248 = n51247 ^ n51244;
  assign n51252 = n51154 ^ n51141;
  assign n51249 = n49264 ^ n41433;
  assign n51250 = n51249 ^ n45520;
  assign n51251 = n51250 ^ n1881;
  assign n51253 = n51252 ^ n51251;
  assign n51297 = n51153 ^ n51152;
  assign n51255 = n49240 ^ n41438;
  assign n51256 = n51255 ^ n45530;
  assign n51257 = n51256 ^ n39891;
  assign n51254 = n51151 ^ n51150;
  assign n51258 = n51257 ^ n51254;
  assign n51286 = n51149 ^ n51142;
  assign n51260 = n48740 ^ n41449;
  assign n51261 = n51260 ^ n45575;
  assign n51262 = n51261 ^ n39902;
  assign n51259 = n51148 ^ n51147;
  assign n51263 = n51262 ^ n51259;
  assign n51275 = n51146 ^ n51145;
  assign n51265 = n48731 ^ n41459;
  assign n51266 = n51265 ^ n45546;
  assign n51267 = n51266 ^ n39933;
  assign n51264 = n51144 ^ n51143;
  assign n51268 = n51267 ^ n51264;
  assign n50770 = n48721 ^ n41463;
  assign n50771 = n50770 ^ n45559;
  assign n50772 = n50771 ^ n39911;
  assign n50769 = n50768 ^ n50767;
  assign n50773 = n50772 ^ n50769;
  assign n50689 = n48714 ^ n41472;
  assign n50690 = n50689 ^ n45552;
  assign n50691 = n50690 ^ n39920;
  assign n50651 = n48710 ^ n41468;
  assign n50652 = n50651 ^ n2543;
  assign n50653 = n50652 ^ n39915;
  assign n50646 = n50645 ^ n48004;
  assign n50647 = n49354 ^ n41810;
  assign n50648 = n50647 ^ n45895;
  assign n50649 = n50648 ^ n2532;
  assign n50650 = n50646 & n50649;
  assign n50654 = n50653 ^ n50650;
  assign n50686 = n50685 ^ n50650;
  assign n50687 = n50654 & ~n50686;
  assign n50688 = n50687 ^ n50653;
  assign n50692 = n50691 ^ n50688;
  assign n50729 = n50728 ^ n50685;
  assign n50730 = n50729 ^ n50688;
  assign n50731 = n50692 & ~n50730;
  assign n50732 = n50731 ^ n50691;
  assign n51269 = n50769 ^ n50732;
  assign n51270 = ~n50773 & n51269;
  assign n51271 = n51270 ^ n50772;
  assign n51272 = n51271 ^ n51264;
  assign n51273 = n51268 & ~n51272;
  assign n51274 = n51273 ^ n51267;
  assign n51276 = n51275 ^ n51274;
  assign n51277 = n48705 ^ n41454;
  assign n51278 = n51277 ^ n45541;
  assign n51279 = n51278 ^ n39907;
  assign n51280 = n51279 ^ n51275;
  assign n51281 = n51276 & ~n51280;
  assign n51282 = n51281 ^ n51279;
  assign n51283 = n51282 ^ n51259;
  assign n51284 = ~n51263 & n51283;
  assign n51285 = n51284 ^ n51262;
  assign n51287 = n51286 ^ n51285;
  assign n51291 = n51290 ^ n51286;
  assign n51292 = n51287 & ~n51291;
  assign n51293 = n51292 ^ n51290;
  assign n51294 = n51293 ^ n51254;
  assign n51295 = ~n51258 & n51294;
  assign n51296 = n51295 ^ n51257;
  assign n51298 = n51297 ^ n51296;
  assign n51299 = n49234 ^ n1745;
  assign n51300 = n51299 ^ n45525;
  assign n51301 = n51300 ^ n39886;
  assign n51302 = n51301 ^ n51297;
  assign n51303 = ~n51298 & n51302;
  assign n51304 = n51303 ^ n51301;
  assign n51305 = n51304 ^ n51252;
  assign n51306 = ~n51253 & n51305;
  assign n51307 = n51306 ^ n51251;
  assign n51308 = n51307 ^ n51244;
  assign n51309 = n51248 & ~n51308;
  assign n51310 = n51309 ^ n51247;
  assign n51312 = n51311 ^ n51310;
  assign n51313 = n49229 ^ n41511;
  assign n51314 = n51313 ^ n45515;
  assign n51315 = n51314 ^ n2021;
  assign n51316 = n51315 ^ n51311;
  assign n51317 = ~n51312 & n51316;
  assign n51318 = n51317 ^ n51315;
  assign n51319 = n51318 ^ n51239;
  assign n51320 = ~n51243 & n51319;
  assign n51321 = n51320 ^ n51242;
  assign n51322 = n51321 ^ n51234;
  assign n51323 = n51238 & ~n51322;
  assign n51324 = n51323 ^ n51237;
  assign n51325 = n51324 ^ n51229;
  assign n51326 = n51233 & ~n51325;
  assign n51327 = n51326 ^ n51232;
  assign n51328 = n51327 ^ n51224;
  assign n51329 = ~n51228 & n51328;
  assign n51330 = n51329 ^ n51227;
  assign n51332 = n51331 ^ n51330;
  assign n51333 = n49205 ^ n41541;
  assign n51334 = n51333 ^ n45501;
  assign n51335 = n51334 ^ n39857;
  assign n51336 = n51335 ^ n51331;
  assign n51337 = ~n51332 & n51336;
  assign n51338 = n51337 ^ n51335;
  assign n51339 = n51338 ^ n51219;
  assign n51340 = n51223 & ~n51339;
  assign n51341 = n51340 ^ n51222;
  assign n51343 = n51342 ^ n51341;
  assign n51344 = n49195 ^ n41408;
  assign n51345 = n51344 ^ n45491;
  assign n51346 = n51345 ^ n39988;
  assign n51347 = n51346 ^ n51342;
  assign n51348 = n51343 & ~n51347;
  assign n51349 = n51348 ^ n51346;
  assign n51215 = n49190 ^ n41555;
  assign n51216 = n51215 ^ n45486;
  assign n51217 = n51216 ^ n39848;
  assign n51166 = ~n51134 & n51165;
  assign n51093 = n51092 ^ n51013;
  assign n51094 = ~n51014 & ~n51093;
  assign n51095 = n51094 ^ n48298;
  assign n50955 = n50394 ^ n48776;
  assign n50956 = n50955 ^ n49973;
  assign n50952 = n50554 ^ n50437;
  assign n50953 = n50952 ^ n50434;
  assign n50949 = n50948 ^ n50818;
  assign n50950 = n50819 & ~n50949;
  assign n50951 = n50950 ^ n50816;
  assign n50954 = n50953 ^ n50951;
  assign n51011 = n50956 ^ n50954;
  assign n51012 = n51011 ^ n48392;
  assign n51133 = n51095 ^ n51012;
  assign n51214 = n51166 ^ n51133;
  assign n51218 = n51217 ^ n51214;
  assign n51793 = n51349 ^ n51218;
  assign n51708 = n51346 ^ n51343;
  assign n51706 = n50857 ^ n50083;
  assign n51128 = n50596 ^ n50408;
  assign n51707 = n51706 ^ n51128;
  assign n51709 = n51708 ^ n51707;
  assign n51783 = n51338 ^ n51223;
  assign n51776 = n51335 ^ n51332;
  assign n51712 = n51327 ^ n51227;
  assign n51713 = n51712 ^ n51224;
  assign n51710 = n50671 ^ n50003;
  assign n50979 = n50582 ^ n50418;
  assign n51711 = n51710 ^ n50979;
  assign n51714 = n51713 ^ n51711;
  assign n51766 = n51324 ^ n51233;
  assign n51759 = n51321 ^ n51238;
  assign n51752 = n51318 ^ n51243;
  assign n51715 = n50380 ^ n49674;
  assign n50808 = n50565 ^ n50562;
  assign n51716 = n51715 ^ n50808;
  assign n51685 = n51315 ^ n51312;
  assign n51717 = n51716 ^ n51685;
  assign n51720 = n51307 ^ n51248;
  assign n51718 = n50366 ^ n49630;
  assign n50812 = n50557 ^ n50432;
  assign n50813 = n50812 ^ n50429;
  assign n51719 = n51718 ^ n50813;
  assign n51721 = n51720 ^ n51719;
  assign n51724 = n50336 ^ n49685;
  assign n51725 = n51724 ^ n50818;
  assign n51723 = n51301 ^ n51298;
  assign n51726 = n51725 ^ n51723;
  assign n51730 = n51293 ^ n51258;
  assign n51674 = n51290 ^ n51287;
  assign n51672 = n50822 ^ n49637;
  assign n51673 = n51672 ^ n50266;
  assign n51675 = n51674 ^ n51673;
  assign n51549 = n51282 ^ n51263;
  assign n51489 = n50160 ^ n49645;
  assign n51490 = n51489 ^ n50929;
  assign n51488 = n51279 ^ n51276;
  assign n51491 = n51490 ^ n51488;
  assign n51481 = n51271 ^ n51268;
  assign n50775 = n49649 ^ n49634;
  assign n50778 = n50777 ^ n50775;
  assign n50774 = n50773 ^ n50732;
  assign n50779 = n50778 ^ n50774;
  assign n51470 = n50729 ^ n50691;
  assign n51471 = n51470 ^ n50688;
  assign n50784 = n50685 ^ n50653;
  assign n50785 = n50784 ^ n50650;
  assign n50782 = n50781 ^ n49619;
  assign n50783 = n50782 ^ n49641;
  assign n50786 = n50785 ^ n50783;
  assign n50791 = n50649 ^ n50646;
  assign n50789 = n50788 ^ n49485;
  assign n50790 = n50789 ^ n49642;
  assign n50792 = n50791 ^ n50790;
  assign n51403 = n50070 ^ n48750;
  assign n51404 = n51403 ^ n48772;
  assign n50993 = n50593 ^ n50413;
  assign n50986 = n50590 ^ n50587;
  assign n50799 = n50750 ^ n48583;
  assign n50800 = n50799 ^ n49367;
  assign n50798 = n50579 ^ n50423;
  assign n50801 = n50800 ^ n50798;
  assign n50804 = n50576 ^ n50573;
  assign n50802 = n50713 ^ n50083;
  assign n50803 = n50802 ^ n49346;
  assign n50805 = n50804 ^ n50803;
  assign n50966 = n50568 ^ n50428;
  assign n50806 = n50634 ^ n49065;
  assign n50807 = n50806 ^ n50025;
  assign n50809 = n50808 ^ n50807;
  assign n50810 = n50612 ^ n48938;
  assign n50811 = n50810 ^ n50003;
  assign n50814 = n50813 ^ n50811;
  assign n50957 = n50956 ^ n50953;
  assign n50958 = ~n50954 & n50957;
  assign n50959 = n50958 ^ n50956;
  assign n50960 = n50959 ^ n50813;
  assign n50961 = ~n50814 & n50960;
  assign n50962 = n50961 ^ n50811;
  assign n50963 = n50962 ^ n50808;
  assign n50964 = n50809 & ~n50963;
  assign n50965 = n50964 ^ n50807;
  assign n50967 = n50966 ^ n50965;
  assign n50968 = n50056 ^ n49127;
  assign n50969 = n50968 ^ n50671;
  assign n50970 = n50969 ^ n50966;
  assign n50971 = ~n50967 & n50970;
  assign n50972 = n50971 ^ n50969;
  assign n50973 = n50972 ^ n50804;
  assign n50974 = ~n50805 & ~n50973;
  assign n50975 = n50974 ^ n50803;
  assign n50976 = n50975 ^ n50798;
  assign n50977 = n50801 & ~n50976;
  assign n50978 = n50977 ^ n50800;
  assign n50980 = n50979 ^ n50978;
  assign n50981 = n50857 ^ n48580;
  assign n50982 = n50981 ^ n49372;
  assign n50983 = n50982 ^ n50979;
  assign n50984 = n50980 & ~n50983;
  assign n50985 = n50984 ^ n50982;
  assign n50987 = n50986 ^ n50985;
  assign n50988 = n49982 ^ n49379;
  assign n50989 = n50988 ^ n48623;
  assign n50990 = n50989 ^ n50986;
  assign n50991 = n50987 & ~n50990;
  assign n50992 = n50991 ^ n50989;
  assign n50994 = n50993 ^ n50992;
  assign n50796 = n50010 ^ n49362;
  assign n50797 = n50796 ^ n48659;
  assign n51125 = n50993 ^ n50797;
  assign n51126 = n50994 & ~n51125;
  assign n51127 = n51126 ^ n50797;
  assign n51129 = n51128 ^ n51127;
  assign n51123 = n49358 ^ n48694;
  assign n51124 = n51123 ^ n50036;
  assign n51398 = n51128 ^ n51124;
  assign n51399 = ~n51129 & n51398;
  assign n51400 = n51399 ^ n51124;
  assign n51402 = n51401 ^ n51400;
  assign n51405 = n51404 ^ n51402;
  assign n51406 = n51405 ^ n47993;
  assign n51130 = n51129 ^ n51124;
  assign n51131 = n51130 ^ n47960;
  assign n50995 = n50994 ^ n50797;
  assign n50996 = n50995 ^ n47964;
  assign n50997 = n50989 ^ n50987;
  assign n50998 = n50997 ^ n47970;
  assign n50999 = n50982 ^ n50980;
  assign n51000 = n50999 ^ n47980;
  assign n51001 = n50975 ^ n50801;
  assign n51002 = n51001 ^ n47974;
  assign n51003 = n50972 ^ n50805;
  assign n51004 = n51003 ^ n48686;
  assign n51005 = n50969 ^ n50967;
  assign n51006 = n51005 ^ n48647;
  assign n51007 = n50962 ^ n50809;
  assign n51008 = n51007 ^ n48613;
  assign n51009 = n50959 ^ n50814;
  assign n51010 = n51009 ^ n48566;
  assign n51096 = n51095 ^ n51011;
  assign n51097 = n51012 & n51096;
  assign n51098 = n51097 ^ n48392;
  assign n51099 = n51098 ^ n51009;
  assign n51100 = n51010 & n51099;
  assign n51101 = n51100 ^ n48566;
  assign n51102 = n51101 ^ n51007;
  assign n51103 = ~n51008 & n51102;
  assign n51104 = n51103 ^ n48613;
  assign n51105 = n51104 ^ n51005;
  assign n51106 = ~n51006 & n51105;
  assign n51107 = n51106 ^ n48647;
  assign n51108 = n51107 ^ n51003;
  assign n51109 = ~n51004 & ~n51108;
  assign n51110 = n51109 ^ n48686;
  assign n51111 = n51110 ^ n51001;
  assign n51112 = n51002 & n51111;
  assign n51113 = n51112 ^ n47974;
  assign n51114 = n51113 ^ n50999;
  assign n51115 = n51000 & n51114;
  assign n51116 = n51115 ^ n47980;
  assign n51117 = n51116 ^ n50997;
  assign n51118 = ~n50998 & ~n51117;
  assign n51119 = n51118 ^ n47970;
  assign n51120 = n51119 ^ n50995;
  assign n51121 = ~n50996 & n51120;
  assign n51122 = n51121 ^ n47964;
  assign n51395 = n51130 ^ n51122;
  assign n51396 = n51131 & ~n51395;
  assign n51397 = n51396 ^ n47960;
  assign n51407 = n51406 ^ n51397;
  assign n51132 = n51131 ^ n51122;
  assign n51167 = ~n51133 & n51166;
  assign n51168 = n51098 ^ n51010;
  assign n51169 = ~n51167 & ~n51168;
  assign n51170 = n51101 ^ n51008;
  assign n51171 = n51169 & ~n51170;
  assign n51172 = n51104 ^ n51006;
  assign n51173 = ~n51171 & n51172;
  assign n51174 = n51107 ^ n51004;
  assign n51175 = n51173 & n51174;
  assign n51176 = n51110 ^ n51002;
  assign n51177 = ~n51175 & ~n51176;
  assign n51178 = n51113 ^ n51000;
  assign n51179 = ~n51177 & ~n51178;
  assign n51180 = n51116 ^ n50998;
  assign n51181 = ~n51179 & n51180;
  assign n51182 = n51119 ^ n50996;
  assign n51183 = ~n51181 & n51182;
  assign n51408 = ~n51132 & n51183;
  assign n51455 = n51407 & ~n51408;
  assign n51451 = n50095 ^ n48771;
  assign n51446 = n49140 ^ n2405;
  assign n51447 = n51446 ^ n45737;
  assign n51448 = n51447 ^ n40231;
  assign n51449 = n51448 ^ n50854;
  assign n51445 = n50621 ^ n50618;
  assign n51450 = n51449 ^ n51445;
  assign n51452 = n51451 ^ n51450;
  assign n51442 = n51404 ^ n51401;
  assign n51443 = n51402 & ~n51442;
  assign n51444 = n51443 ^ n51404;
  assign n51453 = n51452 ^ n51444;
  assign n51439 = n51405 ^ n51397;
  assign n51440 = n51406 & n51439;
  assign n51441 = n51440 ^ n47993;
  assign n51454 = n51453 ^ n51441;
  assign n51456 = n51455 ^ n51454;
  assign n51409 = n51408 ^ n51407;
  assign n51185 = n41784 ^ n1398;
  assign n51186 = n51185 ^ n45845;
  assign n51187 = n51186 ^ n40241;
  assign n51184 = n51183 ^ n51132;
  assign n51188 = n51187 ^ n51184;
  assign n51384 = n51182 ^ n51181;
  assign n51190 = n49155 ^ n1282;
  assign n51191 = n51190 ^ n45856;
  assign n51192 = n51191 ^ n40245;
  assign n51189 = n51180 ^ n51179;
  assign n51193 = n51192 ^ n51189;
  assign n51194 = n51178 ^ n51177;
  assign n51198 = n51197 ^ n51194;
  assign n51200 = n49165 ^ n41384;
  assign n51201 = n51200 ^ n45866;
  assign n51202 = n51201 ^ n40250;
  assign n51199 = n51176 ^ n51175;
  assign n51203 = n51202 ^ n51199;
  assign n51367 = n51174 ^ n51173;
  assign n51205 = n49175 ^ n41394;
  assign n51206 = n51205 ^ n45662;
  assign n51207 = n51206 ^ n809;
  assign n51204 = n51172 ^ n51171;
  assign n51208 = n51207 ^ n51204;
  assign n51356 = n51170 ^ n51169;
  assign n51210 = n49184 ^ n41404;
  assign n51211 = n51210 ^ n45637;
  assign n51212 = n51211 ^ n39999;
  assign n51209 = n51168 ^ n51167;
  assign n51213 = n51212 ^ n51209;
  assign n51350 = n51349 ^ n51214;
  assign n51351 = ~n51218 & n51350;
  assign n51352 = n51351 ^ n51217;
  assign n51353 = n51352 ^ n51209;
  assign n51354 = ~n51213 & n51353;
  assign n51355 = n51354 ^ n51212;
  assign n51357 = n51356 ^ n51355;
  assign n51358 = n49180 ^ n41398;
  assign n51359 = n51358 ^ n45481;
  assign n51360 = n51359 ^ n39843;
  assign n51361 = n51360 ^ n51356;
  assign n51362 = ~n51357 & n51361;
  assign n51363 = n51362 ^ n51360;
  assign n51364 = n51363 ^ n51204;
  assign n51365 = ~n51208 & n51364;
  assign n51366 = n51365 ^ n51207;
  assign n51368 = n51367 ^ n51366;
  assign n51369 = n49170 ^ n41388;
  assign n51370 = n51369 ^ n45668;
  assign n51371 = n51370 ^ n40260;
  assign n51372 = n51371 ^ n51367;
  assign n51373 = ~n51368 & n51372;
  assign n51374 = n51373 ^ n51371;
  assign n51375 = n51374 ^ n51199;
  assign n51376 = ~n51203 & n51375;
  assign n51377 = n51376 ^ n51202;
  assign n51378 = n51377 ^ n51194;
  assign n51379 = n51198 & ~n51378;
  assign n51380 = n51379 ^ n51197;
  assign n51381 = n51380 ^ n51189;
  assign n51382 = n51193 & ~n51381;
  assign n51383 = n51382 ^ n51192;
  assign n51385 = n51384 ^ n51383;
  assign n51386 = n49149 ^ n1300;
  assign n51387 = n51386 ^ n45850;
  assign n51388 = n51387 ^ n40282;
  assign n51389 = n51388 ^ n51384;
  assign n51390 = n51385 & ~n51389;
  assign n51391 = n51390 ^ n51388;
  assign n51392 = n51391 ^ n51184;
  assign n51393 = ~n51188 & n51392;
  assign n51394 = n51393 ^ n51187;
  assign n51410 = n51409 ^ n51394;
  assign n50793 = n49144 ^ n41779;
  assign n50794 = n50793 ^ n45840;
  assign n50795 = n50794 ^ n40235;
  assign n51436 = n51409 ^ n50795;
  assign n51437 = ~n51410 & n51436;
  assign n51438 = n51437 ^ n50795;
  assign n51457 = n51456 ^ n51438;
  assign n51412 = n49648 ^ n48757;
  assign n51413 = n51412 ^ n50887;
  assign n51411 = n51410 ^ n50795;
  assign n51414 = n51413 ^ n51411;
  assign n51426 = n51391 ^ n51188;
  assign n51417 = n50108 ^ n48765;
  assign n51418 = n51417 ^ n50837;
  assign n51419 = n51380 ^ n51193;
  assign n51420 = ~n51418 & n51419;
  assign n51415 = n50833 ^ n49653;
  assign n51416 = n51415 ^ n49404;
  assign n51421 = n51420 ^ n51416;
  assign n51422 = n51388 ^ n51385;
  assign n51423 = n51422 ^ n51416;
  assign n51424 = n51421 & n51423;
  assign n51425 = n51424 ^ n51420;
  assign n51427 = n51426 ^ n51425;
  assign n51428 = n50118 ^ n48759;
  assign n51429 = n51428 ^ n50879;
  assign n51430 = n51429 ^ n51426;
  assign n51431 = n51427 & n51430;
  assign n51432 = n51431 ^ n51429;
  assign n51433 = n51432 ^ n51411;
  assign n51434 = n51414 & n51433;
  assign n51435 = n51434 ^ n51413;
  assign n51458 = n51457 ^ n51435;
  assign n51459 = n50128 ^ n49419;
  assign n51460 = n51459 ^ n50894;
  assign n51461 = n51460 ^ n51457;
  assign n51462 = ~n51458 & ~n51461;
  assign n51463 = n51462 ^ n51460;
  assign n51464 = n51463 ^ n50791;
  assign n51465 = ~n50792 & n51464;
  assign n51466 = n51465 ^ n50790;
  assign n51467 = n51466 ^ n50785;
  assign n51468 = ~n50786 & n51467;
  assign n51469 = n51468 ^ n50783;
  assign n51472 = n51471 ^ n51469;
  assign n51473 = n49711 ^ n49635;
  assign n51474 = n51473 ^ n50913;
  assign n51475 = n51474 ^ n51471;
  assign n51476 = n51472 & n51475;
  assign n51477 = n51476 ^ n51474;
  assign n51478 = n51477 ^ n50774;
  assign n51479 = n50779 & n51478;
  assign n51480 = n51479 ^ n50778;
  assign n51482 = n51481 ^ n51480;
  assign n51483 = n50828 ^ n49704;
  assign n51484 = n51483 ^ n49633;
  assign n51485 = n51484 ^ n51481;
  assign n51486 = n51482 & n51485;
  assign n51487 = n51486 ^ n51484;
  assign n51546 = n51488 ^ n51487;
  assign n51547 = ~n51491 & n51546;
  assign n51548 = n51547 ^ n51490;
  assign n51550 = n51549 ^ n51548;
  assign n51544 = n49699 ^ n49629;
  assign n51545 = n51544 ^ n50824;
  assign n51669 = n51549 ^ n51545;
  assign n51670 = n51550 & ~n51669;
  assign n51671 = n51670 ^ n51545;
  assign n51727 = n51674 ^ n51671;
  assign n51728 = n51675 & n51727;
  assign n51729 = n51728 ^ n51673;
  assign n51731 = n51730 ^ n51729;
  assign n51732 = n50323 ^ n49689;
  assign n51733 = n51732 ^ n50942;
  assign n51734 = n51733 ^ n51730;
  assign n51735 = ~n51731 & n51734;
  assign n51736 = n51735 ^ n51733;
  assign n51737 = n51736 ^ n51723;
  assign n51738 = ~n51726 & n51737;
  assign n51739 = n51738 ^ n51725;
  assign n51722 = n51304 ^ n51253;
  assign n51740 = n51739 ^ n51722;
  assign n51741 = n50350 ^ n49683;
  assign n51742 = n51741 ^ n50953;
  assign n51743 = n51742 ^ n51722;
  assign n51744 = ~n51740 & n51743;
  assign n51745 = n51744 ^ n51742;
  assign n51746 = n51745 ^ n51720;
  assign n51747 = n51721 & n51746;
  assign n51748 = n51747 ^ n51719;
  assign n51749 = n51748 ^ n51685;
  assign n51750 = n51717 & ~n51749;
  assign n51751 = n51750 ^ n51716;
  assign n51753 = n51752 ^ n51751;
  assign n51754 = n50394 ^ n49751;
  assign n51755 = n51754 ^ n50966;
  assign n51756 = n51755 ^ n51752;
  assign n51757 = n51753 & n51756;
  assign n51758 = n51757 ^ n51755;
  assign n51760 = n51759 ^ n51758;
  assign n51761 = n50612 ^ n49823;
  assign n51762 = n51761 ^ n50804;
  assign n51763 = n51762 ^ n51759;
  assign n51764 = n51760 & n51763;
  assign n51765 = n51764 ^ n51762;
  assign n51767 = n51766 ^ n51765;
  assign n51768 = n50634 ^ n49973;
  assign n51769 = n51768 ^ n50798;
  assign n51770 = n51769 ^ n51766;
  assign n51771 = ~n51767 & ~n51770;
  assign n51772 = n51771 ^ n51769;
  assign n51773 = n51772 ^ n51711;
  assign n51774 = ~n51714 & n51773;
  assign n51775 = n51774 ^ n51713;
  assign n51777 = n51776 ^ n51775;
  assign n51778 = n50713 ^ n50025;
  assign n51779 = n51778 ^ n50986;
  assign n51780 = n51779 ^ n51776;
  assign n51781 = n51777 & n51780;
  assign n51782 = n51781 ^ n51779;
  assign n51784 = n51783 ^ n51782;
  assign n51785 = n50750 ^ n50056;
  assign n51786 = n51785 ^ n50993;
  assign n51787 = n51786 ^ n51783;
  assign n51788 = ~n51784 & ~n51787;
  assign n51789 = n51788 ^ n51786;
  assign n51790 = n51789 ^ n51707;
  assign n51791 = ~n51709 & n51790;
  assign n51792 = n51791 ^ n51708;
  assign n51794 = n51793 ^ n51792;
  assign n51880 = n51796 ^ n51794;
  assign n51817 = n51786 ^ n51784;
  assign n51818 = n51817 ^ n49127;
  assign n51819 = n51779 ^ n51777;
  assign n51820 = n51819 ^ n49065;
  assign n51864 = n51772 ^ n51714;
  assign n51859 = n51769 ^ n51767;
  assign n51821 = n51762 ^ n51760;
  assign n51822 = n51821 ^ n48778;
  assign n51823 = n51755 ^ n51753;
  assign n51824 = n51823 ^ n48780;
  assign n51825 = n51748 ^ n51717;
  assign n51826 = n51825 ^ n48784;
  assign n51827 = n51745 ^ n51721;
  assign n51828 = n51827 ^ n48788;
  assign n51829 = n51742 ^ n51740;
  assign n51830 = n51829 ^ n48794;
  assign n51831 = n51736 ^ n51726;
  assign n51832 = n51831 ^ n48799;
  assign n51833 = n51733 ^ n51731;
  assign n51834 = n51833 ^ n48804;
  assign n51676 = n51675 ^ n51671;
  assign n51677 = n51676 ^ n48808;
  assign n51551 = n51550 ^ n51545;
  assign n51552 = n51551 ^ n48812;
  assign n51492 = n51491 ^ n51487;
  assign n51493 = n51492 ^ n48893;
  assign n51494 = n51484 ^ n51482;
  assign n51495 = n51494 ^ n48816;
  assign n51496 = n51477 ^ n50779;
  assign n51497 = n51496 ^ n48180;
  assign n51498 = n51474 ^ n51472;
  assign n51499 = n51498 ^ n48760;
  assign n51500 = n51466 ^ n50786;
  assign n51501 = n51500 ^ n48823;
  assign n51502 = n51463 ^ n50792;
  assign n51503 = n51502 ^ n48766;
  assign n51504 = n51460 ^ n51458;
  assign n51505 = n51504 ^ n48828;
  assign n51506 = n51432 ^ n51414;
  assign n51507 = n51506 ^ n48829;
  assign n51508 = n51429 ^ n51427;
  assign n51509 = n51508 ^ n48773;
  assign n51510 = n51419 ^ n51418;
  assign n51511 = ~n48835 & ~n51510;
  assign n51512 = n51511 ^ n48852;
  assign n51513 = n51422 ^ n51421;
  assign n51514 = n51513 ^ n51511;
  assign n51515 = n51512 & n51514;
  assign n51516 = n51515 ^ n48852;
  assign n51517 = n51516 ^ n51508;
  assign n51518 = ~n51509 & ~n51517;
  assign n51519 = n51518 ^ n48773;
  assign n51520 = n51519 ^ n51506;
  assign n51521 = n51507 & ~n51520;
  assign n51522 = n51521 ^ n48829;
  assign n51523 = n51522 ^ n51504;
  assign n51524 = ~n51505 & ~n51523;
  assign n51525 = n51524 ^ n48828;
  assign n51526 = n51525 ^ n51502;
  assign n51527 = ~n51503 & ~n51526;
  assign n51528 = n51527 ^ n48766;
  assign n51529 = n51528 ^ n51500;
  assign n51530 = n51501 & n51529;
  assign n51531 = n51530 ^ n48823;
  assign n51532 = n51531 ^ n51498;
  assign n51533 = n51499 & n51532;
  assign n51534 = n51533 ^ n48760;
  assign n51535 = n51534 ^ n51496;
  assign n51536 = n51497 & n51535;
  assign n51537 = n51536 ^ n48180;
  assign n51538 = n51537 ^ n51494;
  assign n51539 = n51495 & n51538;
  assign n51540 = n51539 ^ n48816;
  assign n51541 = n51540 ^ n51492;
  assign n51542 = n51493 & ~n51541;
  assign n51543 = n51542 ^ n48893;
  assign n51666 = n51551 ^ n51543;
  assign n51667 = ~n51552 & ~n51666;
  assign n51668 = n51667 ^ n48812;
  assign n51835 = n51676 ^ n51668;
  assign n51836 = n51677 & ~n51835;
  assign n51837 = n51836 ^ n48808;
  assign n51838 = n51837 ^ n51833;
  assign n51839 = ~n51834 & n51838;
  assign n51840 = n51839 ^ n48804;
  assign n51841 = n51840 ^ n51831;
  assign n51842 = ~n51832 & ~n51841;
  assign n51843 = n51842 ^ n48799;
  assign n51844 = n51843 ^ n51829;
  assign n51845 = ~n51830 & ~n51844;
  assign n51846 = n51845 ^ n48794;
  assign n51847 = n51846 ^ n51827;
  assign n51848 = n51828 & n51847;
  assign n51849 = n51848 ^ n48788;
  assign n51850 = n51849 ^ n51825;
  assign n51851 = ~n51826 & n51850;
  assign n51852 = n51851 ^ n48784;
  assign n51853 = n51852 ^ n51823;
  assign n51854 = n51824 & n51853;
  assign n51855 = n51854 ^ n48780;
  assign n51856 = n51855 ^ n51821;
  assign n51857 = n51822 & n51856;
  assign n51858 = n51857 ^ n48778;
  assign n51860 = n51859 ^ n51858;
  assign n51861 = n51859 ^ n48776;
  assign n51862 = ~n51860 & n51861;
  assign n51863 = n51862 ^ n48776;
  assign n51865 = n51864 ^ n51863;
  assign n51866 = n51864 ^ n48938;
  assign n51867 = n51865 & n51866;
  assign n51868 = n51867 ^ n48938;
  assign n51869 = n51868 ^ n51819;
  assign n51870 = n51820 & n51869;
  assign n51871 = n51870 ^ n49065;
  assign n51872 = n51871 ^ n51817;
  assign n51873 = n51818 & ~n51872;
  assign n51874 = n51873 ^ n49127;
  assign n51875 = n51874 ^ n49346;
  assign n51876 = n51789 ^ n51709;
  assign n51877 = n51876 ^ n51874;
  assign n51878 = n51875 & n51877;
  assign n51879 = n51878 ^ n49346;
  assign n51881 = n51880 ^ n51879;
  assign n51938 = n51881 ^ n48583;
  assign n51912 = n51876 ^ n51875;
  assign n51913 = n51871 ^ n51818;
  assign n51914 = n51868 ^ n49065;
  assign n51915 = n51914 ^ n51819;
  assign n51916 = n51865 ^ n48938;
  assign n51917 = n51855 ^ n51822;
  assign n51918 = n51849 ^ n51826;
  assign n51919 = n51843 ^ n51830;
  assign n51920 = n51840 ^ n51832;
  assign n51553 = n51552 ^ n51543;
  assign n51554 = n51540 ^ n51493;
  assign n51555 = n51531 ^ n51499;
  assign n51556 = n51528 ^ n51501;
  assign n51557 = n51525 ^ n51503;
  assign n51558 = n51516 ^ n51509;
  assign n51559 = n51513 ^ n51512;
  assign n51560 = n51558 & n51559;
  assign n51561 = n51519 ^ n51507;
  assign n51562 = ~n51560 & ~n51561;
  assign n51563 = n51522 ^ n51505;
  assign n51564 = ~n51562 & ~n51563;
  assign n51565 = ~n51557 & ~n51564;
  assign n51566 = n51556 & ~n51565;
  assign n51567 = ~n51555 & n51566;
  assign n51568 = n51534 ^ n51497;
  assign n51569 = n51567 & n51568;
  assign n51570 = n51537 ^ n51495;
  assign n51571 = ~n51569 & n51570;
  assign n51572 = ~n51554 & n51571;
  assign n51665 = n51553 & n51572;
  assign n51678 = n51677 ^ n51668;
  assign n51921 = n51665 & n51678;
  assign n51922 = n51837 ^ n51834;
  assign n51923 = n51921 & ~n51922;
  assign n51924 = n51920 & ~n51923;
  assign n51925 = ~n51919 & n51924;
  assign n51926 = n51846 ^ n51828;
  assign n51927 = ~n51925 & n51926;
  assign n51928 = ~n51918 & ~n51927;
  assign n51929 = n51852 ^ n51824;
  assign n51930 = ~n51928 & ~n51929;
  assign n51931 = n51917 & n51930;
  assign n51932 = n51860 ^ n48776;
  assign n51933 = n51931 & ~n51932;
  assign n51934 = n51916 & ~n51933;
  assign n51935 = ~n51915 & n51934;
  assign n51936 = ~n51913 & ~n51935;
  assign n51937 = n51912 & n51936;
  assign n52064 = n51938 ^ n51937;
  assign n51969 = n49877 ^ n869;
  assign n51970 = n51969 ^ n46518;
  assign n51971 = n51970 ^ n40995;
  assign n51968 = n51936 ^ n51912;
  assign n51972 = n51971 ^ n51968;
  assign n51976 = n51935 ^ n51913;
  assign n51973 = n49882 ^ n42099;
  assign n51974 = n51973 ^ n46522;
  assign n51975 = n51974 ^ n41000;
  assign n51977 = n51976 ^ n51975;
  assign n51979 = n49887 ^ n42104;
  assign n51980 = n51979 ^ n46528;
  assign n51981 = n51980 ^ n41005;
  assign n51978 = n51934 ^ n51915;
  assign n51982 = n51981 ^ n51978;
  assign n51984 = n49892 ^ n42109;
  assign n51985 = n51984 ^ n46545;
  assign n51986 = n51985 ^ n41030;
  assign n51983 = n51933 ^ n51916;
  assign n51987 = n51986 ^ n51983;
  assign n51991 = n51932 ^ n51931;
  assign n51988 = n49896 ^ n42114;
  assign n51989 = n51988 ^ n46532;
  assign n51990 = n51989 ^ n41009;
  assign n51992 = n51991 ^ n51990;
  assign n52041 = n51930 ^ n51917;
  assign n51994 = n49907 ^ n42118;
  assign n51995 = n51994 ^ n46115;
  assign n51996 = n51995 ^ n40654;
  assign n51993 = n51929 ^ n51928;
  assign n51997 = n51996 ^ n51993;
  assign n51999 = n49912 ^ n42240;
  assign n52000 = n51999 ^ n46242;
  assign n52001 = n52000 ^ n40512;
  assign n51998 = n51927 ^ n51918;
  assign n52002 = n52001 ^ n51998;
  assign n52004 = n49926 ^ n42229;
  assign n52005 = n52004 ^ n46124;
  assign n52006 = n52005 ^ n40625;
  assign n52003 = n51924 ^ n51919;
  assign n52007 = n52006 ^ n52003;
  assign n52009 = n49627 ^ n42129;
  assign n52010 = n52009 ^ n46130;
  assign n52011 = n52010 ^ n40522;
  assign n52008 = n51923 ^ n51920;
  assign n52012 = n52011 ^ n52008;
  assign n52013 = n51922 ^ n51921;
  assign n2112 = n2111 ^ n2066;
  assign n2149 = n2148 ^ n2112;
  assign n2159 = n2158 ^ n2149;
  assign n52014 = n52013 ^ n2159;
  assign n51680 = n49518 ^ n42133;
  assign n51681 = n51680 ^ n46137;
  assign n51682 = n51681 ^ n2140;
  assign n51679 = n51678 ^ n51665;
  assign n51683 = n51682 ^ n51679;
  assign n51574 = n49598 ^ n46142;
  assign n51575 = n51574 ^ n1965;
  assign n51576 = n51575 ^ n40529;
  assign n51573 = n51572 ^ n51553;
  assign n51577 = n51576 ^ n51573;
  assign n51579 = n49523 ^ n42140;
  assign n51580 = n51579 ^ n46146;
  assign n51581 = n51580 ^ n40534;
  assign n51578 = n51571 ^ n51554;
  assign n51582 = n51581 ^ n51578;
  assign n51651 = n51570 ^ n51569;
  assign n51584 = n49533 ^ n42146;
  assign n51585 = n51584 ^ n46156;
  assign n51586 = n51585 ^ n40538;
  assign n51583 = n51568 ^ n51567;
  assign n51587 = n51586 ^ n51583;
  assign n51640 = n51566 ^ n51555;
  assign n51589 = n49580 ^ n42156;
  assign n51590 = n51589 ^ n46166;
  assign n51591 = n51590 ^ n40548;
  assign n51588 = n51565 ^ n51556;
  assign n51592 = n51591 ^ n51588;
  assign n51629 = n51564 ^ n51557;
  assign n51594 = n49569 ^ n42184;
  assign n51595 = n51594 ^ n46193;
  assign n51596 = n51595 ^ n40580;
  assign n51593 = n51563 ^ n51562;
  assign n51597 = n51596 ^ n51593;
  assign n51599 = n49561 ^ n42165;
  assign n51600 = n51599 ^ n46172;
  assign n51601 = n51600 ^ n40558;
  assign n51598 = n51561 ^ n51560;
  assign n51602 = n51601 ^ n51598;
  assign n51604 = n49552 ^ n42171;
  assign n51605 = n51604 ^ n46181;
  assign n51606 = n51605 ^ n40562;
  assign n51603 = n51559 ^ n51558;
  assign n51607 = n51606 ^ n51603;
  assign n51613 = n49547 ^ n2610;
  assign n51614 = n51613 ^ n46176;
  assign n51615 = n51614 ^ n40565;
  assign n51608 = n50088 ^ n42523;
  assign n51609 = n51608 ^ n46613;
  assign n51610 = n51609 ^ n40771;
  assign n51611 = n51510 ^ n48835;
  assign n51612 = n51610 & n51611;
  assign n51616 = n51615 ^ n51612;
  assign n51617 = n51612 ^ n51559;
  assign n51618 = n51616 & ~n51617;
  assign n51619 = n51618 ^ n51615;
  assign n51620 = n51619 ^ n51603;
  assign n51621 = ~n51607 & n51620;
  assign n51622 = n51621 ^ n51606;
  assign n51623 = n51622 ^ n51598;
  assign n51624 = n51602 & ~n51623;
  assign n51625 = n51624 ^ n51601;
  assign n51626 = n51625 ^ n51593;
  assign n51627 = ~n51597 & n51626;
  assign n51628 = n51627 ^ n51596;
  assign n51630 = n51629 ^ n51628;
  assign n51631 = n49543 ^ n42161;
  assign n51632 = n51631 ^ n46201;
  assign n51633 = n51632 ^ n40553;
  assign n51634 = n51633 ^ n51629;
  assign n51635 = ~n51630 & n51634;
  assign n51636 = n51635 ^ n51633;
  assign n51637 = n51636 ^ n51588;
  assign n51638 = n51592 & ~n51637;
  assign n51639 = n51638 ^ n51591;
  assign n51641 = n51640 ^ n51639;
  assign n51642 = n49538 ^ n42151;
  assign n51643 = n51642 ^ n46162;
  assign n51644 = n51643 ^ n40544;
  assign n51645 = n51644 ^ n51640;
  assign n51646 = ~n51641 & n51645;
  assign n51647 = n51646 ^ n51644;
  assign n51648 = n51647 ^ n51583;
  assign n51649 = ~n51587 & n51648;
  assign n51650 = n51649 ^ n51586;
  assign n51652 = n51651 ^ n51650;
  assign n51653 = n49528 ^ n42204;
  assign n51654 = n51653 ^ n46151;
  assign n51655 = n51654 ^ n40600;
  assign n51656 = n51655 ^ n51651;
  assign n51657 = n51652 & ~n51656;
  assign n51658 = n51657 ^ n51655;
  assign n51659 = n51658 ^ n51578;
  assign n51660 = ~n51582 & n51659;
  assign n51661 = n51660 ^ n51581;
  assign n51662 = n51661 ^ n51573;
  assign n51663 = n51577 & ~n51662;
  assign n51664 = n51663 ^ n51576;
  assign n52015 = n51679 ^ n51664;
  assign n52016 = n51683 & ~n52015;
  assign n52017 = n52016 ^ n51682;
  assign n52018 = n52017 ^ n2159;
  assign n52019 = ~n52014 & ~n52018;
  assign n52020 = n52019 ^ n52013;
  assign n52021 = n52020 ^ n52008;
  assign n52022 = n52012 & n52021;
  assign n52023 = n52022 ^ n52011;
  assign n52024 = n52023 ^ n52003;
  assign n52025 = n52007 & ~n52024;
  assign n52026 = n52025 ^ n52006;
  assign n52030 = n52029 ^ n52026;
  assign n52031 = n51926 ^ n51925;
  assign n52032 = n52031 ^ n52026;
  assign n52033 = n52030 & n52032;
  assign n52034 = n52033 ^ n52029;
  assign n52035 = n52034 ^ n51998;
  assign n52036 = ~n52002 & n52035;
  assign n52037 = n52036 ^ n52001;
  assign n52038 = n52037 ^ n51993;
  assign n52039 = n51997 & ~n52038;
  assign n52040 = n52039 ^ n51996;
  assign n52042 = n52041 ^ n52040;
  assign n52043 = n49902 ^ n42251;
  assign n52044 = n52043 ^ n46269;
  assign n52045 = n52044 ^ n41015;
  assign n52046 = n52045 ^ n52041;
  assign n52047 = ~n52042 & n52046;
  assign n52048 = n52047 ^ n52045;
  assign n52049 = n52048 ^ n51990;
  assign n52050 = ~n51992 & ~n52049;
  assign n52051 = n52050 ^ n51991;
  assign n52052 = n52051 ^ n51983;
  assign n52053 = n51987 & n52052;
  assign n52054 = n52053 ^ n51986;
  assign n52055 = n52054 ^ n51978;
  assign n52056 = n51982 & ~n52055;
  assign n52057 = n52056 ^ n51981;
  assign n52058 = n52057 ^ n51975;
  assign n52059 = n51977 & ~n52058;
  assign n52060 = n52059 ^ n51976;
  assign n52061 = n52060 ^ n51968;
  assign n52062 = n51972 & ~n52061;
  assign n52063 = n52062 ^ n51971;
  assign n52065 = n52064 ^ n52063;
  assign n52066 = n49871 ^ n42437;
  assign n52067 = n52066 ^ n46513;
  assign n52068 = n52067 ^ n1011;
  assign n52069 = n52068 ^ n52064;
  assign n52070 = n52065 & ~n52069;
  assign n52071 = n52070 ^ n52068;
  assign n51939 = ~n51937 & ~n51938;
  assign n51882 = n51880 ^ n48583;
  assign n51883 = ~n51881 & ~n51882;
  assign n51884 = n51883 ^ n48583;
  assign n51910 = n51884 ^ n48580;
  assign n51797 = n51796 ^ n51793;
  assign n51798 = ~n51794 & n51797;
  assign n51799 = n51798 ^ n51796;
  assign n51704 = n51352 ^ n51213;
  assign n51702 = n50010 ^ n49372;
  assign n51703 = n51702 ^ n51445;
  assign n51705 = n51704 ^ n51703;
  assign n51815 = n51799 ^ n51705;
  assign n51911 = n51910 ^ n51815;
  assign n51966 = n51939 ^ n51911;
  assign n51963 = n49867 ^ n42449;
  assign n51964 = n51963 ^ n1022;
  assign n51965 = n51964 ^ n41050;
  assign n51967 = n51966 ^ n51965;
  assign n52873 = n52071 ^ n51967;
  assign n52930 = n52873 ^ n50681;
  assign n52931 = n52930 ^ n51422;
  assign n52350 = n50813 ^ n50336;
  assign n52351 = n52350 ^ n51759;
  assign n52349 = n51655 ^ n51652;
  assign n52352 = n52351 ^ n52349;
  assign n52354 = n50953 ^ n50323;
  assign n52355 = n52354 ^ n51752;
  assign n52353 = n51647 ^ n51587;
  assign n52356 = n52355 ^ n52353;
  assign n52358 = n50818 ^ n50266;
  assign n52359 = n52358 ^ n51685;
  assign n52357 = n51644 ^ n51641;
  assign n52360 = n52359 ^ n52357;
  assign n52362 = n50942 ^ n49629;
  assign n52363 = n52362 ^ n51720;
  assign n52361 = n51636 ^ n51592;
  assign n52364 = n52363 ^ n52361;
  assign n52318 = n50822 ^ n50160;
  assign n52319 = n52318 ^ n51722;
  assign n52317 = n51633 ^ n51630;
  assign n52320 = n52319 ^ n52317;
  assign n52211 = n51625 ^ n51597;
  assign n52208 = n50824 ^ n49633;
  assign n52209 = n52208 ^ n51723;
  assign n52313 = n52211 ^ n52209;
  assign n52197 = n50929 ^ n49634;
  assign n52198 = n52197 ^ n51730;
  assign n52196 = n51622 ^ n51602;
  assign n52199 = n52198 ^ n52196;
  assign n52185 = n50828 ^ n49635;
  assign n52186 = n52185 ^ n51674;
  assign n52184 = n51619 ^ n51607;
  assign n52187 = n52186 ^ n52184;
  assign n52146 = n51615 ^ n51559;
  assign n52147 = n52146 ^ n51612;
  assign n52139 = n51611 ^ n51610;
  assign n52107 = n50781 ^ n50128;
  assign n52108 = n52107 ^ n51481;
  assign n52101 = n50052 ^ n42477;
  assign n52102 = n52101 ^ n46594;
  assign n52103 = n52102 ^ n40976;
  assign n51809 = n51371 ^ n51368;
  assign n51696 = n51363 ^ n51208;
  assign n51694 = n50070 ^ n49362;
  assign n51695 = n51694 ^ n50681;
  assign n51697 = n51696 ^ n51695;
  assign n51700 = n51360 ^ n51357;
  assign n51698 = n50036 ^ n49379;
  assign n51699 = n51698 ^ n50642;
  assign n51701 = n51700 ^ n51699;
  assign n51800 = n51799 ^ n51703;
  assign n51801 = n51705 & ~n51800;
  assign n51802 = n51801 ^ n51704;
  assign n51803 = n51802 ^ n51699;
  assign n51804 = n51701 & n51803;
  assign n51805 = n51804 ^ n51700;
  assign n51806 = n51805 ^ n51696;
  assign n51807 = n51697 & n51806;
  assign n51808 = n51807 ^ n51695;
  assign n51810 = n51809 ^ n51808;
  assign n51692 = n50095 ^ n49358;
  assign n51693 = n51692 ^ n50724;
  assign n51903 = n51809 ^ n51693;
  assign n51904 = n51810 & ~n51903;
  assign n51905 = n51904 ^ n51693;
  assign n51900 = n49664 ^ n48772;
  assign n51901 = n51900 ^ n50763;
  assign n51899 = n51374 ^ n51203;
  assign n51902 = n51901 ^ n51899;
  assign n51906 = n51905 ^ n51902;
  assign n51907 = n51906 ^ n48750;
  assign n51811 = n51810 ^ n51693;
  assign n51812 = n51811 ^ n48694;
  assign n51813 = n51805 ^ n51697;
  assign n51814 = n51813 ^ n48659;
  assign n51888 = n51802 ^ n51701;
  assign n51816 = n51815 ^ n48580;
  assign n51885 = n51884 ^ n51815;
  assign n51886 = n51816 & n51885;
  assign n51887 = n51886 ^ n48580;
  assign n51889 = n51888 ^ n51887;
  assign n51890 = n51887 ^ n48623;
  assign n51891 = ~n51889 & n51890;
  assign n51892 = n51891 ^ n48623;
  assign n51893 = n51892 ^ n51813;
  assign n51894 = n51814 & n51893;
  assign n51895 = n51894 ^ n48659;
  assign n51896 = n51895 ^ n51811;
  assign n51897 = ~n51812 & ~n51896;
  assign n51898 = n51897 ^ n48694;
  assign n51908 = n51907 ^ n51898;
  assign n51909 = n51895 ^ n51812;
  assign n51940 = n51911 & ~n51939;
  assign n51941 = n51889 ^ n48623;
  assign n51942 = ~n51940 & n51941;
  assign n51943 = n51892 ^ n51814;
  assign n51944 = ~n51942 & ~n51943;
  assign n51945 = ~n51909 & n51944;
  assign n52100 = n51908 & ~n51945;
  assign n52104 = n52103 ^ n52100;
  assign n52094 = n49660 ^ n48771;
  assign n52095 = n52094 ^ n50866;
  assign n52091 = n51905 ^ n51901;
  assign n52092 = ~n51902 & n52091;
  assign n52093 = n52092 ^ n51905;
  assign n52096 = n52095 ^ n52093;
  assign n52090 = n51377 ^ n51198;
  assign n52097 = n52096 ^ n52090;
  assign n52087 = n51906 ^ n51898;
  assign n52088 = n51907 & ~n52087;
  assign n52089 = n52088 ^ n48750;
  assign n52098 = n52097 ^ n52089;
  assign n52099 = n52098 ^ n48840;
  assign n52105 = n52104 ^ n52099;
  assign n51946 = n51945 ^ n51908;
  assign n51689 = n50019 ^ n42427;
  assign n51690 = n51689 ^ n46491;
  assign n51691 = n51690 ^ n40981;
  assign n51947 = n51946 ^ n51691;
  assign n51951 = n51944 ^ n51909;
  assign n51948 = n49989 ^ n42468;
  assign n51949 = n51948 ^ n46495;
  assign n51950 = n51949 ^ n41064;
  assign n51952 = n51951 ^ n51950;
  assign n51956 = n51943 ^ n51942;
  assign n51953 = n49670 ^ n42460;
  assign n51954 = n51953 ^ n46501;
  assign n51955 = n51954 ^ n40985;
  assign n51957 = n51956 ^ n51955;
  assign n51961 = n51941 ^ n51940;
  assign n51958 = n49862 ^ n42432;
  assign n51959 = n51958 ^ n46506;
  assign n51960 = n51959 ^ n1154;
  assign n51962 = n51961 ^ n51960;
  assign n52072 = n52071 ^ n51965;
  assign n52073 = ~n51967 & ~n52072;
  assign n52074 = n52073 ^ n51966;
  assign n52075 = n52074 ^ n51960;
  assign n52076 = n51962 & n52075;
  assign n52077 = n52076 ^ n51961;
  assign n52078 = n52077 ^ n51955;
  assign n52079 = n51957 & ~n52078;
  assign n52080 = n52079 ^ n51956;
  assign n52081 = n52080 ^ n51951;
  assign n52082 = ~n51952 & n52081;
  assign n52083 = n52082 ^ n51950;
  assign n52084 = n52083 ^ n51691;
  assign n52085 = n51947 & ~n52084;
  assign n52086 = n52085 ^ n51946;
  assign n52106 = n52105 ^ n52086;
  assign n52109 = n52108 ^ n52106;
  assign n52129 = n50788 ^ n49648;
  assign n52130 = n52129 ^ n50774;
  assign n52112 = n50894 ^ n50118;
  assign n52113 = n52112 ^ n51471;
  assign n52110 = n52080 ^ n51950;
  assign n52111 = n52110 ^ n51951;
  assign n52114 = n52113 ^ n52111;
  assign n52117 = n52074 ^ n51962;
  assign n52118 = n50879 ^ n50108;
  assign n52119 = n52118 ^ n50791;
  assign n52120 = ~n52117 & n52119;
  assign n52115 = n50887 ^ n49653;
  assign n52116 = n52115 ^ n50785;
  assign n52121 = n52120 ^ n52116;
  assign n52122 = n52077 ^ n51957;
  assign n52123 = n52122 ^ n52116;
  assign n52124 = ~n52121 & n52123;
  assign n52125 = n52124 ^ n52120;
  assign n52126 = n52125 ^ n52111;
  assign n52127 = ~n52114 & n52126;
  assign n52128 = n52127 ^ n52113;
  assign n52131 = n52130 ^ n52128;
  assign n52132 = n52083 ^ n51947;
  assign n52133 = n52132 ^ n52128;
  assign n52134 = ~n52131 & ~n52133;
  assign n52135 = n52134 ^ n52130;
  assign n52136 = n52135 ^ n52106;
  assign n52137 = n52109 & n52136;
  assign n52138 = n52137 ^ n52108;
  assign n52140 = n52139 ^ n52138;
  assign n52141 = n50913 ^ n49642;
  assign n52142 = n52141 ^ n51488;
  assign n52143 = n52142 ^ n52139;
  assign n52144 = ~n52140 & ~n52143;
  assign n52145 = n52144 ^ n52142;
  assign n52148 = n52147 ^ n52145;
  assign n51687 = n50777 ^ n49641;
  assign n51688 = n51687 ^ n51549;
  assign n52181 = n52147 ^ n51688;
  assign n52182 = n52148 & ~n52181;
  assign n52183 = n52182 ^ n51688;
  assign n52193 = n52184 ^ n52183;
  assign n52194 = ~n52187 & ~n52193;
  assign n52195 = n52194 ^ n52186;
  assign n52205 = n52196 ^ n52195;
  assign n52206 = n52199 & ~n52205;
  assign n52207 = n52206 ^ n52198;
  assign n52314 = n52211 ^ n52207;
  assign n52315 = ~n52313 & n52314;
  assign n52316 = n52315 ^ n52209;
  assign n52365 = n52319 ^ n52316;
  assign n52366 = ~n52320 & n52365;
  assign n52367 = n52366 ^ n52317;
  assign n52368 = n52367 ^ n52361;
  assign n52369 = ~n52364 & ~n52368;
  assign n52370 = n52369 ^ n52363;
  assign n52371 = n52370 ^ n52359;
  assign n52372 = ~n52360 & ~n52371;
  assign n52373 = n52372 ^ n52357;
  assign n52374 = n52373 ^ n52353;
  assign n52375 = n52356 & n52374;
  assign n52376 = n52375 ^ n52355;
  assign n52377 = n52376 ^ n52349;
  assign n52378 = n52352 & ~n52377;
  assign n52379 = n52378 ^ n52351;
  assign n52345 = n50808 ^ n50350;
  assign n52346 = n52345 ^ n51766;
  assign n52403 = n52379 ^ n52346;
  assign n52347 = n51658 ^ n51582;
  assign n52404 = n52403 ^ n52347;
  assign n52405 = n52404 ^ n49683;
  assign n52406 = n52376 ^ n52352;
  assign n52407 = n52406 ^ n49685;
  assign n52408 = n52373 ^ n52356;
  assign n52409 = n52408 ^ n49689;
  assign n52410 = n52367 ^ n52364;
  assign n52411 = n52410 ^ n49699;
  assign n52210 = n52209 ^ n52207;
  assign n52212 = n52211 ^ n52210;
  assign n52213 = n52212 ^ n49704;
  assign n52200 = n52199 ^ n52195;
  assign n52188 = n52187 ^ n52183;
  assign n52149 = n52148 ^ n51688;
  assign n52150 = n52149 ^ n49619;
  assign n52173 = n52142 ^ n52140;
  assign n52151 = n52135 ^ n52109;
  assign n52152 = n52151 ^ n49419;
  assign n52153 = n52132 ^ n52131;
  assign n52154 = n52153 ^ n48757;
  assign n52155 = n52125 ^ n52114;
  assign n52156 = n52155 ^ n48759;
  assign n52157 = n52119 ^ n52117;
  assign n52158 = n48765 & ~n52157;
  assign n52159 = n52158 ^ n49404;
  assign n52160 = n52122 ^ n52121;
  assign n52161 = n52160 ^ n52158;
  assign n52162 = ~n52159 & n52161;
  assign n52163 = n52162 ^ n49404;
  assign n52164 = n52163 ^ n52155;
  assign n52165 = n52156 & ~n52164;
  assign n52166 = n52165 ^ n48759;
  assign n52167 = n52166 ^ n52153;
  assign n52168 = n52154 & ~n52167;
  assign n52169 = n52168 ^ n48757;
  assign n52170 = n52169 ^ n52151;
  assign n52171 = ~n52152 & ~n52170;
  assign n52172 = n52171 ^ n49419;
  assign n52174 = n52173 ^ n52172;
  assign n52175 = n52173 ^ n49485;
  assign n52176 = n52174 & ~n52175;
  assign n52177 = n52176 ^ n49485;
  assign n52178 = n52177 ^ n52149;
  assign n52179 = n52150 & ~n52178;
  assign n52180 = n52179 ^ n49619;
  assign n52189 = n52188 ^ n52180;
  assign n52190 = n52188 ^ n49711;
  assign n52191 = ~n52189 & n52190;
  assign n52192 = n52191 ^ n49711;
  assign n52201 = n52200 ^ n52192;
  assign n52202 = n52200 ^ n49649;
  assign n52203 = ~n52201 & n52202;
  assign n52204 = n52203 ^ n49649;
  assign n52323 = n52212 ^ n52204;
  assign n52324 = ~n52213 & n52323;
  assign n52325 = n52324 ^ n49704;
  assign n52412 = n52325 ^ n49645;
  assign n52321 = n52320 ^ n52316;
  assign n52413 = n52325 ^ n52321;
  assign n52414 = ~n52412 & n52413;
  assign n52415 = n52414 ^ n49645;
  assign n52416 = n52415 ^ n52410;
  assign n52417 = n52411 & ~n52416;
  assign n52418 = n52417 ^ n49699;
  assign n52419 = n52418 ^ n49637;
  assign n52420 = n52370 ^ n52360;
  assign n52421 = n52420 ^ n52418;
  assign n52422 = n52419 & n52421;
  assign n52423 = n52422 ^ n49637;
  assign n52424 = n52423 ^ n52408;
  assign n52425 = n52409 & n52424;
  assign n52426 = n52425 ^ n49689;
  assign n52427 = n52426 ^ n52406;
  assign n52428 = n52407 & n52427;
  assign n52429 = n52428 ^ n49685;
  assign n52430 = n52429 ^ n52404;
  assign n52431 = ~n52405 & n52430;
  assign n52432 = n52431 ^ n49683;
  assign n52348 = n52347 ^ n52346;
  assign n52380 = n52379 ^ n52347;
  assign n52381 = ~n52348 & ~n52380;
  assign n52382 = n52381 ^ n52346;
  assign n52343 = n51661 ^ n51577;
  assign n52341 = n50966 ^ n50366;
  assign n52342 = n52341 ^ n51713;
  assign n52344 = n52343 ^ n52342;
  assign n52401 = n52382 ^ n52344;
  assign n52402 = n52401 ^ n49630;
  assign n52471 = n52432 ^ n52402;
  assign n52472 = n52429 ^ n52405;
  assign n52473 = n52426 ^ n49685;
  assign n52474 = n52473 ^ n52406;
  assign n52475 = n52423 ^ n49689;
  assign n52476 = n52475 ^ n52408;
  assign n52322 = n52321 ^ n49645;
  assign n52326 = n52325 ^ n52322;
  assign n52214 = n52213 ^ n52204;
  assign n52215 = n52160 ^ n52159;
  assign n52216 = n52163 ^ n48759;
  assign n52217 = n52216 ^ n52155;
  assign n52218 = ~n52215 & n52217;
  assign n52219 = n52166 ^ n52154;
  assign n52220 = ~n52218 & ~n52219;
  assign n52221 = n52169 ^ n49419;
  assign n52222 = n52221 ^ n52151;
  assign n52223 = ~n52220 & ~n52222;
  assign n52224 = n52174 ^ n49485;
  assign n52225 = ~n52223 & ~n52224;
  assign n52226 = n52177 ^ n49619;
  assign n52227 = n52226 ^ n52149;
  assign n52228 = ~n52225 & ~n52227;
  assign n52229 = n52189 ^ n49711;
  assign n52230 = n52228 & ~n52229;
  assign n52231 = n52201 ^ n49649;
  assign n52232 = n52230 & ~n52231;
  assign n52327 = ~n52214 & ~n52232;
  assign n52477 = n52326 & n52327;
  assign n52478 = n52415 ^ n49699;
  assign n52479 = n52478 ^ n52410;
  assign n52480 = n52477 & ~n52479;
  assign n52481 = n52420 ^ n49637;
  assign n52482 = n52481 ^ n52418;
  assign n52483 = n52480 & n52482;
  assign n52484 = ~n52476 & n52483;
  assign n52485 = ~n52474 & ~n52484;
  assign n52486 = ~n52472 & n52485;
  assign n52487 = ~n52471 & ~n52486;
  assign n52433 = n52432 ^ n52401;
  assign n52434 = n52402 & n52433;
  assign n52435 = n52434 ^ n49630;
  assign n52383 = n52382 ^ n52343;
  assign n52384 = n52344 & ~n52383;
  assign n52385 = n52384 ^ n52342;
  assign n52338 = n50804 ^ n50380;
  assign n52339 = n52338 ^ n51776;
  assign n52398 = n52385 ^ n52339;
  assign n51684 = n51683 ^ n51664;
  assign n52399 = n52398 ^ n51684;
  assign n52400 = n52399 ^ n49674;
  assign n52488 = n52435 ^ n52400;
  assign n52489 = ~n52487 & ~n52488;
  assign n52340 = n52339 ^ n51684;
  assign n52386 = n52385 ^ n51684;
  assign n52387 = n52340 & ~n52386;
  assign n52388 = n52387 ^ n52339;
  assign n52336 = n52017 ^ n52014;
  assign n52334 = n50798 ^ n50394;
  assign n52335 = n52334 ^ n51783;
  assign n52337 = n52336 ^ n52335;
  assign n52439 = n52388 ^ n52337;
  assign n52436 = n52435 ^ n52399;
  assign n52437 = n52400 & ~n52436;
  assign n52438 = n52437 ^ n49674;
  assign n52440 = n52439 ^ n52438;
  assign n52490 = n52440 ^ n49751;
  assign n52491 = ~n52489 & ~n52490;
  assign n52441 = n52439 ^ n49751;
  assign n52442 = ~n52440 & ~n52441;
  assign n52443 = n52442 ^ n49751;
  assign n52492 = n52443 ^ n49823;
  assign n52394 = n52020 ^ n52012;
  assign n52392 = n50979 ^ n50612;
  assign n52393 = n52392 ^ n51708;
  assign n52395 = n52394 ^ n52393;
  assign n52389 = n52388 ^ n52336;
  assign n52390 = n52337 & n52389;
  assign n52391 = n52390 ^ n52335;
  assign n52396 = n52395 ^ n52391;
  assign n52493 = n52492 ^ n52396;
  assign n52494 = n52491 & n52493;
  assign n52452 = n52023 ^ n52007;
  assign n52449 = n52393 ^ n52391;
  assign n52450 = ~n52395 & n52449;
  assign n52451 = n52450 ^ n52394;
  assign n52453 = n52452 ^ n52451;
  assign n52447 = n50986 ^ n50634;
  assign n52448 = n52447 ^ n51793;
  assign n52454 = n52453 ^ n52448;
  assign n52397 = n52396 ^ n49823;
  assign n52444 = n52443 ^ n52396;
  assign n52445 = ~n52397 & n52444;
  assign n52446 = n52445 ^ n49823;
  assign n52455 = n52454 ^ n52446;
  assign n52470 = n52455 ^ n49973;
  assign n52679 = n52494 ^ n52470;
  assign n52604 = n50427 ^ n43081;
  assign n52605 = n52604 ^ n46979;
  assign n52606 = n52605 ^ n41408;
  assign n52603 = n52493 ^ n52491;
  assign n52607 = n52606 ^ n52603;
  assign n52609 = n50565 ^ n43086;
  assign n52610 = n52609 ^ n46984;
  assign n52611 = n52610 ^ n41414;
  assign n52608 = n52490 ^ n52489;
  assign n52612 = n52611 ^ n52608;
  assign n52614 = n50432 ^ n42833;
  assign n52615 = n52614 ^ n47114;
  assign n52616 = n52615 ^ n41541;
  assign n52613 = n52488 ^ n52487;
  assign n52617 = n52616 ^ n52613;
  assign n52621 = n52486 ^ n52471;
  assign n52618 = n50437 ^ n42700;
  assign n52619 = n52618 ^ n46989;
  assign n52620 = n52619 ^ n41418;
  assign n52622 = n52621 ^ n52620;
  assign n52624 = n50442 ^ n42705;
  assign n52625 = n52624 ^ n46994;
  assign n52626 = n52625 ^ n41530;
  assign n52623 = n52485 ^ n52472;
  assign n52627 = n52626 ^ n52623;
  assign n52629 = n50447 ^ n2263;
  assign n52630 = n52629 ^ n46999;
  assign n52631 = n52630 ^ n41424;
  assign n52628 = n52484 ^ n52474;
  assign n52632 = n52631 ^ n52628;
  assign n52634 = n50452 ^ n2245;
  assign n52635 = n52634 ^ n47004;
  assign n52636 = n52635 ^ n41519;
  assign n52633 = n52483 ^ n52476;
  assign n52637 = n52636 ^ n52633;
  assign n52650 = n50542 ^ n42714;
  assign n52651 = n52650 ^ n47094;
  assign n52652 = n52651 ^ n41511;
  assign n52639 = n50457 ^ n42719;
  assign n52640 = n52639 ^ n47086;
  assign n52641 = n52640 ^ n41429;
  assign n52638 = n52479 ^ n52477;
  assign n52642 = n52641 ^ n52638;
  assign n52328 = n52327 ^ n52326;
  assign n52309 = n50531 ^ n42793;
  assign n52310 = n52309 ^ n47008;
  assign n52311 = n52310 ^ n41433;
  assign n52643 = n52328 ^ n52311;
  assign n52234 = n50462 ^ n42723;
  assign n52235 = n52234 ^ n47013;
  assign n52236 = n52235 ^ n1745;
  assign n52233 = n52232 ^ n52214;
  assign n52237 = n52236 ^ n52233;
  assign n52239 = n50518 ^ n42782;
  assign n52240 = n52239 ^ n47018;
  assign n52241 = n52240 ^ n41438;
  assign n52238 = n52231 ^ n52230;
  assign n52242 = n52241 ^ n52238;
  assign n52244 = n50467 ^ n42728;
  assign n52245 = n52244 ^ n47024;
  assign n52246 = n52245 ^ n41443;
  assign n52243 = n52229 ^ n52228;
  assign n52247 = n52246 ^ n52243;
  assign n52249 = n50507 ^ n42771;
  assign n52250 = n52249 ^ n47029;
  assign n52251 = n52250 ^ n41449;
  assign n52248 = n52227 ^ n52225;
  assign n52252 = n52251 ^ n52248;
  assign n52289 = n52224 ^ n52223;
  assign n52254 = n50472 ^ n42739;
  assign n52255 = n52254 ^ n47055;
  assign n52256 = n52255 ^ n41459;
  assign n52253 = n52222 ^ n52220;
  assign n52257 = n52256 ^ n52253;
  assign n52259 = n50477 ^ n42743;
  assign n52260 = n52259 ^ n47047;
  assign n52261 = n52260 ^ n41463;
  assign n52258 = n52219 ^ n52218;
  assign n52262 = n52261 ^ n52258;
  assign n52275 = n50481 ^ n42753;
  assign n52276 = n52275 ^ n47033;
  assign n52277 = n52276 ^ n41472;
  assign n52268 = n50484 ^ n42749;
  assign n52269 = n52268 ^ n47036;
  assign n52270 = n52269 ^ n41468;
  assign n52263 = n52157 ^ n48765;
  assign n52264 = n50864 ^ n43204;
  assign n52265 = n52264 ^ n47342;
  assign n52266 = n52265 ^ n41810;
  assign n52267 = ~n52263 & n52266;
  assign n52271 = n52270 ^ n52267;
  assign n52272 = n52267 ^ n52215;
  assign n52273 = n52271 & n52272;
  assign n52274 = n52273 ^ n52270;
  assign n52278 = n52277 ^ n52274;
  assign n52279 = n52217 ^ n52215;
  assign n52280 = n52279 ^ n52274;
  assign n52281 = n52278 & ~n52280;
  assign n52282 = n52281 ^ n52277;
  assign n52283 = n52282 ^ n52258;
  assign n52284 = n52262 & ~n52283;
  assign n52285 = n52284 ^ n52261;
  assign n52286 = n52285 ^ n52253;
  assign n52287 = ~n52257 & n52286;
  assign n52288 = n52287 ^ n52256;
  assign n52290 = n52289 ^ n52288;
  assign n52291 = n50499 ^ n42734;
  assign n52292 = n52291 ^ n47063;
  assign n52293 = n52292 ^ n41454;
  assign n52294 = n52293 ^ n52289;
  assign n52295 = ~n52290 & n52294;
  assign n52296 = n52295 ^ n52293;
  assign n52297 = n52296 ^ n52248;
  assign n52298 = ~n52252 & n52297;
  assign n52299 = n52298 ^ n52251;
  assign n52300 = n52299 ^ n52243;
  assign n52301 = n52247 & ~n52300;
  assign n52302 = n52301 ^ n52246;
  assign n52303 = n52302 ^ n52238;
  assign n52304 = n52242 & ~n52303;
  assign n52305 = n52304 ^ n52241;
  assign n52306 = n52305 ^ n52233;
  assign n52307 = n52237 & ~n52306;
  assign n52308 = n52307 ^ n52236;
  assign n52644 = n52328 ^ n52308;
  assign n52645 = n52643 & ~n52644;
  assign n52646 = n52645 ^ n52311;
  assign n52647 = n52646 ^ n52638;
  assign n52648 = ~n52642 & n52647;
  assign n52649 = n52648 ^ n52641;
  assign n52653 = n52652 ^ n52649;
  assign n52654 = n52482 ^ n52480;
  assign n52655 = n52654 ^ n52649;
  assign n52656 = n52653 & ~n52655;
  assign n52657 = n52656 ^ n52652;
  assign n52658 = n52657 ^ n52633;
  assign n52659 = ~n52637 & n52658;
  assign n52660 = n52659 ^ n52636;
  assign n52661 = n52660 ^ n52628;
  assign n52662 = ~n52632 & n52661;
  assign n52663 = n52662 ^ n52631;
  assign n52664 = n52663 ^ n52623;
  assign n52665 = n52627 & ~n52664;
  assign n52666 = n52665 ^ n52626;
  assign n52667 = n52666 ^ n52621;
  assign n52668 = n52622 & ~n52667;
  assign n52669 = n52668 ^ n52620;
  assign n52670 = n52669 ^ n52613;
  assign n52671 = ~n52617 & n52670;
  assign n52672 = n52671 ^ n52616;
  assign n52673 = n52672 ^ n52608;
  assign n52674 = n52612 & ~n52673;
  assign n52675 = n52674 ^ n52611;
  assign n52676 = n52675 ^ n52603;
  assign n52677 = n52607 & ~n52676;
  assign n52678 = n52677 ^ n52606;
  assign n52680 = n52679 ^ n52678;
  assign n52681 = n50576 ^ n43075;
  assign n52682 = n52681 ^ n46974;
  assign n52683 = n52682 ^ n41555;
  assign n52684 = n52683 ^ n52679;
  assign n52685 = n52680 & ~n52684;
  assign n52686 = n52685 ^ n52683;
  assign n52599 = n50422 ^ n43070;
  assign n52600 = n52599 ^ n46969;
  assign n52601 = n52600 ^ n41404;
  assign n52495 = ~n52470 & n52494;
  assign n52464 = n52031 ^ n52029;
  assign n52465 = n52464 ^ n52026;
  assign n52462 = n50993 ^ n50671;
  assign n52463 = n52462 ^ n51704;
  assign n52466 = n52465 ^ n52463;
  assign n52459 = n52452 ^ n52448;
  assign n52460 = n52453 & n52459;
  assign n52461 = n52460 ^ n52448;
  assign n52467 = n52466 ^ n52461;
  assign n52468 = n52467 ^ n50003;
  assign n52456 = n52454 ^ n49973;
  assign n52457 = ~n52455 & n52456;
  assign n52458 = n52457 ^ n49973;
  assign n52469 = n52468 ^ n52458;
  assign n52598 = n52495 ^ n52469;
  assign n52602 = n52601 ^ n52598;
  assign n52929 = n52686 ^ n52602;
  assign n52932 = n52931 ^ n52929;
  assign n53076 = n52683 ^ n52680;
  assign n52935 = n52675 ^ n52607;
  assign n52933 = n52090 ^ n51445;
  assign n52774 = n52060 ^ n51972;
  assign n52934 = n52933 ^ n52774;
  assign n52936 = n52935 ^ n52934;
  assign n52939 = n52672 ^ n52612;
  assign n52728 = n52057 ^ n51977;
  assign n52937 = n52728 ^ n51401;
  assign n52938 = n52937 ^ n51899;
  assign n52940 = n52939 ^ n52938;
  assign n52577 = n52054 ^ n51982;
  assign n52942 = n52577 ^ n51128;
  assign n52943 = n52942 ^ n51809;
  assign n52941 = n52669 ^ n52617;
  assign n52944 = n52943 ^ n52941;
  assign n52562 = n52051 ^ n51987;
  assign n52947 = n52562 ^ n51696;
  assign n52948 = n52947 ^ n50993;
  assign n52945 = n52666 ^ n52620;
  assign n52946 = n52945 ^ n52621;
  assign n52949 = n52948 ^ n52946;
  assign n52952 = n52663 ^ n52627;
  assign n52950 = n51700 ^ n50986;
  assign n52548 = n52048 ^ n51992;
  assign n52951 = n52950 ^ n52548;
  assign n52953 = n52952 ^ n52951;
  assign n52534 = n52045 ^ n52042;
  assign n52956 = n52534 ^ n50979;
  assign n52957 = n52956 ^ n51704;
  assign n52954 = n52660 ^ n52631;
  assign n52955 = n52954 ^ n52628;
  assign n52958 = n52957 ^ n52955;
  assign n52960 = n51793 ^ n50798;
  assign n52520 = n52037 ^ n51997;
  assign n52961 = n52960 ^ n52520;
  assign n52959 = n52657 ^ n52637;
  assign n52962 = n52961 ^ n52959;
  assign n52966 = n52465 ^ n51783;
  assign n52967 = n52966 ^ n50966;
  assign n52965 = n52646 ^ n52642;
  assign n52968 = n52967 ^ n52965;
  assign n52969 = n51776 ^ n50808;
  assign n52970 = n52969 ^ n52452;
  assign n52312 = n52311 ^ n52308;
  assign n52329 = n52328 ^ n52312;
  assign n52971 = n52970 ^ n52329;
  assign n52972 = n52336 ^ n51766;
  assign n52973 = n52972 ^ n50953;
  assign n52899 = n52302 ^ n52242;
  assign n52974 = n52973 ^ n52899;
  assign n52975 = n51752 ^ n50942;
  assign n52976 = n52975 ^ n52343;
  assign n52911 = n52296 ^ n52251;
  assign n52912 = n52911 ^ n52248;
  assign n52977 = n52976 ^ n52912;
  assign n52978 = n51685 ^ n50822;
  assign n52979 = n52978 ^ n52347;
  assign n52917 = n52293 ^ n52290;
  assign n52980 = n52979 ^ n52917;
  assign n52983 = n51720 ^ n50824;
  assign n52984 = n52983 ^ n52349;
  assign n52981 = n52285 ^ n52256;
  assign n52982 = n52981 ^ n52253;
  assign n52985 = n52984 ^ n52982;
  assign n53011 = n52282 ^ n52261;
  assign n53012 = n53011 ^ n52258;
  assign n52988 = n52279 ^ n52278;
  assign n52986 = n51723 ^ n50828;
  assign n52987 = n52986 ^ n52357;
  assign n52989 = n52988 ^ n52987;
  assign n52992 = n52270 ^ n52215;
  assign n52993 = n52992 ^ n52267;
  assign n52990 = n51730 ^ n50777;
  assign n52991 = n52990 ^ n52361;
  assign n52994 = n52993 ^ n52991;
  assign n52996 = n51674 ^ n50913;
  assign n52997 = n52996 ^ n52317;
  assign n52995 = n52266 ^ n52263;
  assign n52998 = n52997 ^ n52995;
  assign n52496 = n52469 & ~n52495;
  assign n52505 = n52034 ^ n52002;
  assign n52503 = n51128 ^ n50713;
  assign n52504 = n52503 ^ n51700;
  assign n52506 = n52505 ^ n52504;
  assign n52500 = n52465 ^ n52461;
  assign n52501 = ~n52466 & n52500;
  assign n52502 = n52501 ^ n52463;
  assign n52507 = n52506 ^ n52502;
  assign n52497 = n52467 ^ n52458;
  assign n52498 = n52468 & ~n52497;
  assign n52499 = n52498 ^ n50003;
  assign n52508 = n52507 ^ n52499;
  assign n52509 = n52508 ^ n50025;
  assign n52510 = n52496 & n52509;
  assign n52518 = n51401 ^ n50750;
  assign n52519 = n52518 ^ n51696;
  assign n52521 = n52520 ^ n52519;
  assign n52515 = n52504 ^ n52502;
  assign n52516 = n52506 & n52515;
  assign n52517 = n52516 ^ n52505;
  assign n52522 = n52521 ^ n52517;
  assign n52511 = n52507 ^ n50025;
  assign n52512 = n52508 & n52511;
  assign n52513 = n52512 ^ n50025;
  assign n52514 = n52513 ^ n50056;
  assign n52523 = n52522 ^ n52514;
  assign n52524 = ~n52510 & ~n52523;
  assign n52532 = n51445 ^ n50857;
  assign n52533 = n52532 ^ n51809;
  assign n52535 = n52534 ^ n52533;
  assign n52529 = n52520 ^ n52517;
  assign n52530 = n52521 & n52529;
  assign n52531 = n52530 ^ n52519;
  assign n52536 = n52535 ^ n52531;
  assign n52537 = n52536 ^ n50083;
  assign n52525 = n52522 ^ n50056;
  assign n52526 = n52522 ^ n52513;
  assign n52527 = ~n52525 & n52526;
  assign n52528 = n52527 ^ n50056;
  assign n52538 = n52537 ^ n52528;
  assign n52539 = n52524 & ~n52538;
  assign n52546 = n50642 ^ n49982;
  assign n52547 = n52546 ^ n51899;
  assign n52549 = n52548 ^ n52547;
  assign n52543 = n52534 ^ n52531;
  assign n52544 = ~n52535 & ~n52543;
  assign n52545 = n52544 ^ n52533;
  assign n52550 = n52549 ^ n52545;
  assign n52551 = n52550 ^ n49367;
  assign n52540 = n52536 ^ n52528;
  assign n52541 = ~n52537 & n52540;
  assign n52542 = n52541 ^ n50083;
  assign n52552 = n52551 ^ n52542;
  assign n52553 = ~n52539 & n52552;
  assign n52559 = n52548 ^ n52545;
  assign n52560 = n52549 & ~n52559;
  assign n52561 = n52560 ^ n52547;
  assign n52563 = n52562 ^ n52561;
  assign n52557 = n50681 ^ n50010;
  assign n52558 = n52557 ^ n52090;
  assign n52564 = n52563 ^ n52558;
  assign n52565 = n52564 ^ n49372;
  assign n52554 = n52550 ^ n52542;
  assign n52555 = ~n52551 & n52554;
  assign n52556 = n52555 ^ n49367;
  assign n52566 = n52565 ^ n52556;
  assign n52567 = ~n52553 & n52566;
  assign n52574 = n50724 ^ n50036;
  assign n52575 = n52574 ^ n51419;
  assign n52571 = n52562 ^ n52558;
  assign n52572 = ~n52563 & n52571;
  assign n52573 = n52572 ^ n52558;
  assign n52576 = n52575 ^ n52573;
  assign n52578 = n52577 ^ n52576;
  assign n52579 = n52578 ^ n49379;
  assign n52568 = n52564 ^ n52556;
  assign n52569 = n52565 & n52568;
  assign n52570 = n52569 ^ n49372;
  assign n52580 = n52579 ^ n52570;
  assign n52718 = ~n52567 & ~n52580;
  assign n52726 = n50763 ^ n50070;
  assign n52727 = n52726 ^ n51422;
  assign n52729 = n52728 ^ n52727;
  assign n52722 = n52577 ^ n52575;
  assign n52723 = n52577 ^ n52573;
  assign n52724 = ~n52722 & n52723;
  assign n52725 = n52724 ^ n52575;
  assign n52730 = n52729 ^ n52725;
  assign n52731 = n52730 ^ n49362;
  assign n52719 = n52578 ^ n52570;
  assign n52720 = ~n52579 & n52719;
  assign n52721 = n52720 ^ n49379;
  assign n52732 = n52731 ^ n52721;
  assign n52765 = ~n52718 & ~n52732;
  assign n52772 = n50866 ^ n50095;
  assign n52773 = n52772 ^ n51426;
  assign n52775 = n52774 ^ n52773;
  assign n52769 = n52727 ^ n52725;
  assign n52770 = n52729 & n52769;
  assign n52771 = n52770 ^ n52728;
  assign n52776 = n52775 ^ n52771;
  assign n52766 = n52730 ^ n52721;
  assign n52767 = n52731 & ~n52766;
  assign n52768 = n52767 ^ n49362;
  assign n52777 = n52776 ^ n52768;
  assign n52778 = n52777 ^ n49358;
  assign n52792 = n52765 & n52778;
  assign n52800 = n52774 ^ n52771;
  assign n52801 = ~n52775 & ~n52800;
  assign n52802 = n52801 ^ n52773;
  assign n52798 = n52068 ^ n52065;
  assign n52796 = n50837 ^ n49664;
  assign n52797 = n52796 ^ n51411;
  assign n52799 = n52798 ^ n52797;
  assign n52803 = n52802 ^ n52799;
  assign n52793 = n52776 ^ n49358;
  assign n52794 = ~n52777 & ~n52793;
  assign n52795 = n52794 ^ n49358;
  assign n52804 = n52803 ^ n52795;
  assign n52805 = n52804 ^ n48772;
  assign n52881 = ~n52792 & ~n52805;
  assign n52877 = n50743 ^ n43160;
  assign n52878 = n52877 ^ n47289;
  assign n52879 = n52878 ^ n2405;
  assign n52871 = n50833 ^ n49660;
  assign n52872 = n52871 ^ n51457;
  assign n52874 = n52873 ^ n52872;
  assign n52868 = n52802 ^ n52797;
  assign n52869 = ~n52799 & n52868;
  assign n52870 = n52869 ^ n52802;
  assign n52875 = n52874 ^ n52870;
  assign n52864 = n52803 ^ n48772;
  assign n52865 = n52804 & n52864;
  assign n52866 = n52865 ^ n48772;
  assign n52867 = n52866 ^ n48771;
  assign n52876 = n52875 ^ n52867;
  assign n52880 = n52879 ^ n52876;
  assign n52882 = n52881 ^ n52880;
  assign n52807 = n50722 ^ n43044;
  assign n52808 = n52807 ^ n47322;
  assign n52809 = n52808 ^ n41779;
  assign n52806 = n52805 ^ n52792;
  assign n52810 = n52809 ^ n52806;
  assign n52779 = n52778 ^ n52765;
  assign n52761 = n50679 ^ n43048;
  assign n52762 = n52761 ^ n47169;
  assign n52763 = n52762 ^ n41784;
  assign n52788 = n52779 ^ n52763;
  assign n52733 = n52732 ^ n52718;
  assign n1254 = n1253 ^ n1199;
  assign n1291 = n1290 ^ n1254;
  assign n1301 = n1300 ^ n1291;
  assign n52734 = n52733 ^ n1301;
  assign n52581 = n52580 ^ n52567;
  assign n52331 = n50621 ^ n43053;
  assign n52332 = n52331 ^ n46939;
  assign n52333 = n52332 ^ n1282;
  assign n52582 = n52581 ^ n52333;
  assign n52707 = n50402 ^ n1098;
  assign n52708 = n52707 ^ n46944;
  assign n52709 = n52708 ^ n41595;
  assign n52584 = n50407 ^ n43121;
  assign n52585 = n52584 ^ n46949;
  assign n52586 = n52585 ^ n41384;
  assign n52583 = n52552 ^ n52539;
  assign n52587 = n52586 ^ n52583;
  assign n52589 = n50412 ^ n43061;
  assign n52590 = n52589 ^ n46954;
  assign n52591 = n52590 ^ n41388;
  assign n52588 = n52538 ^ n52524;
  assign n52592 = n52591 ^ n52588;
  assign n52693 = n52523 ^ n52510;
  assign n52594 = n50417 ^ n43066;
  assign n52595 = n52594 ^ n46964;
  assign n52596 = n52595 ^ n41398;
  assign n52593 = n52509 ^ n52496;
  assign n52597 = n52596 ^ n52593;
  assign n52687 = n52686 ^ n52598;
  assign n52688 = n52602 & ~n52687;
  assign n52689 = n52688 ^ n52601;
  assign n52690 = n52689 ^ n52593;
  assign n52691 = ~n52597 & n52690;
  assign n52692 = n52691 ^ n52596;
  assign n52694 = n52693 ^ n52692;
  assign n52695 = n50590 ^ n43110;
  assign n52696 = n52695 ^ n46959;
  assign n52697 = n52696 ^ n41394;
  assign n52698 = n52697 ^ n52693;
  assign n52699 = ~n52694 & n52698;
  assign n52700 = n52699 ^ n52697;
  assign n52701 = n52700 ^ n52588;
  assign n52702 = ~n52592 & n52701;
  assign n52703 = n52702 ^ n52591;
  assign n52704 = n52703 ^ n52583;
  assign n52705 = n52587 & ~n52704;
  assign n52706 = n52705 ^ n52586;
  assign n52710 = n52709 ^ n52706;
  assign n52711 = n52566 ^ n52553;
  assign n52712 = n52711 ^ n52706;
  assign n52713 = n52710 & n52712;
  assign n52714 = n52713 ^ n52709;
  assign n52715 = n52714 ^ n52581;
  assign n52716 = ~n52582 & n52715;
  assign n52717 = n52716 ^ n52333;
  assign n52758 = n52733 ^ n52717;
  assign n52759 = n52734 & ~n52758;
  assign n52760 = n52759 ^ n1301;
  assign n52789 = n52779 ^ n52760;
  assign n52790 = n52788 & ~n52789;
  assign n52791 = n52790 ^ n52763;
  assign n52861 = n52806 ^ n52791;
  assign n52862 = ~n52810 & n52861;
  assign n52863 = n52862 ^ n52809;
  assign n52883 = n52882 ^ n52863;
  assign n52764 = n52763 ^ n52760;
  assign n52780 = n52779 ^ n52764;
  assign n52755 = n51481 ^ n50894;
  assign n52756 = n52755 ^ n52184;
  assign n52815 = n52780 ^ n52756;
  assign n52738 = n51471 ^ n50879;
  assign n52739 = n52738 ^ n52139;
  assign n52740 = n52714 ^ n52333;
  assign n52741 = n52740 ^ n52581;
  assign n52742 = n52739 & ~n52741;
  assign n52736 = n50887 ^ n50774;
  assign n52737 = n52736 ^ n52147;
  assign n52743 = n52742 ^ n52737;
  assign n52735 = n52734 ^ n52717;
  assign n52752 = n52737 ^ n52735;
  assign n52753 = ~n52743 & n52752;
  assign n52754 = n52753 ^ n52742;
  assign n52816 = n52780 ^ n52754;
  assign n52817 = ~n52815 & ~n52816;
  assign n52818 = n52817 ^ n52756;
  assign n52812 = n51488 ^ n50788;
  assign n52813 = n52812 ^ n52196;
  assign n52857 = n52818 ^ n52813;
  assign n52811 = n52810 ^ n52791;
  assign n52858 = n52818 ^ n52811;
  assign n52859 = ~n52857 & ~n52858;
  assign n52860 = n52859 ^ n52813;
  assign n52884 = n52883 ^ n52860;
  assign n52855 = n51549 ^ n50781;
  assign n52856 = n52855 ^ n52211;
  assign n52999 = n52883 ^ n52856;
  assign n53000 = n52884 & n52999;
  assign n53001 = n53000 ^ n52856;
  assign n53002 = n53001 ^ n52995;
  assign n53003 = n52998 & ~n53002;
  assign n53004 = n53003 ^ n52997;
  assign n53005 = n53004 ^ n52993;
  assign n53006 = n52994 & ~n53005;
  assign n53007 = n53006 ^ n52991;
  assign n53008 = n53007 ^ n52987;
  assign n53009 = ~n52989 & ~n53008;
  assign n53010 = n53009 ^ n52988;
  assign n53013 = n53012 ^ n53010;
  assign n53014 = n51722 ^ n50929;
  assign n53015 = n53014 ^ n52353;
  assign n53016 = n53015 ^ n53012;
  assign n53017 = ~n53013 & n53016;
  assign n53018 = n53017 ^ n53015;
  assign n53019 = n53018 ^ n52982;
  assign n53020 = ~n52985 & n53019;
  assign n53021 = n53020 ^ n52984;
  assign n53022 = n53021 ^ n52917;
  assign n53023 = n52980 & ~n53022;
  assign n53024 = n53023 ^ n52979;
  assign n53025 = n53024 ^ n52976;
  assign n53026 = ~n52977 & ~n53025;
  assign n53027 = n53026 ^ n52912;
  assign n52906 = n52299 ^ n52247;
  assign n53028 = n53027 ^ n52906;
  assign n53029 = n51759 ^ n50818;
  assign n53030 = n53029 ^ n51684;
  assign n53031 = n53030 ^ n52906;
  assign n53032 = n53028 & n53031;
  assign n53033 = n53032 ^ n53030;
  assign n53034 = n53033 ^ n52899;
  assign n53035 = ~n52974 & ~n53034;
  assign n53036 = n53035 ^ n52973;
  assign n52894 = n52305 ^ n52237;
  assign n53037 = n53036 ^ n52894;
  assign n53038 = n52394 ^ n51713;
  assign n53039 = n53038 ^ n50813;
  assign n53040 = n53039 ^ n52894;
  assign n53041 = n53037 & ~n53040;
  assign n53042 = n53041 ^ n53039;
  assign n53043 = n53042 ^ n52329;
  assign n53044 = n52971 & n53043;
  assign n53045 = n53044 ^ n52970;
  assign n53046 = n53045 ^ n52967;
  assign n53047 = n52968 & n53046;
  assign n53048 = n53047 ^ n52965;
  assign n52963 = n52654 ^ n52652;
  assign n52964 = n52963 ^ n52649;
  assign n53049 = n53048 ^ n52964;
  assign n53050 = n52505 ^ n50804;
  assign n53051 = n53050 ^ n51708;
  assign n53052 = n53051 ^ n52964;
  assign n53053 = n53049 & n53052;
  assign n53054 = n53053 ^ n53051;
  assign n53055 = n53054 ^ n52959;
  assign n53056 = ~n52962 & n53055;
  assign n53057 = n53056 ^ n52961;
  assign n53058 = n53057 ^ n52955;
  assign n53059 = n52958 & n53058;
  assign n53060 = n53059 ^ n52957;
  assign n53061 = n53060 ^ n52951;
  assign n53062 = ~n52953 & ~n53061;
  assign n53063 = n53062 ^ n52952;
  assign n53064 = n53063 ^ n52946;
  assign n53065 = n52949 & ~n53064;
  assign n53066 = n53065 ^ n52948;
  assign n53067 = n53066 ^ n52941;
  assign n53068 = n52944 & n53067;
  assign n53069 = n53068 ^ n52943;
  assign n53070 = n53069 ^ n52939;
  assign n53071 = ~n52940 & n53070;
  assign n53072 = n53071 ^ n52938;
  assign n53073 = n53072 ^ n52934;
  assign n53074 = n52936 & n53073;
  assign n53075 = n53074 ^ n52935;
  assign n53077 = n53076 ^ n53075;
  assign n53078 = n51419 ^ n50642;
  assign n53079 = n53078 ^ n52798;
  assign n53080 = n53079 ^ n53076;
  assign n53081 = n53077 & ~n53080;
  assign n53082 = n53081 ^ n53079;
  assign n53083 = n53082 ^ n52929;
  assign n53084 = ~n52932 & ~n53083;
  assign n53085 = n53084 ^ n52931;
  assign n52926 = n52117 ^ n50724;
  assign n52927 = n52926 ^ n51426;
  assign n53219 = n53085 ^ n52927;
  assign n52925 = n52689 ^ n52597;
  assign n53220 = n53219 ^ n52925;
  assign n53291 = n53220 ^ n50036;
  assign n53100 = n53082 ^ n52932;
  assign n53101 = n53100 ^ n50010;
  assign n53102 = n53079 ^ n53077;
  assign n53103 = n53102 ^ n49982;
  assign n53104 = n53072 ^ n52936;
  assign n53105 = n53104 ^ n50857;
  assign n53106 = n53069 ^ n52938;
  assign n53107 = n53106 ^ n52939;
  assign n53108 = n53107 ^ n50750;
  assign n53109 = n53066 ^ n52944;
  assign n53110 = n53109 ^ n50713;
  assign n53111 = n53063 ^ n52948;
  assign n53112 = n53111 ^ n52946;
  assign n53113 = n53112 ^ n50671;
  assign n53114 = n53060 ^ n52953;
  assign n53115 = n53114 ^ n50634;
  assign n53116 = n53057 ^ n52958;
  assign n53117 = n53116 ^ n50612;
  assign n53118 = n53054 ^ n52961;
  assign n53119 = n53118 ^ n52959;
  assign n53120 = n53119 ^ n50394;
  assign n53186 = n53051 ^ n53049;
  assign n53121 = n53045 ^ n52968;
  assign n53122 = n53121 ^ n50366;
  assign n53123 = n53042 ^ n52971;
  assign n53124 = n53123 ^ n50350;
  assign n53125 = n53039 ^ n53037;
  assign n53126 = n53125 ^ n50336;
  assign n53127 = n53033 ^ n52973;
  assign n53128 = n53127 ^ n52899;
  assign n53129 = n53128 ^ n50323;
  assign n53130 = n53030 ^ n53028;
  assign n53131 = n53130 ^ n50266;
  assign n53132 = n53024 ^ n52977;
  assign n53133 = n53132 ^ n49629;
  assign n53162 = n53021 ^ n52979;
  assign n53163 = n53162 ^ n52917;
  assign n53134 = n53018 ^ n52985;
  assign n53135 = n53134 ^ n49633;
  assign n53136 = n53015 ^ n53013;
  assign n53137 = n53136 ^ n49634;
  assign n53138 = n53004 ^ n52994;
  assign n53139 = n53138 ^ n49641;
  assign n52814 = n52813 ^ n52811;
  assign n52819 = n52818 ^ n52814;
  assign n52757 = n52756 ^ n52754;
  assign n52781 = n52780 ^ n52757;
  assign n52782 = n52781 ^ n50118;
  assign n52745 = n52741 ^ n52739;
  assign n52746 = n50108 & ~n52745;
  assign n52747 = n52746 ^ n49653;
  assign n52744 = n52743 ^ n52735;
  assign n52749 = n52746 ^ n52744;
  assign n52750 = ~n52747 & n52749;
  assign n52751 = n52750 ^ n49653;
  assign n52785 = n52781 ^ n52751;
  assign n52786 = ~n52782 & ~n52785;
  assign n52787 = n52786 ^ n50118;
  assign n52820 = n52819 ^ n52787;
  assign n52886 = n52819 ^ n49648;
  assign n52887 = ~n52820 & ~n52886;
  assign n52888 = n52887 ^ n49648;
  assign n52889 = n52888 ^ n50128;
  assign n52885 = n52884 ^ n52856;
  assign n53140 = n52888 ^ n52885;
  assign n53141 = n52889 & n53140;
  assign n53142 = n53141 ^ n50128;
  assign n53143 = n53142 ^ n49642;
  assign n53144 = n53001 ^ n52998;
  assign n53145 = n53144 ^ n53142;
  assign n53146 = ~n53143 & ~n53145;
  assign n53147 = n53146 ^ n49642;
  assign n53148 = n53147 ^ n53138;
  assign n53149 = ~n53139 & n53148;
  assign n53150 = n53149 ^ n49641;
  assign n53151 = n53150 ^ n49635;
  assign n53152 = n53007 ^ n52989;
  assign n53153 = n53152 ^ n53150;
  assign n53154 = n53151 & ~n53153;
  assign n53155 = n53154 ^ n49635;
  assign n53156 = n53155 ^ n53136;
  assign n53157 = ~n53137 & ~n53156;
  assign n53158 = n53157 ^ n49634;
  assign n53159 = n53158 ^ n53134;
  assign n53160 = n53135 & ~n53159;
  assign n53161 = n53160 ^ n49633;
  assign n53164 = n53163 ^ n53161;
  assign n53165 = n53163 ^ n50160;
  assign n53166 = n53164 & ~n53165;
  assign n53167 = n53166 ^ n50160;
  assign n53168 = n53167 ^ n53132;
  assign n53169 = ~n53133 & ~n53168;
  assign n53170 = n53169 ^ n49629;
  assign n53171 = n53170 ^ n53130;
  assign n53172 = n53131 & n53171;
  assign n53173 = n53172 ^ n50266;
  assign n53174 = n53173 ^ n53128;
  assign n53175 = ~n53129 & ~n53174;
  assign n53176 = n53175 ^ n50323;
  assign n53177 = n53176 ^ n53125;
  assign n53178 = n53126 & ~n53177;
  assign n53179 = n53178 ^ n50336;
  assign n53180 = n53179 ^ n53123;
  assign n53181 = ~n53124 & n53180;
  assign n53182 = n53181 ^ n50350;
  assign n53183 = n53182 ^ n53121;
  assign n53184 = ~n53122 & ~n53183;
  assign n53185 = n53184 ^ n50366;
  assign n53187 = n53186 ^ n53185;
  assign n53188 = n53186 ^ n50380;
  assign n53189 = ~n53187 & ~n53188;
  assign n53190 = n53189 ^ n50380;
  assign n53191 = n53190 ^ n53119;
  assign n53192 = ~n53120 & n53191;
  assign n53193 = n53192 ^ n50394;
  assign n53194 = n53193 ^ n53116;
  assign n53195 = ~n53117 & ~n53194;
  assign n53196 = n53195 ^ n50612;
  assign n53197 = n53196 ^ n53114;
  assign n53198 = ~n53115 & n53197;
  assign n53199 = n53198 ^ n50634;
  assign n53200 = n53199 ^ n53112;
  assign n53201 = ~n53113 & n53200;
  assign n53202 = n53201 ^ n50671;
  assign n53203 = n53202 ^ n53109;
  assign n53204 = n53110 & n53203;
  assign n53205 = n53204 ^ n50713;
  assign n53206 = n53205 ^ n53107;
  assign n53207 = ~n53108 & ~n53206;
  assign n53208 = n53207 ^ n50750;
  assign n53209 = n53208 ^ n53104;
  assign n53210 = n53105 & ~n53209;
  assign n53211 = n53210 ^ n50857;
  assign n53212 = n53211 ^ n53102;
  assign n53213 = n53103 & ~n53212;
  assign n53214 = n53213 ^ n49982;
  assign n53215 = n53214 ^ n53100;
  assign n53216 = ~n53101 & ~n53215;
  assign n53217 = n53216 ^ n50010;
  assign n53292 = n53291 ^ n53217;
  assign n53241 = n53214 ^ n53101;
  assign n53242 = n53211 ^ n53103;
  assign n53243 = n53205 ^ n53108;
  assign n53244 = n53202 ^ n53110;
  assign n53245 = n53199 ^ n53113;
  assign n53246 = n53196 ^ n53115;
  assign n53247 = n53167 ^ n53133;
  assign n53248 = n53164 ^ n50160;
  assign n53249 = n53147 ^ n53139;
  assign n53250 = n53144 ^ n53143;
  assign n52748 = n52747 ^ n52744;
  assign n52783 = n52782 ^ n52751;
  assign n52784 = ~n52748 & ~n52783;
  assign n52821 = n52820 ^ n49648;
  assign n52854 = ~n52784 & ~n52821;
  assign n52890 = n52889 ^ n52885;
  assign n53251 = ~n52854 & ~n52890;
  assign n53252 = n53250 & ~n53251;
  assign n53253 = n53249 & ~n53252;
  assign n53254 = n53152 ^ n53151;
  assign n53255 = n53253 & ~n53254;
  assign n53256 = n53155 ^ n49634;
  assign n53257 = n53256 ^ n53136;
  assign n53258 = n53255 & n53257;
  assign n53259 = n53158 ^ n53135;
  assign n53260 = ~n53258 & ~n53259;
  assign n53261 = n53248 & n53260;
  assign n53262 = n53247 & n53261;
  assign n53263 = n53170 ^ n53131;
  assign n53264 = n53262 & n53263;
  assign n53265 = n53173 ^ n53129;
  assign n53266 = n53264 & n53265;
  assign n53267 = n53176 ^ n50336;
  assign n53268 = n53267 ^ n53125;
  assign n53269 = ~n53266 & ~n53268;
  assign n53270 = n53179 ^ n50350;
  assign n53271 = n53270 ^ n53123;
  assign n53272 = n53269 & n53271;
  assign n53273 = n53182 ^ n50366;
  assign n53274 = n53273 ^ n53121;
  assign n53275 = ~n53272 & ~n53274;
  assign n53276 = n53187 ^ n50380;
  assign n53277 = ~n53275 & ~n53276;
  assign n53278 = n53190 ^ n53120;
  assign n53279 = ~n53277 & ~n53278;
  assign n53280 = n53193 ^ n53117;
  assign n53281 = n53279 & ~n53280;
  assign n53282 = n53246 & n53281;
  assign n53283 = ~n53245 & ~n53282;
  assign n53284 = n53244 & n53283;
  assign n53285 = ~n53243 & ~n53284;
  assign n53286 = n53208 ^ n50857;
  assign n53287 = n53286 ^ n53104;
  assign n53288 = n53285 & ~n53287;
  assign n53289 = n53242 & ~n53288;
  assign n53290 = n53241 & ~n53289;
  assign n53313 = n53292 ^ n53290;
  assign n53317 = n53316 ^ n53313;
  assign n53490 = n51202 ^ n43509;
  assign n53491 = n53490 ^ n47725;
  assign n53492 = n53491 ^ n42449;
  assign n53319 = n51371 ^ n43513;
  assign n53320 = n53319 ^ n47730;
  assign n53321 = n53320 ^ n42437;
  assign n53318 = n53288 ^ n53242;
  assign n53322 = n53321 ^ n53318;
  assign n53326 = n53287 ^ n53285;
  assign n53323 = n51207 ^ n43519;
  assign n53324 = n53323 ^ n47905;
  assign n53325 = n53324 ^ n869;
  assign n53327 = n53326 ^ n53325;
  assign n53329 = n51360 ^ n43694;
  assign n53330 = n53329 ^ n47735;
  assign n53331 = n53330 ^ n42099;
  assign n53328 = n53284 ^ n53243;
  assign n53332 = n53331 ^ n53328;
  assign n53334 = n47740 ^ n43524;
  assign n53335 = n53334 ^ n51212;
  assign n53336 = n53335 ^ n42104;
  assign n53333 = n53283 ^ n53244;
  assign n53337 = n53336 ^ n53333;
  assign n53339 = n51217 ^ n43529;
  assign n53340 = n53339 ^ n47891;
  assign n53341 = n53340 ^ n42109;
  assign n53338 = n53282 ^ n53245;
  assign n53342 = n53341 ^ n53338;
  assign n53344 = n51346 ^ n43533;
  assign n53345 = n53344 ^ n47883;
  assign n53346 = n53345 ^ n42114;
  assign n53343 = n53281 ^ n53246;
  assign n53347 = n53346 ^ n53343;
  assign n53351 = n53280 ^ n53279;
  assign n53348 = n51222 ^ n43539;
  assign n53349 = n53348 ^ n47875;
  assign n53350 = n53349 ^ n42251;
  assign n53352 = n53351 ^ n53350;
  assign n53354 = n51335 ^ n43674;
  assign n53355 = n53354 ^ n47867;
  assign n53356 = n53355 ^ n42118;
  assign n53353 = n53278 ^ n53277;
  assign n53357 = n53356 ^ n53353;
  assign n53359 = n51227 ^ n43666;
  assign n53360 = n53359 ^ n47859;
  assign n53361 = n53360 ^ n42240;
  assign n53358 = n53276 ^ n53275;
  assign n53362 = n53361 ^ n53358;
  assign n53364 = n51232 ^ n43544;
  assign n53365 = n53364 ^ n47745;
  assign n53366 = n53365 ^ n42124;
  assign n53363 = n53274 ^ n53272;
  assign n53367 = n53366 ^ n53363;
  assign n53369 = n51237 ^ n43549;
  assign n53370 = n53369 ^ n47750;
  assign n53371 = n53370 ^ n42229;
  assign n53368 = n53271 ^ n53269;
  assign n53372 = n53371 ^ n53368;
  assign n53449 = n53268 ^ n53266;
  assign n53374 = n51315 ^ n43559;
  assign n53375 = n53374 ^ n47842;
  assign n53376 = n53375 ^ n2111;
  assign n53373 = n53265 ^ n53264;
  assign n53377 = n53376 ^ n53373;
  assign n53381 = n53263 ^ n53262;
  assign n53378 = n51247 ^ n43564;
  assign n53379 = n53378 ^ n1976;
  assign n53380 = n53379 ^ n42133;
  assign n53382 = n53381 ^ n53380;
  assign n53386 = n53261 ^ n53247;
  assign n53383 = n51251 ^ n43643;
  assign n53384 = n53383 ^ n47759;
  assign n53385 = n53384 ^ n1965;
  assign n53387 = n53386 ^ n53385;
  assign n53391 = n53260 ^ n53248;
  assign n53388 = n51301 ^ n1811;
  assign n53389 = n53388 ^ n47765;
  assign n53390 = n53389 ^ n42140;
  assign n53392 = n53391 ^ n53390;
  assign n53394 = n51257 ^ n43568;
  assign n53395 = n53394 ^ n47770;
  assign n53396 = n53395 ^ n42204;
  assign n53393 = n53259 ^ n53258;
  assign n53397 = n53396 ^ n53393;
  assign n53398 = n53257 ^ n53255;
  assign n53402 = n53401 ^ n53398;
  assign n53404 = n51262 ^ n43574;
  assign n53405 = n53404 ^ n47779;
  assign n53406 = n53405 ^ n42151;
  assign n53403 = n53254 ^ n53253;
  assign n53407 = n53406 ^ n53403;
  assign n53411 = n53252 ^ n53249;
  assign n53408 = n51279 ^ n43616;
  assign n53409 = n53408 ^ n47785;
  assign n53410 = n53409 ^ n42156;
  assign n53412 = n53411 ^ n53410;
  assign n53417 = n51267 ^ n43579;
  assign n53418 = n53417 ^ n47811;
  assign n53419 = n53418 ^ n42161;
  assign n52891 = n52890 ^ n52854;
  assign n52850 = n50772 ^ n43584;
  assign n52851 = n52850 ^ n47790;
  assign n52852 = n52851 ^ n42184;
  assign n53413 = n52891 ^ n52852;
  assign n52823 = n50691 ^ n43589;
  assign n52824 = n52823 ^ n47798;
  assign n52825 = n52824 ^ n42165;
  assign n52822 = n52821 ^ n52784;
  assign n52826 = n52825 ^ n52822;
  assign n52828 = n50653 ^ n43598;
  assign n52829 = n52828 ^ n2621;
  assign n52830 = n52829 ^ n42171;
  assign n52827 = n52783 ^ n52748;
  assign n52831 = n52830 ^ n52827;
  assign n52837 = n50649 ^ n43593;
  assign n52838 = n52837 ^ n47206;
  assign n52839 = n52838 ^ n2610;
  assign n52832 = n51448 ^ n2468;
  assign n52833 = n52832 ^ n47942;
  assign n52834 = n52833 ^ n42523;
  assign n52835 = n52745 ^ n50108;
  assign n52836 = n52834 & ~n52835;
  assign n52840 = n52839 ^ n52836;
  assign n52841 = n52836 ^ n52748;
  assign n52842 = n52840 & n52841;
  assign n52843 = n52842 ^ n52839;
  assign n52844 = n52843 ^ n52827;
  assign n52845 = ~n52831 & n52844;
  assign n52846 = n52845 ^ n52830;
  assign n52847 = n52846 ^ n52822;
  assign n52848 = n52826 & ~n52847;
  assign n52849 = n52848 ^ n52825;
  assign n53414 = n52891 ^ n52849;
  assign n53415 = ~n53413 & n53414;
  assign n53416 = n53415 ^ n52852;
  assign n53420 = n53419 ^ n53416;
  assign n53421 = n53251 ^ n53250;
  assign n53422 = n53421 ^ n53416;
  assign n53423 = n53420 & n53422;
  assign n53424 = n53423 ^ n53419;
  assign n53425 = n53424 ^ n53411;
  assign n53426 = n53412 & ~n53425;
  assign n53427 = n53426 ^ n53410;
  assign n53428 = n53427 ^ n53403;
  assign n53429 = n53407 & ~n53428;
  assign n53430 = n53429 ^ n53406;
  assign n53431 = n53430 ^ n53398;
  assign n53432 = ~n53402 & n53431;
  assign n53433 = n53432 ^ n53401;
  assign n53434 = n53433 ^ n53393;
  assign n53435 = n53397 & ~n53434;
  assign n53436 = n53435 ^ n53396;
  assign n53437 = n53436 ^ n53391;
  assign n53438 = n53392 & ~n53437;
  assign n53439 = n53438 ^ n53390;
  assign n53440 = n53439 ^ n53386;
  assign n53441 = n53387 & ~n53440;
  assign n53442 = n53441 ^ n53385;
  assign n53443 = n53442 ^ n53381;
  assign n53444 = n53382 & ~n53443;
  assign n53445 = n53444 ^ n53380;
  assign n53446 = n53445 ^ n53373;
  assign n53447 = n53377 & ~n53446;
  assign n53448 = n53447 ^ n53376;
  assign n53450 = n53449 ^ n53448;
  assign n53451 = n51242 ^ n43554;
  assign n53452 = n53451 ^ n47755;
  assign n53453 = n53452 ^ n42129;
  assign n53454 = n53453 ^ n53449;
  assign n53455 = n53450 & ~n53454;
  assign n53456 = n53455 ^ n53453;
  assign n53457 = n53456 ^ n53368;
  assign n53458 = ~n53372 & n53457;
  assign n53459 = n53458 ^ n53371;
  assign n53460 = n53459 ^ n53363;
  assign n53461 = n53367 & ~n53460;
  assign n53462 = n53461 ^ n53366;
  assign n53463 = n53462 ^ n53358;
  assign n53464 = ~n53362 & n53463;
  assign n53465 = n53464 ^ n53361;
  assign n53466 = n53465 ^ n53353;
  assign n53467 = n53357 & ~n53466;
  assign n53468 = n53467 ^ n53356;
  assign n53469 = n53468 ^ n53350;
  assign n53470 = ~n53352 & ~n53469;
  assign n53471 = n53470 ^ n53351;
  assign n53472 = n53471 ^ n53343;
  assign n53473 = n53347 & n53472;
  assign n53474 = n53473 ^ n53346;
  assign n53475 = n53474 ^ n53338;
  assign n53476 = ~n53342 & n53475;
  assign n53477 = n53476 ^ n53341;
  assign n53478 = n53477 ^ n53333;
  assign n53479 = ~n53337 & n53478;
  assign n53480 = n53479 ^ n53336;
  assign n53481 = n53480 ^ n53328;
  assign n53482 = n53332 & ~n53481;
  assign n53483 = n53482 ^ n53331;
  assign n53484 = n53483 ^ n53325;
  assign n53485 = ~n53327 & ~n53484;
  assign n53486 = n53485 ^ n53326;
  assign n53487 = n53486 ^ n53318;
  assign n53488 = n53322 & n53487;
  assign n53489 = n53488 ^ n53321;
  assign n53493 = n53492 ^ n53489;
  assign n53494 = n53289 ^ n53241;
  assign n53495 = n53494 ^ n53489;
  assign n53496 = n53493 & n53495;
  assign n53497 = n53496 ^ n53492;
  assign n53498 = n53497 ^ n53313;
  assign n53499 = n53317 & ~n53498;
  assign n53500 = n53499 ^ n53316;
  assign n53309 = n51192 ^ n1390;
  assign n53310 = n53309 ^ n47922;
  assign n53311 = n53310 ^ n42460;
  assign n53218 = n53217 ^ n50036;
  assign n53221 = n53220 ^ n53217;
  assign n53222 = n53218 & n53221;
  assign n53223 = n53222 ^ n50036;
  assign n52928 = n52927 ^ n52925;
  assign n53086 = n53085 ^ n52925;
  assign n53087 = n52928 & ~n53086;
  assign n53088 = n53087 ^ n52927;
  assign n52922 = n51411 ^ n50763;
  assign n52923 = n52922 ^ n52122;
  assign n52921 = n52697 ^ n52694;
  assign n52924 = n52923 ^ n52921;
  assign n53098 = n53088 ^ n52924;
  assign n53099 = n53098 ^ n50070;
  assign n53294 = n53223 ^ n53099;
  assign n53293 = ~n53290 & n53292;
  assign n53308 = n53294 ^ n53293;
  assign n53312 = n53311 ^ n53308;
  assign n53549 = n53500 ^ n53312;
  assign n53544 = n53497 ^ n53317;
  assign n53545 = n52184 ^ n51471;
  assign n53546 = n53545 ^ n52995;
  assign n53547 = n53544 & n53546;
  assign n53542 = n52993 ^ n50774;
  assign n53543 = n53542 ^ n52196;
  assign n53548 = n53547 ^ n53543;
  assign n53596 = n53549 ^ n53548;
  assign n53593 = n53546 ^ n53544;
  assign n53594 = n50879 & n53593;
  assign n53595 = n53594 ^ n50887;
  assign n53646 = n53596 ^ n53595;
  assign n53597 = n53596 ^ n53594;
  assign n53598 = n53595 & n53597;
  assign n53599 = n53598 ^ n50887;
  assign n53550 = n53549 ^ n53543;
  assign n53551 = n53548 & n53550;
  assign n53552 = n53551 ^ n53547;
  assign n53539 = n52988 ^ n52211;
  assign n53540 = n53539 ^ n51481;
  assign n53590 = n53552 ^ n53540;
  assign n53501 = n53500 ^ n53308;
  assign n53502 = ~n53312 & n53501;
  assign n53503 = n53502 ^ n53311;
  assign n53304 = n51388 ^ n42468;
  assign n53305 = n53304 ^ n47715;
  assign n53306 = n53305 ^ n1408;
  assign n53537 = n53503 ^ n53306;
  assign n53224 = n53223 ^ n53098;
  assign n53225 = n53099 & n53224;
  assign n53226 = n53225 ^ n50070;
  assign n53095 = n52700 ^ n52592;
  assign n53092 = n52111 ^ n51457;
  assign n53093 = n53092 ^ n50866;
  assign n53089 = n53088 ^ n52921;
  assign n53090 = n52924 & n53089;
  assign n53091 = n53090 ^ n52923;
  assign n53094 = n53093 ^ n53091;
  assign n53096 = n53095 ^ n53094;
  assign n53097 = n53096 ^ n50095;
  assign n53296 = n53226 ^ n53097;
  assign n53295 = ~n53293 & n53294;
  assign n53303 = n53296 ^ n53295;
  assign n53538 = n53537 ^ n53303;
  assign n53591 = n53590 ^ n53538;
  assign n53592 = n53591 ^ n50894;
  assign n53647 = n53599 ^ n53592;
  assign n53648 = n53646 & ~n53647;
  assign n53600 = n53599 ^ n53591;
  assign n53601 = n53592 & ~n53600;
  assign n53602 = n53601 ^ n50894;
  assign n53541 = n53540 ^ n53538;
  assign n53553 = n53552 ^ n53538;
  assign n53554 = n53541 & n53553;
  assign n53555 = n53554 ^ n53540;
  assign n53307 = n53306 ^ n53303;
  assign n53504 = n53503 ^ n53303;
  assign n53505 = ~n53307 & n53504;
  assign n53506 = n53505 ^ n53306;
  assign n53299 = n51187 ^ n43849;
  assign n53300 = n53299 ^ n47933;
  assign n53301 = n53300 ^ n42427;
  assign n53534 = n53506 ^ n53301;
  assign n53297 = n53295 & ~n53296;
  assign n53235 = n52132 ^ n50791;
  assign n53236 = n53235 ^ n50837;
  assign n53234 = n52703 ^ n52587;
  assign n53237 = n53236 ^ n53234;
  assign n53230 = n53095 ^ n53093;
  assign n53231 = n53095 ^ n53091;
  assign n53232 = n53230 & n53231;
  assign n53233 = n53232 ^ n53093;
  assign n53238 = n53237 ^ n53233;
  assign n53239 = n53238 ^ n49664;
  assign n53227 = n53226 ^ n53096;
  assign n53228 = n53097 & n53227;
  assign n53229 = n53228 ^ n50095;
  assign n53240 = n53239 ^ n53229;
  assign n53298 = n53297 ^ n53240;
  assign n53535 = n53534 ^ n53298;
  assign n53532 = n53012 ^ n51488;
  assign n53533 = n53532 ^ n52317;
  assign n53536 = n53535 ^ n53533;
  assign n53588 = n53555 ^ n53536;
  assign n53589 = n53588 ^ n50788;
  assign n53649 = n53602 ^ n53589;
  assign n53650 = ~n53648 & n53649;
  assign n53603 = n53602 ^ n53588;
  assign n53604 = n53589 & n53603;
  assign n53605 = n53604 ^ n50788;
  assign n53556 = n53555 ^ n53533;
  assign n53557 = n53536 & ~n53556;
  assign n53558 = n53557 ^ n53535;
  assign n53529 = n52361 ^ n51549;
  assign n53530 = n53529 ^ n52982;
  assign n53524 = n50795 ^ n43877;
  assign n53525 = n53524 ^ n47710;
  assign n53526 = n53525 ^ n42477;
  assign n53518 = n52871 ^ n50785;
  assign n53517 = n52711 ^ n52710;
  assign n53519 = n53518 ^ n53517;
  assign n53514 = n53234 ^ n53233;
  assign n53515 = ~n53237 & n53514;
  assign n53516 = n53515 ^ n53236;
  assign n53520 = n53519 ^ n53516;
  assign n53511 = n53238 ^ n53229;
  assign n53512 = n53239 & ~n53511;
  assign n53513 = n53512 ^ n49664;
  assign n53521 = n53520 ^ n53513;
  assign n53522 = n53521 ^ n52106;
  assign n53510 = ~n53240 & ~n53297;
  assign n53523 = n53522 ^ n53510;
  assign n53527 = n53526 ^ n53523;
  assign n53302 = n53301 ^ n53298;
  assign n53507 = n53506 ^ n53298;
  assign n53508 = ~n53302 & n53507;
  assign n53509 = n53508 ^ n53301;
  assign n53528 = n53527 ^ n53509;
  assign n53531 = n53530 ^ n53528;
  assign n53586 = n53558 ^ n53531;
  assign n53587 = n53586 ^ n50781;
  assign n53645 = n53605 ^ n53587;
  assign n53760 = n53650 ^ n53645;
  assign n53756 = n51601 ^ n44335;
  assign n53757 = n53756 ^ n48117;
  assign n53758 = n53757 ^ n42739;
  assign n53748 = n51606 ^ n44340;
  assign n53749 = n53748 ^ n48133;
  assign n53750 = n53749 ^ n42743;
  assign n53740 = n51615 ^ n44345;
  assign n53741 = n53740 ^ n48121;
  assign n53742 = n53741 ^ n42753;
  assign n53733 = n51610 ^ n43752;
  assign n53734 = n53733 ^ n48124;
  assign n53735 = n53734 ^ n42749;
  assign n53728 = n52103 ^ n44520;
  assign n53729 = n53728 ^ n48675;
  assign n53730 = n53729 ^ n43204;
  assign n53731 = n53593 ^ n50879;
  assign n53732 = n53730 & n53731;
  assign n53736 = n53735 ^ n53732;
  assign n53737 = n53732 ^ n53646;
  assign n53738 = n53736 & ~n53737;
  assign n53739 = n53738 ^ n53735;
  assign n53743 = n53742 ^ n53739;
  assign n53744 = n53647 ^ n53646;
  assign n53745 = n53744 ^ n53739;
  assign n53746 = n53743 & ~n53745;
  assign n53747 = n53746 ^ n53742;
  assign n53751 = n53750 ^ n53747;
  assign n53752 = n53649 ^ n53648;
  assign n53753 = n53752 ^ n53747;
  assign n53754 = n53751 & n53753;
  assign n53755 = n53754 ^ n53750;
  assign n53759 = n53758 ^ n53755;
  assign n53845 = n53760 ^ n53759;
  assign n54978 = n53845 ^ n52912;
  assign n53639 = n53424 ^ n53412;
  assign n54979 = n54978 ^ n53639;
  assign n53885 = n52577 ^ n51700;
  assign n53886 = n53885 ^ n53076;
  assign n53827 = n53456 ^ n53371;
  assign n53828 = n53827 ^ n53368;
  assign n53887 = n53886 ^ n53828;
  assign n53888 = n52935 ^ n52562;
  assign n53889 = n53888 ^ n51704;
  assign n53833 = n53453 ^ n53450;
  assign n53890 = n53889 ^ n53833;
  assign n53893 = n53445 ^ n53377;
  assign n53891 = n52939 ^ n51793;
  assign n53892 = n53891 ^ n52548;
  assign n53894 = n53893 ^ n53892;
  assign n53897 = n52941 ^ n52534;
  assign n53898 = n53897 ^ n51708;
  assign n53895 = n53442 ^ n53380;
  assign n53896 = n53895 ^ n53381;
  assign n53899 = n53898 ^ n53896;
  assign n53902 = n52946 ^ n51783;
  assign n53903 = n53902 ^ n52520;
  assign n53900 = n53439 ^ n53385;
  assign n53901 = n53900 ^ n53386;
  assign n53904 = n53903 ^ n53901;
  assign n53809 = n53433 ^ n53397;
  assign n53687 = n52959 ^ n51766;
  assign n53688 = n53687 ^ n52452;
  assign n53686 = n53430 ^ n53402;
  assign n53689 = n53688 ^ n53686;
  assign n53673 = n52394 ^ n51759;
  assign n53674 = n53673 ^ n52964;
  assign n53672 = n53427 ^ n53407;
  assign n53675 = n53674 ^ n53672;
  assign n53637 = n52336 ^ n51752;
  assign n53638 = n53637 ^ n52965;
  assign n53640 = n53639 ^ n53638;
  assign n53577 = n53421 ^ n53420;
  assign n52893 = n52343 ^ n51720;
  assign n52895 = n52894 ^ n52893;
  assign n52853 = n52852 ^ n52849;
  assign n52892 = n52891 ^ n52853;
  assign n52896 = n52895 ^ n52892;
  assign n52900 = n52899 ^ n51722;
  assign n52901 = n52900 ^ n52347;
  assign n52897 = n52846 ^ n52825;
  assign n52898 = n52897 ^ n52822;
  assign n52902 = n52901 ^ n52898;
  assign n52905 = n52349 ^ n51723;
  assign n52907 = n52906 ^ n52905;
  assign n52903 = n52843 ^ n52830;
  assign n52904 = n52903 ^ n52827;
  assign n52908 = n52907 ^ n52904;
  assign n52913 = n52912 ^ n51730;
  assign n52914 = n52913 ^ n52353;
  assign n52909 = n52839 ^ n52748;
  assign n52910 = n52909 ^ n52836;
  assign n52915 = n52914 ^ n52910;
  assign n52918 = n52917 ^ n51674;
  assign n52919 = n52918 ^ n52357;
  assign n52916 = n52835 ^ n52834;
  assign n52920 = n52919 ^ n52916;
  assign n53559 = n53558 ^ n53528;
  assign n53560 = n53531 & n53559;
  assign n53561 = n53560 ^ n53530;
  assign n53562 = n53561 ^ n52916;
  assign n53563 = n52920 & n53562;
  assign n53564 = n53563 ^ n52919;
  assign n53565 = n53564 ^ n52910;
  assign n53566 = n52915 & ~n53565;
  assign n53567 = n53566 ^ n52914;
  assign n53568 = n53567 ^ n52904;
  assign n53569 = n52908 & ~n53568;
  assign n53570 = n53569 ^ n52907;
  assign n53571 = n53570 ^ n52898;
  assign n53572 = n52902 & n53571;
  assign n53573 = n53572 ^ n52901;
  assign n53574 = n53573 ^ n52892;
  assign n53575 = ~n52896 & n53574;
  assign n53576 = n53575 ^ n52895;
  assign n53578 = n53577 ^ n53576;
  assign n51686 = n51685 ^ n51684;
  assign n52330 = n52329 ^ n51686;
  assign n53634 = n53577 ^ n52330;
  assign n53635 = n53578 & ~n53634;
  assign n53636 = n53635 ^ n52330;
  assign n53669 = n53638 ^ n53636;
  assign n53670 = ~n53640 & n53669;
  assign n53671 = n53670 ^ n53639;
  assign n53683 = n53672 ^ n53671;
  assign n53684 = ~n53675 & ~n53683;
  assign n53685 = n53684 ^ n53674;
  assign n53806 = n53686 ^ n53685;
  assign n53807 = n53689 & ~n53806;
  assign n53808 = n53807 ^ n53688;
  assign n53810 = n53809 ^ n53808;
  assign n53804 = n52955 ^ n52465;
  assign n53805 = n53804 ^ n51713;
  assign n53905 = n53809 ^ n53805;
  assign n53906 = n53810 & ~n53905;
  assign n53907 = n53906 ^ n53805;
  assign n53837 = n53436 ^ n53390;
  assign n53838 = n53837 ^ n53391;
  assign n53908 = n53907 ^ n53838;
  assign n53909 = n52952 ^ n52505;
  assign n53910 = n53909 ^ n51776;
  assign n53911 = n53910 ^ n53838;
  assign n53912 = n53908 & ~n53911;
  assign n53913 = n53912 ^ n53910;
  assign n53914 = n53913 ^ n53901;
  assign n53915 = n53904 & n53914;
  assign n53916 = n53915 ^ n53903;
  assign n53917 = n53916 ^ n53896;
  assign n53918 = n53899 & ~n53917;
  assign n53919 = n53918 ^ n53898;
  assign n53920 = n53919 ^ n53893;
  assign n53921 = n53894 & ~n53920;
  assign n53922 = n53921 ^ n53892;
  assign n53923 = n53922 ^ n53833;
  assign n53924 = ~n53890 & n53923;
  assign n53925 = n53924 ^ n53889;
  assign n53926 = n53925 ^ n53828;
  assign n53927 = n53887 & n53926;
  assign n53928 = n53927 ^ n53886;
  assign n53882 = n52728 ^ n51696;
  assign n53883 = n53882 ^ n52929;
  assign n53820 = n53459 ^ n53366;
  assign n53821 = n53820 ^ n53363;
  assign n53884 = n53883 ^ n53821;
  assign n54019 = n53928 ^ n53884;
  assign n53983 = n53925 ^ n53887;
  assign n53984 = n53983 ^ n50986;
  assign n53985 = n53922 ^ n53890;
  assign n53986 = n53985 ^ n50979;
  assign n53987 = n53919 ^ n53892;
  assign n53988 = n53987 ^ n53893;
  assign n53989 = n53988 ^ n50798;
  assign n53990 = n53916 ^ n53899;
  assign n53991 = n53990 ^ n50804;
  assign n53992 = n53913 ^ n53903;
  assign n53993 = n53992 ^ n53901;
  assign n53994 = n53993 ^ n50966;
  assign n53995 = n53910 ^ n53908;
  assign n53996 = n53995 ^ n50808;
  assign n53811 = n53810 ^ n53805;
  assign n53812 = n53811 ^ n50813;
  assign n53690 = n53689 ^ n53685;
  assign n53691 = n53690 ^ n50953;
  assign n53676 = n53675 ^ n53671;
  assign n53641 = n53640 ^ n53636;
  assign n53579 = n53578 ^ n52330;
  assign n53580 = n53579 ^ n50822;
  assign n53625 = n53573 ^ n52895;
  assign n53626 = n53625 ^ n52892;
  assign n53615 = n53567 ^ n52908;
  assign n53581 = n53564 ^ n52915;
  assign n53582 = n53581 ^ n50777;
  assign n53583 = n53561 ^ n52919;
  assign n53584 = n53583 ^ n52916;
  assign n53585 = n53584 ^ n50913;
  assign n53606 = n53605 ^ n53586;
  assign n53607 = n53587 & ~n53606;
  assign n53608 = n53607 ^ n50781;
  assign n53609 = n53608 ^ n53584;
  assign n53610 = n53585 & n53609;
  assign n53611 = n53610 ^ n50913;
  assign n53612 = n53611 ^ n53581;
  assign n53613 = ~n53582 & n53612;
  assign n53614 = n53613 ^ n50777;
  assign n53616 = n53615 ^ n53614;
  assign n53617 = n53615 ^ n50828;
  assign n53618 = n53616 & n53617;
  assign n53619 = n53618 ^ n50828;
  assign n53620 = n53619 ^ n50929;
  assign n53621 = n53570 ^ n52902;
  assign n53622 = n53621 ^ n53619;
  assign n53623 = ~n53620 & ~n53622;
  assign n53624 = n53623 ^ n50929;
  assign n53627 = n53626 ^ n53624;
  assign n53628 = n53626 ^ n50824;
  assign n53629 = n53627 & n53628;
  assign n53630 = n53629 ^ n50824;
  assign n53631 = n53630 ^ n53579;
  assign n53632 = n53580 & ~n53631;
  assign n53633 = n53632 ^ n50822;
  assign n53642 = n53641 ^ n53633;
  assign n53666 = n53641 ^ n50942;
  assign n53667 = ~n53642 & n53666;
  assign n53668 = n53667 ^ n50942;
  assign n53677 = n53676 ^ n53668;
  assign n53680 = n53676 ^ n50818;
  assign n53681 = ~n53677 & ~n53680;
  assign n53682 = n53681 ^ n50818;
  assign n53801 = n53690 ^ n53682;
  assign n53802 = ~n53691 & n53801;
  assign n53803 = n53802 ^ n50953;
  assign n53997 = n53811 ^ n53803;
  assign n53998 = ~n53812 & ~n53997;
  assign n53999 = n53998 ^ n50813;
  assign n54000 = n53999 ^ n53995;
  assign n54001 = n53996 & n54000;
  assign n54002 = n54001 ^ n50808;
  assign n54003 = n54002 ^ n53993;
  assign n54004 = ~n53994 & n54003;
  assign n54005 = n54004 ^ n50966;
  assign n54006 = n54005 ^ n53990;
  assign n54007 = n53991 & ~n54006;
  assign n54008 = n54007 ^ n50804;
  assign n54009 = n54008 ^ n53988;
  assign n54010 = ~n53989 & ~n54009;
  assign n54011 = n54010 ^ n50798;
  assign n54012 = n54011 ^ n53985;
  assign n54013 = ~n53986 & ~n54012;
  assign n54014 = n54013 ^ n50979;
  assign n54015 = n54014 ^ n53983;
  assign n54016 = n53984 & ~n54015;
  assign n54017 = n54016 ^ n50986;
  assign n54018 = n54017 ^ n50993;
  assign n54065 = n54019 ^ n54018;
  assign n54066 = n54011 ^ n53986;
  assign n54067 = n54002 ^ n50966;
  assign n54068 = n54067 ^ n53993;
  assign n53813 = n53812 ^ n53803;
  assign n53643 = n53642 ^ n50942;
  assign n53644 = n53608 ^ n53585;
  assign n53651 = n53645 & ~n53650;
  assign n53652 = ~n53644 & ~n53651;
  assign n53653 = n53611 ^ n50777;
  assign n53654 = n53653 ^ n53581;
  assign n53655 = ~n53652 & n53654;
  assign n53656 = n53616 ^ n50828;
  assign n53657 = n53655 & ~n53656;
  assign n53658 = n53621 ^ n50929;
  assign n53659 = n53658 ^ n53619;
  assign n53660 = n53657 & ~n53659;
  assign n53661 = n53627 ^ n50824;
  assign n53662 = ~n53660 & n53661;
  assign n53663 = n53630 ^ n53580;
  assign n53664 = n53662 & ~n53663;
  assign n53665 = ~n53643 & n53664;
  assign n53678 = n53677 ^ n50818;
  assign n53679 = n53665 & n53678;
  assign n53692 = n53691 ^ n53682;
  assign n53814 = n53679 & ~n53692;
  assign n54069 = n53813 & ~n53814;
  assign n54070 = n53999 ^ n53996;
  assign n54071 = n54069 & n54070;
  assign n54072 = ~n54068 & ~n54071;
  assign n54073 = n54005 ^ n50804;
  assign n54074 = n54073 ^ n53990;
  assign n54075 = ~n54072 & ~n54074;
  assign n54076 = n54008 ^ n53989;
  assign n54077 = ~n54075 & ~n54076;
  assign n54078 = n54066 & n54077;
  assign n54079 = n54014 ^ n50986;
  assign n54080 = n54079 ^ n53983;
  assign n54081 = n54078 & n54080;
  assign n54082 = ~n54065 & ~n54081;
  assign n54020 = n54019 ^ n54017;
  assign n54021 = n54018 & ~n54020;
  assign n54022 = n54021 ^ n50993;
  assign n53929 = n53928 ^ n53883;
  assign n53930 = ~n53884 & ~n53929;
  assign n53931 = n53930 ^ n53821;
  assign n53880 = n53462 ^ n53362;
  assign n53878 = n52774 ^ n51809;
  assign n53879 = n53878 ^ n52925;
  assign n53881 = n53880 ^ n53879;
  assign n53981 = n53931 ^ n53881;
  assign n53982 = n53981 ^ n51128;
  assign n54083 = n54022 ^ n53982;
  assign n54084 = n54082 & n54083;
  assign n54023 = n54022 ^ n53981;
  assign n54024 = ~n53982 & ~n54023;
  assign n54025 = n54024 ^ n51128;
  assign n54085 = n54025 ^ n51401;
  assign n53936 = n53465 ^ n53357;
  assign n53876 = n52798 ^ n51899;
  assign n53877 = n53876 ^ n52921;
  assign n53978 = n53936 ^ n53877;
  assign n53932 = n53931 ^ n53880;
  assign n53933 = n53881 & n53932;
  assign n53934 = n53933 ^ n53879;
  assign n53979 = n53978 ^ n53934;
  assign n54086 = n54085 ^ n53979;
  assign n54087 = ~n54084 & n54086;
  assign n53942 = n52873 ^ n52090;
  assign n53943 = n53942 ^ n53095;
  assign n53940 = n53468 ^ n53352;
  assign n53935 = n53934 ^ n53877;
  assign n53937 = n53936 ^ n53934;
  assign n53938 = ~n53935 & n53937;
  assign n53939 = n53938 ^ n53877;
  assign n53941 = n53940 ^ n53939;
  assign n54029 = n53943 ^ n53941;
  assign n53980 = n53979 ^ n51401;
  assign n54026 = n54025 ^ n53979;
  assign n54027 = ~n53980 & ~n54026;
  assign n54028 = n54027 ^ n51401;
  assign n54030 = n54029 ^ n54028;
  assign n54088 = n54030 ^ n51445;
  assign n54089 = n54087 & ~n54088;
  assign n53950 = n53234 ^ n51419;
  assign n53951 = n53950 ^ n52117;
  assign n53947 = n53471 ^ n53346;
  assign n53948 = n53947 ^ n53343;
  assign n53944 = n53943 ^ n53940;
  assign n53945 = n53941 & ~n53944;
  assign n53946 = n53945 ^ n53943;
  assign n53949 = n53948 ^ n53946;
  assign n54034 = n53951 ^ n53949;
  assign n54031 = n54029 ^ n51445;
  assign n54032 = n54030 & ~n54031;
  assign n54033 = n54032 ^ n51445;
  assign n54035 = n54034 ^ n54033;
  assign n54064 = n54035 ^ n50642;
  assign n54207 = n54089 ^ n54064;
  assign n54199 = n54088 ^ n54087;
  assign n54125 = n51981 ^ n44271;
  assign n54126 = n54125 ^ n48452;
  assign n54127 = n54126 ^ n43110;
  assign n54124 = n54086 ^ n54084;
  assign n54128 = n54127 ^ n54124;
  assign n54188 = n51986 ^ n44276;
  assign n54189 = n54188 ^ n48457;
  assign n54190 = n54189 ^ n43066;
  assign n54180 = n54081 ^ n54065;
  assign n54130 = n52045 ^ n44425;
  assign n54131 = n54130 ^ n48468;
  assign n54132 = n54131 ^ n43075;
  assign n54129 = n54080 ^ n54078;
  assign n54133 = n54132 ^ n54129;
  assign n54135 = n51996 ^ n44285;
  assign n54136 = n54135 ^ n48530;
  assign n54137 = n54136 ^ n43081;
  assign n54134 = n54077 ^ n54066;
  assign n54138 = n54137 ^ n54134;
  assign n54142 = n54076 ^ n54075;
  assign n54139 = n52001 ^ n44291;
  assign n54140 = n54139 ^ n48473;
  assign n54141 = n54140 ^ n43086;
  assign n54143 = n54142 ^ n54141;
  assign n54144 = n54074 ^ n54072;
  assign n54148 = n54147 ^ n54144;
  assign n54160 = n54071 ^ n54068;
  assign n54152 = n54070 ^ n54069;
  assign n54149 = n52011 ^ n44306;
  assign n54150 = n54149 ^ n48488;
  assign n54151 = n54150 ^ n42705;
  assign n54153 = n54152 ^ n54151;
  assign n53815 = n53814 ^ n53813;
  assign n53694 = n51682 ^ n44313;
  assign n53695 = n53694 ^ n48495;
  assign n53696 = n53695 ^ n2245;
  assign n53693 = n53692 ^ n53679;
  assign n53697 = n53696 ^ n53693;
  assign n53790 = n53678 ^ n53665;
  assign n53699 = n51581 ^ n44320;
  assign n53700 = n53699 ^ n48178;
  assign n53701 = n53700 ^ n42719;
  assign n53698 = n53664 ^ n53643;
  assign n53702 = n53701 ^ n53698;
  assign n53706 = n53663 ^ n53662;
  assign n53703 = n51655 ^ n44390;
  assign n53704 = n53703 ^ n48087;
  assign n53705 = n53704 ^ n42793;
  assign n53707 = n53706 ^ n53705;
  assign n53709 = n51586 ^ n44382;
  assign n53710 = n53709 ^ n48092;
  assign n53711 = n53710 ^ n42723;
  assign n53708 = n53661 ^ n53660;
  assign n53712 = n53711 ^ n53708;
  assign n53714 = n51644 ^ n44374;
  assign n53715 = n53714 ^ n48097;
  assign n53716 = n53715 ^ n42782;
  assign n53713 = n53659 ^ n53657;
  assign n53717 = n53716 ^ n53713;
  assign n53721 = n53656 ^ n53655;
  assign n53718 = n51591 ^ n44325;
  assign n53719 = n53718 ^ n48102;
  assign n53720 = n53719 ^ n42728;
  assign n53722 = n53721 ^ n53720;
  assign n53726 = n53654 ^ n53652;
  assign n53723 = n51633 ^ n44363;
  assign n53724 = n53723 ^ n48107;
  assign n53725 = n53724 ^ n42771;
  assign n53727 = n53726 ^ n53725;
  assign n53764 = n53651 ^ n53644;
  assign n53761 = n53760 ^ n53755;
  assign n53762 = n53759 & ~n53761;
  assign n53763 = n53762 ^ n53758;
  assign n53765 = n53764 ^ n53763;
  assign n53766 = n51596 ^ n44330;
  assign n53767 = n53766 ^ n48112;
  assign n53768 = n53767 ^ n42734;
  assign n53769 = n53768 ^ n53764;
  assign n53770 = ~n53765 & n53769;
  assign n53771 = n53770 ^ n53768;
  assign n53772 = n53771 ^ n53725;
  assign n53773 = n53727 & ~n53772;
  assign n53774 = n53773 ^ n53726;
  assign n53775 = n53774 ^ n53720;
  assign n53776 = n53722 & ~n53775;
  assign n53777 = n53776 ^ n53721;
  assign n53778 = n53777 ^ n53713;
  assign n53779 = n53717 & ~n53778;
  assign n53780 = n53779 ^ n53716;
  assign n53781 = n53780 ^ n53708;
  assign n53782 = ~n53712 & n53781;
  assign n53783 = n53782 ^ n53711;
  assign n53784 = n53783 ^ n53705;
  assign n53785 = ~n53707 & ~n53784;
  assign n53786 = n53785 ^ n53706;
  assign n53787 = n53786 ^ n53698;
  assign n53788 = ~n53702 & ~n53787;
  assign n53789 = n53788 ^ n53701;
  assign n53791 = n53790 ^ n53789;
  assign n53792 = n51576 ^ n2055;
  assign n53793 = n53792 ^ n48500;
  assign n53794 = n53793 ^ n42714;
  assign n53795 = n53794 ^ n53790;
  assign n53796 = ~n53791 & n53795;
  assign n53797 = n53796 ^ n53794;
  assign n53798 = n53797 ^ n53693;
  assign n53799 = ~n53697 & n53798;
  assign n53800 = n53799 ^ n53696;
  assign n53816 = n53815 ^ n53800;
  assign n2217 = n2216 ^ n2159;
  assign n2254 = n2253 ^ n2217;
  assign n2264 = n2263 ^ n2254;
  assign n54154 = n53815 ^ n2264;
  assign n54155 = ~n53816 & n54154;
  assign n54156 = n54155 ^ n2264;
  assign n54157 = n54156 ^ n54151;
  assign n54158 = ~n54153 & ~n54157;
  assign n54159 = n54158 ^ n54152;
  assign n54161 = n54160 ^ n54159;
  assign n54162 = n52006 ^ n44301;
  assign n54163 = n54162 ^ n48483;
  assign n54164 = n54163 ^ n42700;
  assign n54165 = n54164 ^ n54160;
  assign n54166 = n54161 & n54165;
  assign n54167 = n54166 ^ n54164;
  assign n54168 = n54167 ^ n54144;
  assign n54169 = ~n54148 & n54168;
  assign n54170 = n54169 ^ n54147;
  assign n54171 = n54170 ^ n54142;
  assign n54172 = n54143 & ~n54171;
  assign n54173 = n54172 ^ n54141;
  assign n54174 = n54173 ^ n54134;
  assign n54175 = n54138 & ~n54174;
  assign n54176 = n54175 ^ n54137;
  assign n54177 = n54176 ^ n54129;
  assign n54178 = n54133 & ~n54177;
  assign n54179 = n54178 ^ n54132;
  assign n54181 = n54180 ^ n54179;
  assign n54182 = n51990 ^ n44280;
  assign n54183 = n54182 ^ n48462;
  assign n54184 = n54183 ^ n43070;
  assign n54185 = n54184 ^ n54180;
  assign n54186 = n54181 & ~n54185;
  assign n54187 = n54186 ^ n54184;
  assign n54191 = n54190 ^ n54187;
  assign n54192 = n54083 ^ n54082;
  assign n54193 = n54192 ^ n54187;
  assign n54194 = n54191 & n54193;
  assign n54195 = n54194 ^ n54190;
  assign n54196 = n54195 ^ n54124;
  assign n54197 = ~n54128 & n54196;
  assign n54198 = n54197 ^ n54127;
  assign n54200 = n54199 ^ n54198;
  assign n54201 = n51975 ^ n44266;
  assign n54202 = n54201 ^ n48448;
  assign n54203 = n54202 ^ n43061;
  assign n54204 = n54203 ^ n54199;
  assign n54205 = n54200 & ~n54204;
  assign n54206 = n54205 ^ n54203;
  assign n54208 = n54207 ^ n54206;
  assign n54209 = n51971 ^ n941;
  assign n54210 = n54209 ^ n48443;
  assign n54211 = n54210 ^ n43121;
  assign n54212 = n54211 ^ n54207;
  assign n54213 = ~n54208 & n54212;
  assign n54214 = n54213 ^ n54211;
  assign n54120 = n52068 ^ n44448;
  assign n54121 = n54120 ^ n48438;
  assign n54122 = n54121 ^ n1098;
  assign n54036 = n54034 ^ n50642;
  assign n54037 = ~n54035 & ~n54036;
  assign n54038 = n54037 ^ n50642;
  assign n53952 = n53951 ^ n53948;
  assign n53953 = n53949 & n53952;
  assign n53954 = n53953 ^ n53951;
  assign n53871 = n53517 ^ n51422;
  assign n53872 = n53871 ^ n52122;
  assign n53975 = n53954 ^ n53872;
  assign n53873 = n53474 ^ n53341;
  assign n53874 = n53873 ^ n53338;
  assign n53976 = n53975 ^ n53874;
  assign n53977 = n53976 ^ n50681;
  assign n54091 = n54038 ^ n53977;
  assign n54090 = n54064 & ~n54089;
  assign n54119 = n54091 ^ n54090;
  assign n54123 = n54122 ^ n54119;
  assign n54968 = n54214 ^ n54123;
  assign n54969 = n54968 ^ n52993;
  assign n54970 = n54969 ^ n44797;
  assign n54942 = n54211 ^ n54208;
  assign n54939 = n52995 ^ n52139;
  assign n54940 = n54939 ^ n53535;
  assign n54863 = n54203 ^ n54200;
  assign n54861 = n52883 ^ n52106;
  assign n54862 = n54861 ^ n53538;
  assign n54864 = n54863 ^ n54862;
  assign n54619 = n53549 ^ n52132;
  assign n54620 = n54619 ^ n52811;
  assign n54617 = n54195 ^ n54127;
  assign n54618 = n54617 ^ n54124;
  assign n54621 = n54620 ^ n54618;
  assign n54600 = n52780 ^ n52111;
  assign n54601 = n54600 ^ n53544;
  assign n54599 = n54192 ^ n54191;
  assign n54602 = n54601 ^ n54599;
  assign n54233 = n53494 ^ n53492;
  assign n54234 = n54233 ^ n53489;
  assign n54586 = n54234 ^ n52122;
  assign n54587 = n54586 ^ n52735;
  assign n54585 = n54184 ^ n54181;
  assign n54588 = n54587 ^ n54585;
  assign n54573 = n54176 ^ n54132;
  assign n54574 = n54573 ^ n54129;
  assign n54056 = n53486 ^ n53321;
  assign n54057 = n54056 ^ n53318;
  assign n54571 = n54057 ^ n52117;
  assign n54572 = n54571 ^ n52741;
  assign n54575 = n54574 ^ n54572;
  assign n53967 = n53483 ^ n53327;
  assign n54553 = n53967 ^ n53517;
  assign n54554 = n54553 ^ n52873;
  assign n54552 = n54173 ^ n54138;
  assign n54555 = n54554 ^ n54552;
  assign n54490 = n53234 ^ n52798;
  assign n53866 = n53480 ^ n53332;
  assign n54491 = n54490 ^ n53866;
  assign n54488 = n54170 ^ n54141;
  assign n54489 = n54488 ^ n54142;
  assign n54492 = n54491 ^ n54489;
  assign n53869 = n53477 ^ n53337;
  assign n54481 = n53869 ^ n53095;
  assign n54482 = n54481 ^ n52774;
  assign n54480 = n54167 ^ n54148;
  assign n54483 = n54482 ^ n54480;
  assign n54469 = n54164 ^ n54161;
  assign n54467 = n53874 ^ n52921;
  assign n54468 = n54467 ^ n52728;
  assign n54470 = n54469 ^ n54468;
  assign n54354 = n54156 ^ n54153;
  assign n54351 = n53948 ^ n52577;
  assign n54352 = n54351 ^ n52925;
  assign n54463 = n54354 ^ n54352;
  assign n54332 = n53794 ^ n53791;
  assign n53824 = n53786 ^ n53702;
  assign n53822 = n52939 ^ n52520;
  assign n53823 = n53822 ^ n53821;
  assign n53825 = n53824 ^ n53823;
  assign n53829 = n53828 ^ n52505;
  assign n53830 = n53829 ^ n52941;
  assign n53826 = n53783 ^ n53707;
  assign n53831 = n53830 ^ n53826;
  assign n53834 = n52946 ^ n52465;
  assign n53835 = n53834 ^ n53833;
  assign n53832 = n53780 ^ n53712;
  assign n53836 = n53835 ^ n53832;
  assign n54315 = n53777 ^ n53716;
  assign n54316 = n54315 ^ n53713;
  assign n54308 = n53774 ^ n53722;
  assign n54301 = n53771 ^ n53727;
  assign n53841 = n53768 ^ n53765;
  assign n53839 = n53838 ^ n52964;
  assign n53840 = n53839 ^ n51684;
  assign n53842 = n53841 ^ n53840;
  assign n53843 = n53809 ^ n52965;
  assign n53844 = n53843 ^ n52343;
  assign n53846 = n53845 ^ n53844;
  assign n53849 = n52347 ^ n52329;
  assign n53850 = n53849 ^ n53686;
  assign n53847 = n53752 ^ n53750;
  assign n53848 = n53847 ^ n53747;
  assign n53851 = n53850 ^ n53848;
  assign n53854 = n52894 ^ n52349;
  assign n53855 = n53854 ^ n53672;
  assign n53852 = n53744 ^ n53742;
  assign n53853 = n53852 ^ n53739;
  assign n53856 = n53855 ^ n53853;
  assign n53859 = n53639 ^ n52899;
  assign n53860 = n53859 ^ n52353;
  assign n53857 = n53735 ^ n53646;
  assign n53858 = n53857 ^ n53732;
  assign n53861 = n53860 ^ n53858;
  assign n53863 = n52906 ^ n52357;
  assign n53864 = n53863 ^ n53577;
  assign n53862 = n53731 ^ n53730;
  assign n53865 = n53864 ^ n53862;
  assign n54251 = n52912 ^ n52892;
  assign n54252 = n54251 ^ n52361;
  assign n54058 = n52811 ^ n50791;
  assign n54059 = n54058 ^ n52139;
  assign n54060 = n54059 ^ n54057;
  assign n53968 = n52780 ^ n52106;
  assign n53969 = n53968 ^ n51457;
  assign n53970 = n53969 ^ n53967;
  assign n53867 = n52111 ^ n51426;
  assign n53868 = n53867 ^ n52741;
  assign n53870 = n53869 ^ n53868;
  assign n53875 = n53874 ^ n53872;
  assign n53955 = n53954 ^ n53874;
  assign n53956 = ~n53875 & ~n53955;
  assign n53957 = n53956 ^ n53872;
  assign n53958 = n53957 ^ n53868;
  assign n53959 = n53870 & n53958;
  assign n53960 = n53959 ^ n53869;
  assign n53961 = n53960 ^ n53866;
  assign n53962 = n52132 ^ n51411;
  assign n53963 = n53962 ^ n52735;
  assign n53964 = n53963 ^ n53866;
  assign n53965 = n53961 & n53964;
  assign n53966 = n53965 ^ n53963;
  assign n54053 = n53967 ^ n53966;
  assign n54054 = ~n53970 & n54053;
  assign n54055 = n54054 ^ n53969;
  assign n54061 = n54060 ^ n54055;
  assign n54062 = n54061 ^ n50837;
  assign n53971 = n53970 ^ n53966;
  assign n53972 = n53971 ^ n50866;
  assign n54045 = n53963 ^ n53961;
  assign n53973 = n53957 ^ n53870;
  assign n53974 = n53973 ^ n50724;
  assign n54039 = n54038 ^ n53976;
  assign n54040 = ~n53977 & n54039;
  assign n54041 = n54040 ^ n50681;
  assign n54042 = n54041 ^ n53973;
  assign n54043 = ~n53974 & n54042;
  assign n54044 = n54043 ^ n50724;
  assign n54046 = n54045 ^ n54044;
  assign n54047 = n54045 ^ n50763;
  assign n54048 = ~n54046 & ~n54047;
  assign n54049 = n54048 ^ n50763;
  assign n54050 = n54049 ^ n53971;
  assign n54051 = ~n53972 & n54050;
  assign n54052 = n54051 ^ n50866;
  assign n54063 = n54062 ^ n54052;
  assign n54092 = ~n54090 & n54091;
  assign n54093 = n54041 ^ n53974;
  assign n54094 = ~n54092 & ~n54093;
  assign n54095 = n54046 ^ n50763;
  assign n54096 = ~n54094 & n54095;
  assign n54097 = n54049 ^ n53972;
  assign n54098 = n54096 & ~n54097;
  assign n54248 = n54063 & ~n54098;
  assign n54244 = n51691 ^ n44484;
  assign n54245 = n54244 ^ n48642;
  assign n54246 = n54245 ^ n43160;
  assign n54239 = n52147 ^ n50785;
  assign n54240 = n54239 ^ n52883;
  assign n54235 = n54057 ^ n54055;
  assign n54236 = n54060 & n54235;
  assign n54237 = n54236 ^ n54059;
  assign n54238 = n54237 ^ n54234;
  assign n54241 = n54240 ^ n54238;
  assign n54242 = n54241 ^ n50833;
  assign n54230 = n54061 ^ n54052;
  assign n54231 = ~n54062 & ~n54230;
  assign n54232 = n54231 ^ n50837;
  assign n54243 = n54242 ^ n54232;
  assign n54247 = n54246 ^ n54243;
  assign n54249 = n54248 ^ n54247;
  assign n54100 = n51950 ^ n43760;
  assign n54101 = n54100 ^ n48603;
  assign n54102 = n54101 ^ n43044;
  assign n54099 = n54098 ^ n54063;
  assign n54103 = n54102 ^ n54099;
  assign n54107 = n54097 ^ n54096;
  assign n54104 = n51955 ^ n44251;
  assign n54105 = n54104 ^ n48578;
  assign n54106 = n54105 ^ n43048;
  assign n54108 = n54107 ^ n54106;
  assign n54110 = n51960 ^ n44255;
  assign n54111 = n54110 ^ n48186;
  assign n54112 = n54111 ^ n1253;
  assign n54109 = n54095 ^ n54094;
  assign n54113 = n54112 ^ n54109;
  assign n54115 = n51965 ^ n44260;
  assign n54116 = n54115 ^ n1109;
  assign n54117 = n54116 ^ n43053;
  assign n54114 = n54093 ^ n54092;
  assign n54118 = n54117 ^ n54114;
  assign n54215 = n54214 ^ n54119;
  assign n54216 = ~n54123 & n54215;
  assign n54217 = n54216 ^ n54122;
  assign n54218 = n54217 ^ n54114;
  assign n54219 = ~n54118 & n54218;
  assign n54220 = n54219 ^ n54117;
  assign n54221 = n54220 ^ n54109;
  assign n54222 = ~n54113 & n54221;
  assign n54223 = n54222 ^ n54112;
  assign n54224 = n54223 ^ n54106;
  assign n54225 = ~n54108 & ~n54224;
  assign n54226 = n54225 ^ n54107;
  assign n54227 = n54226 ^ n54099;
  assign n54228 = n54103 & n54227;
  assign n54229 = n54228 ^ n54102;
  assign n54250 = n54249 ^ n54229;
  assign n54253 = n54252 ^ n54250;
  assign n54255 = n52917 ^ n52898;
  assign n54256 = n54255 ^ n52317;
  assign n54254 = n54226 ^ n54103;
  assign n54257 = n54256 ^ n54254;
  assign n54270 = n52982 ^ n52904;
  assign n54271 = n54270 ^ n52211;
  assign n54259 = n52910 ^ n52196;
  assign n54260 = n54259 ^ n53012;
  assign n54258 = n54220 ^ n54113;
  assign n54261 = n54260 ^ n54258;
  assign n54262 = n52988 ^ n52916;
  assign n54263 = n54262 ^ n52184;
  assign n54264 = n54217 ^ n54117;
  assign n54265 = n54264 ^ n54114;
  assign n54266 = n54263 & ~n54265;
  assign n54267 = n54266 ^ n54258;
  assign n54268 = ~n54261 & ~n54267;
  assign n54269 = n54268 ^ n54266;
  assign n54272 = n54271 ^ n54269;
  assign n54273 = n54223 ^ n54108;
  assign n54274 = n54273 ^ n54269;
  assign n54275 = ~n54272 & n54274;
  assign n54276 = n54275 ^ n54271;
  assign n54277 = n54276 ^ n54254;
  assign n54278 = ~n54257 & ~n54277;
  assign n54279 = n54278 ^ n54256;
  assign n54280 = n54279 ^ n54250;
  assign n54281 = n54253 & ~n54280;
  assign n54282 = n54281 ^ n54252;
  assign n54283 = n54282 ^ n53862;
  assign n54284 = ~n53865 & ~n54283;
  assign n54285 = n54284 ^ n53864;
  assign n54286 = n54285 ^ n53858;
  assign n54287 = ~n53861 & n54286;
  assign n54288 = n54287 ^ n53860;
  assign n54289 = n54288 ^ n53853;
  assign n54290 = ~n53856 & n54289;
  assign n54291 = n54290 ^ n53855;
  assign n54292 = n54291 ^ n53848;
  assign n54293 = ~n53851 & ~n54292;
  assign n54294 = n54293 ^ n53850;
  assign n54295 = n54294 ^ n53845;
  assign n54296 = ~n53846 & ~n54295;
  assign n54297 = n54296 ^ n53844;
  assign n54298 = n54297 ^ n53841;
  assign n54299 = n53842 & n54298;
  assign n54300 = n54299 ^ n53840;
  assign n54302 = n54301 ^ n54300;
  assign n54303 = n53901 ^ n52959;
  assign n54304 = n54303 ^ n52336;
  assign n54305 = n54304 ^ n54301;
  assign n54306 = ~n54302 & n54305;
  assign n54307 = n54306 ^ n54304;
  assign n54309 = n54308 ^ n54307;
  assign n54310 = n52955 ^ n52394;
  assign n54311 = n54310 ^ n53896;
  assign n54312 = n54311 ^ n54308;
  assign n54313 = ~n54309 & n54312;
  assign n54314 = n54313 ^ n54311;
  assign n54317 = n54316 ^ n54314;
  assign n54318 = n52952 ^ n52452;
  assign n54319 = n54318 ^ n53893;
  assign n54320 = n54319 ^ n54316;
  assign n54321 = ~n54317 & n54320;
  assign n54322 = n54321 ^ n54319;
  assign n54323 = n54322 ^ n53832;
  assign n54324 = ~n53836 & n54323;
  assign n54325 = n54324 ^ n53835;
  assign n54326 = n54325 ^ n53826;
  assign n54327 = n53831 & n54326;
  assign n54328 = n54327 ^ n53830;
  assign n54329 = n54328 ^ n53824;
  assign n54330 = n53825 & n54329;
  assign n54331 = n54330 ^ n53823;
  assign n54333 = n54332 ^ n54331;
  assign n54334 = n53880 ^ n52534;
  assign n54335 = n54334 ^ n52935;
  assign n54336 = n54335 ^ n54332;
  assign n54337 = ~n54333 & ~n54336;
  assign n54338 = n54337 ^ n54335;
  assign n53818 = n53797 ^ n53696;
  assign n53819 = n53818 ^ n53693;
  assign n54339 = n54338 ^ n53819;
  assign n54340 = n53076 ^ n52548;
  assign n54341 = n54340 ^ n53936;
  assign n54342 = n54341 ^ n53819;
  assign n54343 = ~n54339 & ~n54342;
  assign n54344 = n54343 ^ n54341;
  assign n53817 = n53816 ^ n2264;
  assign n54345 = n54344 ^ n53817;
  assign n54346 = n53940 ^ n52929;
  assign n54347 = n54346 ^ n52562;
  assign n54348 = n54347 ^ n53817;
  assign n54349 = ~n54345 & n54348;
  assign n54350 = n54349 ^ n54347;
  assign n54464 = n54354 ^ n54350;
  assign n54465 = ~n54463 & n54464;
  assign n54466 = n54465 ^ n54352;
  assign n54477 = n54468 ^ n54466;
  assign n54478 = n54470 & n54477;
  assign n54479 = n54478 ^ n54469;
  assign n54493 = n54480 ^ n54479;
  assign n54494 = ~n54483 & ~n54493;
  assign n54495 = n54494 ^ n54482;
  assign n54556 = n54495 ^ n54489;
  assign n54557 = ~n54492 & ~n54556;
  assign n54558 = n54557 ^ n54491;
  assign n54576 = n54558 ^ n54552;
  assign n54577 = ~n54555 & n54576;
  assign n54578 = n54577 ^ n54554;
  assign n54589 = n54578 ^ n54572;
  assign n54590 = ~n54575 & ~n54589;
  assign n54591 = n54590 ^ n54574;
  assign n54596 = n54591 ^ n54585;
  assign n54597 = n54588 & n54596;
  assign n54598 = n54597 ^ n54587;
  assign n54614 = n54599 ^ n54598;
  assign n54615 = n54602 & ~n54614;
  assign n54616 = n54615 ^ n54601;
  assign n54858 = n54618 ^ n54616;
  assign n54859 = ~n54621 & ~n54858;
  assign n54860 = n54859 ^ n54620;
  assign n54936 = n54862 ^ n54860;
  assign n54937 = ~n54864 & ~n54936;
  assign n54938 = n54937 ^ n54863;
  assign n54941 = n54940 ^ n54938;
  assign n54943 = n54942 ^ n54941;
  assign n54865 = n54864 ^ n54860;
  assign n54932 = n54865 ^ n51457;
  assign n54622 = n54621 ^ n54616;
  assign n54623 = n54622 ^ n51411;
  assign n54592 = n54591 ^ n54588;
  assign n54559 = n54558 ^ n54555;
  assign n54566 = n54559 ^ n52090;
  assign n54496 = n54495 ^ n54492;
  assign n54471 = n54470 ^ n54466;
  assign n54353 = n54352 ^ n54350;
  assign n54355 = n54354 ^ n54353;
  assign n54356 = n54355 ^ n51700;
  assign n54357 = n54347 ^ n54345;
  assign n54358 = n54357 ^ n51704;
  assign n54359 = n54341 ^ n54339;
  assign n54360 = n54359 ^ n51793;
  assign n54361 = n54335 ^ n54333;
  assign n54362 = n54361 ^ n51708;
  assign n54363 = n54328 ^ n53825;
  assign n54364 = n54363 ^ n51783;
  assign n54365 = n54325 ^ n53830;
  assign n54366 = n54365 ^ n53826;
  assign n54367 = n54366 ^ n51776;
  assign n54368 = n54322 ^ n53836;
  assign n54369 = n54368 ^ n51713;
  assign n54370 = n54319 ^ n54317;
  assign n54371 = n54370 ^ n51766;
  assign n54372 = n54311 ^ n54309;
  assign n54373 = n54372 ^ n51759;
  assign n54374 = n54304 ^ n54302;
  assign n54375 = n54374 ^ n51752;
  assign n54428 = n54297 ^ n53842;
  assign n54376 = n54294 ^ n53844;
  assign n54377 = n54376 ^ n53845;
  assign n54378 = n54377 ^ n51720;
  assign n54419 = n54291 ^ n53850;
  assign n54420 = n54419 ^ n53848;
  assign n54379 = n54288 ^ n53856;
  assign n54380 = n54379 ^ n51723;
  assign n54381 = n54285 ^ n53861;
  assign n54382 = n54381 ^ n51730;
  assign n54383 = n54282 ^ n53865;
  assign n54384 = n54383 ^ n51674;
  assign n54404 = n54279 ^ n54252;
  assign n54405 = n54404 ^ n54250;
  assign n54385 = n54276 ^ n54257;
  assign n54386 = n54385 ^ n51488;
  assign n54395 = n54273 ^ n54271;
  assign n54396 = n54395 ^ n54269;
  assign n54387 = n54265 ^ n54263;
  assign n54388 = n51471 & ~n54387;
  assign n54389 = n54388 ^ n50774;
  assign n54390 = n54266 ^ n54260;
  assign n54391 = n54390 ^ n54258;
  assign n54392 = n54391 ^ n54388;
  assign n54393 = ~n54389 & ~n54392;
  assign n54394 = n54393 ^ n50774;
  assign n54397 = n54396 ^ n54394;
  assign n54398 = n54396 ^ n51481;
  assign n54399 = n54397 & n54398;
  assign n54400 = n54399 ^ n51481;
  assign n54401 = n54400 ^ n54385;
  assign n54402 = ~n54386 & ~n54401;
  assign n54403 = n54402 ^ n51488;
  assign n54406 = n54405 ^ n54403;
  assign n54407 = n54405 ^ n51549;
  assign n54408 = n54406 & ~n54407;
  assign n54409 = n54408 ^ n51549;
  assign n54410 = n54409 ^ n54383;
  assign n54411 = n54384 & ~n54410;
  assign n54412 = n54411 ^ n51674;
  assign n54413 = n54412 ^ n54381;
  assign n54414 = ~n54382 & n54413;
  assign n54415 = n54414 ^ n51730;
  assign n54416 = n54415 ^ n54379;
  assign n54417 = n54380 & n54416;
  assign n54418 = n54417 ^ n51723;
  assign n54421 = n54420 ^ n54418;
  assign n54422 = n54420 ^ n51722;
  assign n54423 = ~n54421 & ~n54422;
  assign n54424 = n54423 ^ n51722;
  assign n54425 = n54424 ^ n54377;
  assign n54426 = ~n54378 & ~n54425;
  assign n54427 = n54426 ^ n51720;
  assign n54429 = n54428 ^ n54427;
  assign n54430 = n54427 ^ n51685;
  assign n54431 = n54429 & n54430;
  assign n54432 = n54431 ^ n51685;
  assign n54433 = n54432 ^ n54374;
  assign n54434 = ~n54375 & ~n54433;
  assign n54435 = n54434 ^ n51752;
  assign n54436 = n54435 ^ n54372;
  assign n54437 = n54373 & n54436;
  assign n54438 = n54437 ^ n51759;
  assign n54439 = n54438 ^ n54370;
  assign n54440 = n54371 & ~n54439;
  assign n54441 = n54440 ^ n51766;
  assign n54442 = n54441 ^ n54368;
  assign n54443 = n54369 & n54442;
  assign n54444 = n54443 ^ n51713;
  assign n54445 = n54444 ^ n54366;
  assign n54446 = n54367 & n54445;
  assign n54447 = n54446 ^ n51776;
  assign n54448 = n54447 ^ n54363;
  assign n54449 = ~n54364 & n54448;
  assign n54450 = n54449 ^ n51783;
  assign n54451 = n54450 ^ n54361;
  assign n54452 = n54362 & n54451;
  assign n54453 = n54452 ^ n51708;
  assign n54454 = n54453 ^ n54359;
  assign n54455 = ~n54360 & n54454;
  assign n54456 = n54455 ^ n51793;
  assign n54457 = n54456 ^ n54357;
  assign n54458 = ~n54358 & n54457;
  assign n54459 = n54458 ^ n51704;
  assign n54460 = n54459 ^ n54355;
  assign n54461 = ~n54356 & ~n54460;
  assign n54462 = n54461 ^ n51700;
  assign n54472 = n54471 ^ n54462;
  assign n54473 = n54471 ^ n51696;
  assign n54474 = ~n54472 & ~n54473;
  assign n54475 = n54474 ^ n51696;
  assign n54476 = n54475 ^ n51809;
  assign n54484 = n54483 ^ n54479;
  assign n54485 = n54484 ^ n54475;
  assign n54486 = ~n54476 & n54485;
  assign n54487 = n54486 ^ n51809;
  assign n54497 = n54496 ^ n54487;
  assign n54560 = n54496 ^ n51899;
  assign n54561 = n54497 & n54560;
  assign n54562 = n54561 ^ n51899;
  assign n54567 = n54562 ^ n54559;
  assign n54568 = n54566 & n54567;
  assign n54569 = n54568 ^ n52090;
  assign n54570 = n54569 ^ n51419;
  assign n54579 = n54578 ^ n54575;
  assign n54582 = n54579 ^ n54569;
  assign n54583 = n54570 & ~n54582;
  assign n54584 = n54583 ^ n51419;
  assign n54593 = n54592 ^ n54584;
  assign n54605 = n54592 ^ n51422;
  assign n54606 = ~n54593 & ~n54605;
  assign n54607 = n54606 ^ n51422;
  assign n54610 = n54607 ^ n51426;
  assign n54603 = n54602 ^ n54598;
  assign n54611 = n54607 ^ n54603;
  assign n54612 = n54610 & ~n54611;
  assign n54613 = n54612 ^ n51426;
  assign n54854 = n54622 ^ n54613;
  assign n54855 = n54623 & n54854;
  assign n54856 = n54855 ^ n51411;
  assign n54933 = n54865 ^ n54856;
  assign n54934 = ~n54932 & n54933;
  assign n54935 = n54934 ^ n51457;
  assign n54944 = n54943 ^ n54935;
  assign n54945 = n54944 ^ n50791;
  assign n54498 = n54497 ^ n51899;
  assign n54499 = n54472 ^ n51696;
  assign n54500 = n54453 ^ n51793;
  assign n54501 = n54500 ^ n54359;
  assign n54502 = n54450 ^ n51708;
  assign n54503 = n54502 ^ n54361;
  assign n54504 = n54415 ^ n54380;
  assign n54505 = n54397 ^ n51481;
  assign n54506 = n54391 ^ n54389;
  assign n54507 = n54505 & n54506;
  assign n54508 = n54400 ^ n54386;
  assign n54509 = ~n54507 & ~n54508;
  assign n54510 = n54406 ^ n51549;
  assign n54511 = ~n54509 & ~n54510;
  assign n54512 = n54409 ^ n54384;
  assign n54513 = ~n54511 & ~n54512;
  assign n54514 = n54412 ^ n54382;
  assign n54515 = ~n54513 & ~n54514;
  assign n54516 = n54504 & n54515;
  assign n54517 = n54421 ^ n51722;
  assign n54518 = n54516 & n54517;
  assign n54519 = n54424 ^ n54378;
  assign n54520 = ~n54518 & n54519;
  assign n54521 = n54429 ^ n51685;
  assign n54522 = n54520 & ~n54521;
  assign n54523 = n54432 ^ n51752;
  assign n54524 = n54523 ^ n54374;
  assign n54525 = n54522 & ~n54524;
  assign n54526 = n54435 ^ n51759;
  assign n54527 = n54526 ^ n54372;
  assign n54528 = n54525 & ~n54527;
  assign n54529 = n54438 ^ n51766;
  assign n54530 = n54529 ^ n54370;
  assign n54531 = n54528 & n54530;
  assign n54532 = n54441 ^ n51713;
  assign n54533 = n54532 ^ n54368;
  assign n54534 = ~n54531 & ~n54533;
  assign n54535 = n54444 ^ n51776;
  assign n54536 = n54535 ^ n54366;
  assign n54537 = n54534 & n54536;
  assign n54538 = n54447 ^ n54364;
  assign n54539 = ~n54537 & ~n54538;
  assign n54540 = ~n54503 & ~n54539;
  assign n54541 = n54501 & ~n54540;
  assign n54542 = n54456 ^ n51704;
  assign n54543 = n54542 ^ n54357;
  assign n54544 = n54541 & n54543;
  assign n54545 = n54459 ^ n54356;
  assign n54546 = n54544 & n54545;
  assign n54547 = n54499 & ~n54546;
  assign n54548 = n54484 ^ n51809;
  assign n54549 = n54548 ^ n54475;
  assign n54550 = n54547 & n54549;
  assign n54551 = n54498 & ~n54550;
  assign n54563 = n54562 ^ n52090;
  assign n54564 = n54563 ^ n54559;
  assign n54565 = n54551 & ~n54564;
  assign n54580 = n54579 ^ n54570;
  assign n54581 = ~n54565 & ~n54580;
  assign n54594 = n54593 ^ n51422;
  assign n54595 = ~n54581 & ~n54594;
  assign n54604 = n54603 ^ n51426;
  assign n54608 = n54607 ^ n54604;
  assign n54609 = ~n54595 & n54608;
  assign n54624 = n54623 ^ n54613;
  assign n54853 = ~n54609 & ~n54624;
  assign n54857 = n54856 ^ n51457;
  assign n54866 = n54865 ^ n54857;
  assign n54946 = n54853 & ~n54866;
  assign n54965 = n54945 & ~n54946;
  assign n54966 = n54965 ^ n43877;
  assign n54967 = n54966 ^ n52809;
  assign n54971 = n54970 ^ n54967;
  assign n54972 = n54971 ^ n49140;
  assign n54973 = n54972 ^ n54239;
  assign n54961 = n54942 ^ n54940;
  assign n54962 = n54942 ^ n54938;
  assign n54963 = n54961 & n54962;
  assign n54964 = n54963 ^ n54940;
  assign n54974 = n54973 ^ n54964;
  assign n54958 = n54943 ^ n50791;
  assign n54959 = n54944 & ~n54958;
  assign n54960 = n54959 ^ n50791;
  assign n54975 = n54974 ^ n54960;
  assign n54976 = n54975 ^ n53528;
  assign n54948 = n52763 ^ n44800;
  assign n54949 = n54948 ^ n49144;
  assign n54950 = n54949 ^ n43849;
  assign n54947 = n54946 ^ n54945;
  assign n54951 = n54950 ^ n54947;
  assign n54867 = n54866 ^ n54853;
  assign n54626 = n52333 ^ n45175;
  assign n54627 = n54626 ^ n49149;
  assign n54628 = n54627 ^ n1390;
  assign n54625 = n54624 ^ n54609;
  assign n54629 = n54628 ^ n54625;
  assign n54631 = n52709 ^ n1188;
  assign n54632 = n54631 ^ n49155;
  assign n54633 = n54632 ^ n43725;
  assign n54630 = n54608 ^ n54595;
  assign n54634 = n54633 ^ n54630;
  assign n54638 = n54594 ^ n54581;
  assign n54635 = n52586 ^ n45056;
  assign n54636 = n54635 ^ n49160;
  assign n54637 = n54636 ^ n43509;
  assign n54639 = n54638 ^ n54637;
  assign n54641 = n52591 ^ n45161;
  assign n54642 = n54641 ^ n49165;
  assign n54643 = n54642 ^ n43513;
  assign n54640 = n54580 ^ n54565;
  assign n54644 = n54643 ^ n54640;
  assign n54833 = n54564 ^ n54551;
  assign n54648 = n54550 ^ n54498;
  assign n54645 = n52596 ^ n45150;
  assign n54646 = n54645 ^ n49175;
  assign n54647 = n54646 ^ n43694;
  assign n54649 = n54648 ^ n54647;
  assign n54822 = n54549 ^ n54547;
  assign n54651 = n52683 ^ n45071;
  assign n54652 = n54651 ^ n49184;
  assign n54653 = n54652 ^ n43529;
  assign n54650 = n54546 ^ n54499;
  assign n54654 = n54653 ^ n54650;
  assign n54811 = n54545 ^ n54544;
  assign n54656 = n52611 ^ n45128;
  assign n54657 = n54656 ^ n49195;
  assign n54658 = n54657 ^ n43539;
  assign n54655 = n54543 ^ n54541;
  assign n54659 = n54658 ^ n54655;
  assign n54663 = n54540 ^ n54501;
  assign n54660 = n52616 ^ n45120;
  assign n54661 = n54660 ^ n49200;
  assign n54662 = n54661 ^ n43674;
  assign n54664 = n54663 ^ n54662;
  assign n54668 = n54539 ^ n54503;
  assign n54665 = n52620 ^ n45076;
  assign n54666 = n54665 ^ n49205;
  assign n54667 = n54666 ^ n43666;
  assign n54669 = n54668 ^ n54667;
  assign n54671 = n52626 ^ n45081;
  assign n54672 = n54671 ^ n49210;
  assign n54673 = n54672 ^ n43544;
  assign n54670 = n54538 ^ n54537;
  assign n54674 = n54673 ^ n54670;
  assign n54676 = n52631 ^ n45086;
  assign n54677 = n54676 ^ n49215;
  assign n54678 = n54677 ^ n43549;
  assign n54675 = n54536 ^ n54534;
  assign n54679 = n54678 ^ n54675;
  assign n54681 = n52636 ^ n45091;
  assign n54682 = n54681 ^ n49220;
  assign n54683 = n54682 ^ n43554;
  assign n54680 = n54533 ^ n54531;
  assign n54684 = n54683 ^ n54680;
  assign n54686 = n52652 ^ n45096;
  assign n54687 = n54686 ^ n49225;
  assign n54688 = n54687 ^ n43559;
  assign n54685 = n54530 ^ n54528;
  assign n54689 = n54688 ^ n54685;
  assign n54782 = n54527 ^ n54525;
  assign n54774 = n52311 ^ n44645;
  assign n54775 = n54774 ^ n49272;
  assign n54776 = n54775 ^ n43643;
  assign n54691 = n52236 ^ n44719;
  assign n54692 = n54691 ^ n49264;
  assign n54693 = n54692 ^ n1811;
  assign n54690 = n54521 ^ n54520;
  assign n54694 = n54693 ^ n54690;
  assign n54763 = n54519 ^ n54518;
  assign n54755 = n54517 ^ n54516;
  assign n54696 = n52251 ^ n44654;
  assign n54697 = n54696 ^ n49245;
  assign n54698 = n54697 ^ n43574;
  assign n54695 = n54515 ^ n54504;
  assign n54699 = n54698 ^ n54695;
  assign n54703 = n54514 ^ n54513;
  assign n54700 = n52293 ^ n44697;
  assign n54701 = n54700 ^ n48740;
  assign n54702 = n54701 ^ n43616;
  assign n54704 = n54703 ^ n54702;
  assign n54741 = n54512 ^ n54511;
  assign n54733 = n54510 ^ n54509;
  assign n54706 = n52277 ^ n44669;
  assign n54707 = n54706 ^ n48721;
  assign n54708 = n54707 ^ n43589;
  assign n54705 = n54508 ^ n54507;
  assign n54709 = n54708 ^ n54705;
  assign n54722 = n52270 ^ n44679;
  assign n54723 = n54722 ^ n48714;
  assign n54724 = n54723 ^ n43598;
  assign n54715 = n52266 ^ n44674;
  assign n54716 = n54715 ^ n48710;
  assign n54717 = n54716 ^ n43593;
  assign n54710 = n52879 ^ n45247;
  assign n54711 = n54710 ^ n49354;
  assign n54712 = n54711 ^ n2468;
  assign n54713 = n54387 ^ n51471;
  assign n54714 = n54712 & ~n54713;
  assign n54718 = n54717 ^ n54714;
  assign n54719 = n54714 ^ n54506;
  assign n54720 = n54718 & ~n54719;
  assign n54721 = n54720 ^ n54717;
  assign n54725 = n54724 ^ n54721;
  assign n54726 = n54506 ^ n54505;
  assign n54727 = n54726 ^ n54721;
  assign n54728 = n54725 & n54727;
  assign n54729 = n54728 ^ n54724;
  assign n54730 = n54729 ^ n54705;
  assign n54731 = n54709 & ~n54730;
  assign n54732 = n54731 ^ n54708;
  assign n54734 = n54733 ^ n54732;
  assign n54735 = n52261 ^ n44665;
  assign n54736 = n54735 ^ n48731;
  assign n54737 = n54736 ^ n43584;
  assign n54738 = n54737 ^ n54733;
  assign n54739 = n54734 & ~n54738;
  assign n54740 = n54739 ^ n54737;
  assign n54742 = n54741 ^ n54740;
  assign n54743 = n52256 ^ n44660;
  assign n54744 = n54743 ^ n48705;
  assign n54745 = n54744 ^ n43579;
  assign n54746 = n54745 ^ n54741;
  assign n54747 = ~n54742 & n54746;
  assign n54748 = n54747 ^ n54745;
  assign n54749 = n54748 ^ n54702;
  assign n54750 = ~n54704 & ~n54749;
  assign n54751 = n54750 ^ n54703;
  assign n54752 = n54751 ^ n54695;
  assign n54753 = ~n54699 & ~n54752;
  assign n54754 = n54753 ^ n54698;
  assign n54756 = n54755 ^ n54754;
  assign n54757 = n52246 ^ n44708;
  assign n54758 = n54757 ^ n49240;
  assign n54759 = n54758 ^ n43627;
  assign n54760 = n54759 ^ n54755;
  assign n54761 = n54756 & ~n54760;
  assign n54762 = n54761 ^ n54759;
  assign n54764 = n54763 ^ n54762;
  assign n54765 = n52241 ^ n44650;
  assign n54766 = n54765 ^ n49234;
  assign n54767 = n54766 ^ n43568;
  assign n54768 = n54767 ^ n54762;
  assign n54769 = n54764 & n54768;
  assign n54770 = n54769 ^ n54767;
  assign n54771 = n54770 ^ n54690;
  assign n54772 = ~n54694 & n54771;
  assign n54773 = n54772 ^ n54693;
  assign n54777 = n54776 ^ n54773;
  assign n54778 = n54524 ^ n54522;
  assign n54779 = n54778 ^ n54776;
  assign n54780 = ~n54777 & ~n54779;
  assign n54781 = n54780 ^ n54778;
  assign n54783 = n54782 ^ n54781;
  assign n54784 = n52641 ^ n44743;
  assign n54785 = n54784 ^ n49229;
  assign n54786 = n54785 ^ n43564;
  assign n54787 = n54786 ^ n54782;
  assign n54788 = ~n54783 & ~n54787;
  assign n54789 = n54788 ^ n54786;
  assign n54790 = n54789 ^ n54685;
  assign n54791 = n54689 & ~n54790;
  assign n54792 = n54791 ^ n54688;
  assign n54793 = n54792 ^ n54680;
  assign n54794 = ~n54684 & n54793;
  assign n54795 = n54794 ^ n54683;
  assign n54796 = n54795 ^ n54675;
  assign n54797 = ~n54679 & n54796;
  assign n54798 = n54797 ^ n54678;
  assign n54799 = n54798 ^ n54670;
  assign n54800 = n54674 & ~n54799;
  assign n54801 = n54800 ^ n54673;
  assign n54802 = n54801 ^ n54668;
  assign n54803 = ~n54669 & n54802;
  assign n54804 = n54803 ^ n54667;
  assign n54805 = n54804 ^ n54662;
  assign n54806 = ~n54664 & ~n54805;
  assign n54807 = n54806 ^ n54663;
  assign n54808 = n54807 ^ n54655;
  assign n54809 = n54659 & n54808;
  assign n54810 = n54809 ^ n54658;
  assign n54812 = n54811 ^ n54810;
  assign n54813 = n52606 ^ n45136;
  assign n54814 = n54813 ^ n49190;
  assign n54815 = n54814 ^ n43533;
  assign n54816 = n54815 ^ n54811;
  assign n54817 = ~n54812 & n54816;
  assign n54818 = n54817 ^ n54815;
  assign n54819 = n54818 ^ n54650;
  assign n54820 = n54654 & ~n54819;
  assign n54821 = n54820 ^ n54653;
  assign n54823 = n54822 ^ n54821;
  assign n54824 = n52601 ^ n45066;
  assign n54825 = n54824 ^ n49180;
  assign n54826 = n54825 ^ n43524;
  assign n54827 = n54826 ^ n54822;
  assign n54828 = n54823 & ~n54827;
  assign n54829 = n54828 ^ n54826;
  assign n54830 = n54829 ^ n54647;
  assign n54831 = ~n54649 & ~n54830;
  assign n54832 = n54831 ^ n54648;
  assign n54834 = n54833 ^ n54832;
  assign n54835 = n52697 ^ n45061;
  assign n54836 = n54835 ^ n49170;
  assign n54837 = n54836 ^ n43519;
  assign n54838 = n54837 ^ n54833;
  assign n54839 = ~n54834 & ~n54838;
  assign n54840 = n54839 ^ n54837;
  assign n54841 = n54840 ^ n54640;
  assign n54842 = ~n54644 & n54841;
  assign n54843 = n54842 ^ n54643;
  assign n54844 = n54843 ^ n54637;
  assign n54845 = n54639 & ~n54844;
  assign n54846 = n54845 ^ n54638;
  assign n54847 = n54846 ^ n54630;
  assign n54848 = n54634 & ~n54847;
  assign n54849 = n54848 ^ n54633;
  assign n54850 = n54849 ^ n54625;
  assign n54851 = n54629 & ~n54850;
  assign n54852 = n54851 ^ n54628;
  assign n54868 = n54867 ^ n54852;
  assign n1362 = n1361 ^ n1301;
  assign n1399 = n1398 ^ n1362;
  assign n1409 = n1408 ^ n1399;
  assign n54952 = n54867 ^ n1409;
  assign n54953 = n54868 & ~n54952;
  assign n54954 = n54953 ^ n1409;
  assign n54955 = n54954 ^ n54947;
  assign n54956 = n54951 & ~n54955;
  assign n54957 = n54956 ^ n54950;
  assign n54977 = n54976 ^ n54957;
  assign n54980 = n54979 ^ n54977;
  assign n54999 = n53577 ^ n52917;
  assign n55000 = n54999 ^ n53848;
  assign n54983 = n54846 ^ n54633;
  assign n54984 = n54983 ^ n54630;
  assign n54985 = n53862 ^ n52988;
  assign n54986 = n54985 ^ n52904;
  assign n54987 = n54984 & ~n54986;
  assign n54981 = n53012 ^ n52898;
  assign n54982 = n54981 ^ n53858;
  assign n54988 = n54987 ^ n54982;
  assign n54989 = n54849 ^ n54629;
  assign n54990 = n54989 ^ n54982;
  assign n54991 = n54988 & ~n54990;
  assign n54992 = n54991 ^ n54987;
  assign n54869 = n54868 ^ n1409;
  assign n54993 = n54992 ^ n54869;
  assign n54994 = n53853 ^ n52982;
  assign n54995 = n54994 ^ n52892;
  assign n54996 = n54995 ^ n54869;
  assign n54997 = n54993 & ~n54996;
  assign n54998 = n54997 ^ n54995;
  assign n55001 = n55000 ^ n54998;
  assign n55002 = n54954 ^ n54951;
  assign n55003 = n55002 ^ n54998;
  assign n55004 = n55001 & ~n55003;
  assign n55005 = n55004 ^ n55000;
  assign n55006 = n55005 ^ n54977;
  assign n55007 = ~n54980 & ~n55006;
  assign n55008 = n55007 ^ n54979;
  assign n54929 = n53841 ^ n53672;
  assign n54930 = n54929 ^ n52906;
  assign n54928 = n54713 ^ n54712;
  assign n54931 = n54930 ^ n54928;
  assign n55108 = n55008 ^ n54931;
  assign n55084 = n55005 ^ n54979;
  assign n55085 = n55084 ^ n54977;
  assign n55086 = n55085 ^ n52361;
  assign n55087 = n55002 ^ n55000;
  assign n55088 = n55087 ^ n54998;
  assign n55089 = n55088 ^ n52317;
  assign n55090 = n54995 ^ n54993;
  assign n55091 = n55090 ^ n52211;
  assign n55092 = n54986 ^ n54984;
  assign n55093 = ~n52184 & ~n55092;
  assign n55094 = n55093 ^ n52196;
  assign n55095 = n54989 ^ n54988;
  assign n55096 = n55095 ^ n55093;
  assign n55097 = n55094 & ~n55096;
  assign n55098 = n55097 ^ n52196;
  assign n55099 = n55098 ^ n55090;
  assign n55100 = n55091 & n55099;
  assign n55101 = n55100 ^ n52211;
  assign n55102 = n55101 ^ n55088;
  assign n55103 = n55089 & n55102;
  assign n55104 = n55103 ^ n52317;
  assign n55105 = n55104 ^ n55085;
  assign n55106 = ~n55086 & n55105;
  assign n55107 = n55106 ^ n52361;
  assign n55109 = n55108 ^ n55107;
  assign n55177 = n55109 ^ n52357;
  assign n55178 = n55095 ^ n55094;
  assign n55179 = n55098 ^ n55091;
  assign n55180 = ~n55178 & ~n55179;
  assign n55181 = n55101 ^ n55089;
  assign n55182 = ~n55180 & ~n55181;
  assign n55183 = n55104 ^ n55086;
  assign n55184 = ~n55182 & n55183;
  assign n55185 = n55177 & ~n55184;
  assign n55110 = n55108 ^ n52357;
  assign n55111 = ~n55109 & n55110;
  assign n55112 = n55111 ^ n52357;
  assign n55009 = n55008 ^ n54928;
  assign n55010 = ~n54931 & ~n55009;
  assign n55011 = n55010 ^ n54930;
  assign n54925 = n54301 ^ n52899;
  assign n54926 = n54925 ^ n53686;
  assign n55081 = n55011 ^ n54926;
  assign n54923 = n54717 ^ n54506;
  assign n54924 = n54923 ^ n54714;
  assign n55082 = n55081 ^ n54924;
  assign n55083 = n55082 ^ n52353;
  assign n55186 = n55112 ^ n55083;
  assign n55187 = ~n55185 & ~n55186;
  assign n54927 = n54926 ^ n54924;
  assign n55012 = n55011 ^ n54924;
  assign n55013 = ~n54927 & ~n55012;
  assign n55014 = n55013 ^ n54926;
  assign n54920 = n53809 ^ n52894;
  assign n54921 = n54920 ^ n54308;
  assign n55116 = n55014 ^ n54921;
  assign n54918 = n54726 ^ n54724;
  assign n54919 = n54918 ^ n54721;
  assign n55117 = n55116 ^ n54919;
  assign n55113 = n55112 ^ n55082;
  assign n55114 = n55083 & n55113;
  assign n55115 = n55114 ^ n52353;
  assign n55118 = n55117 ^ n55115;
  assign n55188 = n55118 ^ n52349;
  assign n55189 = n55187 & ~n55188;
  assign n55119 = n55117 ^ n52349;
  assign n55120 = n55118 & ~n55119;
  assign n55121 = n55120 ^ n52349;
  assign n54922 = n54921 ^ n54919;
  assign n55015 = n55014 ^ n54919;
  assign n55016 = ~n54922 & ~n55015;
  assign n55017 = n55016 ^ n54921;
  assign n54915 = n54316 ^ n53838;
  assign n54916 = n54915 ^ n52329;
  assign n54913 = n54729 ^ n54708;
  assign n54914 = n54913 ^ n54705;
  assign n54917 = n54916 ^ n54914;
  assign n55079 = n55017 ^ n54917;
  assign n55080 = n55079 ^ n52347;
  assign n55190 = n55121 ^ n55080;
  assign n55191 = n55189 & ~n55190;
  assign n55122 = n55121 ^ n55079;
  assign n55123 = ~n55080 & n55122;
  assign n55124 = n55123 ^ n52347;
  assign n55018 = n55017 ^ n54914;
  assign n55019 = n54917 & ~n55018;
  assign n55020 = n55019 ^ n54916;
  assign n54910 = n53832 ^ n52965;
  assign n54911 = n54910 ^ n53901;
  assign n55076 = n55020 ^ n54911;
  assign n54909 = n54737 ^ n54734;
  assign n55077 = n55076 ^ n54909;
  assign n55078 = n55077 ^ n52343;
  assign n55176 = n55124 ^ n55078;
  assign n55321 = n55191 ^ n55176;
  assign n55325 = n55324 ^ n55321;
  assign n55329 = n55190 ^ n55189;
  assign n55326 = n53406 ^ n45530;
  assign n55327 = n55326 ^ n49533;
  assign n55328 = n55327 ^ n44374;
  assign n55330 = n55329 ^ n55328;
  assign n55383 = n55188 ^ n55187;
  assign n55332 = n53419 ^ n45575;
  assign n55333 = n55332 ^ n49580;
  assign n55334 = n55333 ^ n44363;
  assign n55331 = n55186 ^ n55185;
  assign n55335 = n55334 ^ n55331;
  assign n55337 = n52852 ^ n45541;
  assign n55338 = n55337 ^ n49543;
  assign n55339 = n55338 ^ n44330;
  assign n55336 = n55184 ^ n55177;
  assign n55340 = n55339 ^ n55336;
  assign n55342 = n52825 ^ n45546;
  assign n55343 = n55342 ^ n49569;
  assign n55344 = n55343 ^ n44335;
  assign n55341 = n55183 ^ n55182;
  assign n55345 = n55344 ^ n55341;
  assign n55366 = n52830 ^ n45559;
  assign n55367 = n55366 ^ n49561;
  assign n55368 = n55367 ^ n44340;
  assign n55358 = n55179 ^ n55178;
  assign n55351 = n52834 ^ n2543;
  assign n55352 = n55351 ^ n49547;
  assign n55353 = n55352 ^ n43752;
  assign n55346 = n53526 ^ n45895;
  assign n55347 = n55346 ^ n50088;
  assign n55348 = n55347 ^ n44520;
  assign n55349 = n55092 ^ n52184;
  assign n55350 = n55348 & n55349;
  assign n55354 = n55353 ^ n55350;
  assign n55355 = n55350 ^ n55178;
  assign n55356 = n55354 & n55355;
  assign n55357 = n55356 ^ n55353;
  assign n55359 = n55358 ^ n55357;
  assign n55360 = n52839 ^ n45552;
  assign n55361 = n55360 ^ n49552;
  assign n55362 = n55361 ^ n44345;
  assign n55363 = n55362 ^ n55357;
  assign n55364 = n55359 & n55363;
  assign n55365 = n55364 ^ n55362;
  assign n55369 = n55368 ^ n55365;
  assign n55370 = n55181 ^ n55180;
  assign n55371 = n55370 ^ n55365;
  assign n55372 = n55369 & ~n55371;
  assign n55373 = n55372 ^ n55368;
  assign n55374 = n55373 ^ n55341;
  assign n55375 = n55345 & ~n55374;
  assign n55376 = n55375 ^ n55344;
  assign n55377 = n55376 ^ n55336;
  assign n55378 = ~n55340 & n55377;
  assign n55379 = n55378 ^ n55339;
  assign n55380 = n55379 ^ n55331;
  assign n55381 = ~n55335 & n55380;
  assign n55382 = n55381 ^ n55334;
  assign n55384 = n55383 ^ n55382;
  assign n55385 = n53410 ^ n45536;
  assign n55386 = n55385 ^ n49538;
  assign n55387 = n55386 ^ n44325;
  assign n55388 = n55387 ^ n55383;
  assign n55389 = ~n55384 & n55388;
  assign n55390 = n55389 ^ n55387;
  assign n55391 = n55390 ^ n55328;
  assign n55392 = n55330 & ~n55391;
  assign n55393 = n55392 ^ n55329;
  assign n55394 = n55393 ^ n55321;
  assign n55395 = ~n55325 & n55394;
  assign n55396 = n55395 ^ n55324;
  assign n55317 = n53396 ^ n45520;
  assign n55318 = n55317 ^ n49523;
  assign n55319 = n55318 ^ n44390;
  assign n54912 = n54911 ^ n54909;
  assign n55021 = n55020 ^ n54909;
  assign n55022 = ~n54912 & n55021;
  assign n55023 = n55022 ^ n54911;
  assign n54906 = n53896 ^ n52964;
  assign n54907 = n54906 ^ n53826;
  assign n54905 = n54745 ^ n54742;
  assign n54908 = n54907 ^ n54905;
  assign n55128 = n55023 ^ n54908;
  assign n55125 = n55124 ^ n55077;
  assign n55126 = ~n55078 & ~n55125;
  assign n55127 = n55126 ^ n52343;
  assign n55129 = n55128 ^ n55127;
  assign n55193 = n55129 ^ n51684;
  assign n55192 = n55176 & ~n55191;
  assign n55316 = n55193 ^ n55192;
  assign n55320 = n55319 ^ n55316;
  assign n55765 = n55396 ^ n55320;
  assign n55057 = n54792 ^ n54684;
  assign n55511 = n55057 ^ n54469;
  assign n55512 = n55511 ^ n53821;
  assign n55509 = n55393 ^ n55324;
  assign n55510 = n55509 ^ n55321;
  assign n55513 = n55512 ^ n55510;
  assign n55048 = n54789 ^ n54689;
  assign n55515 = n55048 ^ n53828;
  assign n55516 = n55515 ^ n54354;
  assign n55514 = n55390 ^ n55330;
  assign n55517 = n55516 ^ n55514;
  assign n55752 = n55387 ^ n55384;
  assign n55745 = n55379 ^ n55335;
  assign n55738 = n54332 ^ n53896;
  assign n54885 = n54770 ^ n54693;
  assign n54886 = n54885 ^ n54690;
  assign n55739 = n55738 ^ n54886;
  assign n54890 = n54767 ^ n54764;
  assign n55519 = n54890 ^ n53824;
  assign n55520 = n55519 ^ n53901;
  assign n55518 = n55373 ^ n55345;
  assign n55521 = n55520 ^ n55518;
  assign n55728 = n55370 ^ n55369;
  assign n55721 = n55362 ^ n55359;
  assign n55713 = n55353 ^ n55178;
  assign n55714 = n55713 ^ n55350;
  assign n55706 = n55349 ^ n55348;
  assign n55670 = n53301 ^ n45737;
  assign n55671 = n55670 ^ n50052;
  assign n55672 = n55671 ^ n44484;
  assign n55642 = n52995 ^ n52916;
  assign n55643 = n55642 ^ n54254;
  assign n55620 = n54273 ^ n53528;
  assign n55621 = n55620 ^ n52883;
  assign n55619 = n54837 ^ n54834;
  assign n55622 = n55621 ^ n55619;
  assign n55599 = n54258 ^ n53535;
  assign n55600 = n55599 ^ n52811;
  assign n55477 = n54829 ^ n54649;
  assign n55601 = n55600 ^ n55477;
  assign n55581 = n53538 ^ n52780;
  assign n55582 = n55581 ^ n54265;
  assign n55483 = n54826 ^ n54823;
  assign n55583 = n55582 ^ n55483;
  assign n55535 = n54942 ^ n52741;
  assign n55536 = n55535 ^ n53544;
  assign n55447 = n54863 ^ n54234;
  assign n55448 = n55447 ^ n53517;
  assign n55445 = n54807 ^ n54658;
  assign n55446 = n55445 ^ n54655;
  assign n55449 = n55448 ^ n55446;
  assign n55249 = n54804 ^ n54664;
  assign n55234 = n53967 ^ n53095;
  assign n55235 = n55234 ^ n54599;
  assign n55233 = n54801 ^ n54669;
  assign n55236 = n55235 ^ n55233;
  assign n55221 = n54798 ^ n54674;
  assign n55218 = n54585 ^ n52921;
  assign n55219 = n55218 ^ n53866;
  assign n55229 = n55221 ^ n55219;
  assign n55168 = n54795 ^ n54679;
  assign n55055 = n54552 ^ n53874;
  assign n55056 = n55055 ^ n52929;
  assign n55058 = n55057 ^ n55056;
  assign n54876 = n53940 ^ n52935;
  assign n54877 = n54876 ^ n54480;
  assign n54875 = n54786 ^ n54783;
  assign n54878 = n54877 ^ n54875;
  assign n54880 = n53936 ^ n52939;
  assign n54881 = n54880 ^ n54469;
  assign n54879 = n54778 ^ n54777;
  assign n54882 = n54881 ^ n54879;
  assign n54883 = n54354 ^ n52941;
  assign n54884 = n54883 ^ n53880;
  assign n54887 = n54886 ^ n54884;
  assign n54888 = n53821 ^ n53817;
  assign n54889 = n54888 ^ n52946;
  assign n54891 = n54890 ^ n54889;
  assign n54893 = n53828 ^ n52952;
  assign n54894 = n54893 ^ n53819;
  assign n54892 = n54759 ^ n54756;
  assign n54895 = n54894 ^ n54892;
  assign n54898 = n54751 ^ n54698;
  assign n54899 = n54898 ^ n54695;
  assign n54896 = n54332 ^ n53833;
  assign n54897 = n54896 ^ n52955;
  assign n54900 = n54899 ^ n54897;
  assign n54902 = n53824 ^ n52959;
  assign n54903 = n54902 ^ n53893;
  assign n54901 = n54748 ^ n54704;
  assign n54904 = n54903 ^ n54901;
  assign n55024 = n55023 ^ n54905;
  assign n55025 = ~n54908 & ~n55024;
  assign n55026 = n55025 ^ n54907;
  assign n55027 = n55026 ^ n54901;
  assign n55028 = n54904 & ~n55027;
  assign n55029 = n55028 ^ n54903;
  assign n55030 = n55029 ^ n54897;
  assign n55031 = n54900 & n55030;
  assign n55032 = n55031 ^ n54899;
  assign n55033 = n55032 ^ n54892;
  assign n55034 = ~n54895 & n55033;
  assign n55035 = n55034 ^ n54894;
  assign n55036 = n55035 ^ n54890;
  assign n55037 = ~n54891 & n55036;
  assign n55038 = n55037 ^ n54889;
  assign n55039 = n55038 ^ n54884;
  assign n55040 = n54887 & n55039;
  assign n55041 = n55040 ^ n54886;
  assign n55042 = n55041 ^ n54879;
  assign n55043 = n54882 & ~n55042;
  assign n55044 = n55043 ^ n54881;
  assign n55045 = n55044 ^ n54875;
  assign n55046 = n54878 & n55045;
  assign n55047 = n55046 ^ n54877;
  assign n55049 = n55048 ^ n55047;
  assign n55050 = n54489 ^ n53076;
  assign n55051 = n55050 ^ n53948;
  assign n55052 = n55051 ^ n55048;
  assign n55053 = ~n55049 & n55052;
  assign n55054 = n55053 ^ n55051;
  assign n55165 = n55057 ^ n55054;
  assign n55166 = n55058 & n55165;
  assign n55167 = n55166 ^ n55056;
  assign n55169 = n55168 ^ n55167;
  assign n55163 = n54574 ^ n52925;
  assign n55164 = n55163 ^ n53869;
  assign n55215 = n55168 ^ n55164;
  assign n55216 = ~n55169 & ~n55215;
  assign n55217 = n55216 ^ n55164;
  assign n55230 = n55221 ^ n55217;
  assign n55231 = ~n55229 & ~n55230;
  assign n55232 = n55231 ^ n55219;
  assign n55246 = n55233 ^ n55232;
  assign n55247 = n55236 & ~n55246;
  assign n55248 = n55247 ^ n55235;
  assign n55250 = n55249 ^ n55248;
  assign n55244 = n54057 ^ n53234;
  assign n55245 = n55244 ^ n54618;
  assign n55442 = n55249 ^ n55245;
  assign n55443 = ~n55250 & ~n55442;
  assign n55444 = n55443 ^ n55245;
  assign n55532 = n55446 ^ n55444;
  assign n55533 = n55449 & n55532;
  assign n55534 = n55533 ^ n55448;
  assign n55537 = n55536 ^ n55534;
  assign n55530 = n54815 ^ n54810;
  assign n55531 = n55530 ^ n54811;
  assign n55555 = n55536 ^ n55531;
  assign n55556 = n55537 & n55555;
  assign n55557 = n55556 ^ n55534;
  assign n55487 = n54818 ^ n54654;
  assign n55558 = n55557 ^ n55487;
  assign n55553 = n54968 ^ n52735;
  assign n55554 = n55553 ^ n53549;
  assign n55578 = n55554 ^ n55487;
  assign n55579 = n55558 & n55578;
  assign n55580 = n55579 ^ n55554;
  assign n55596 = n55580 ^ n55483;
  assign n55597 = ~n55583 & n55596;
  assign n55598 = n55597 ^ n55582;
  assign n55616 = n55598 ^ n55477;
  assign n55617 = n55601 & n55616;
  assign n55618 = n55617 ^ n55600;
  assign n55638 = n55619 ^ n55618;
  assign n55639 = n55622 & n55638;
  assign n55640 = n55639 ^ n55621;
  assign n55470 = n54840 ^ n54644;
  assign n55641 = n55640 ^ n55470;
  assign n55644 = n55643 ^ n55641;
  assign n55645 = n55644 ^ n52139;
  assign n55623 = n55622 ^ n55618;
  assign n55602 = n55601 ^ n55598;
  assign n55584 = n55583 ^ n55580;
  assign n55585 = n55584 ^ n52111;
  assign n55559 = n55558 ^ n55554;
  assign n55560 = n55559 ^ n52122;
  assign n55538 = n55537 ^ n55531;
  assign n55539 = n55538 ^ n52117;
  assign n55450 = n55449 ^ n55444;
  assign n55451 = n55450 ^ n52873;
  assign n55251 = n55250 ^ n55245;
  assign n55237 = n55236 ^ n55232;
  assign n55238 = n55237 ^ n52774;
  assign n55220 = n55219 ^ n55217;
  assign n55222 = n55221 ^ n55220;
  assign n55170 = n55169 ^ n55164;
  assign n55211 = n55170 ^ n52577;
  assign n55059 = n55058 ^ n55054;
  assign n55060 = n55059 ^ n52562;
  assign n55061 = n55051 ^ n55049;
  assign n55062 = n55061 ^ n52548;
  assign n55063 = n55044 ^ n54877;
  assign n55064 = n55063 ^ n54875;
  assign n55065 = n55064 ^ n52534;
  assign n55066 = n55041 ^ n54882;
  assign n55067 = n55066 ^ n52520;
  assign n55068 = n55038 ^ n54887;
  assign n55069 = n55068 ^ n52505;
  assign n55070 = n55035 ^ n54891;
  assign n55071 = n55070 ^ n52465;
  assign n55072 = n55032 ^ n54895;
  assign n55073 = n55072 ^ n52452;
  assign n55074 = n55026 ^ n54904;
  assign n55075 = n55074 ^ n52336;
  assign n55130 = n55128 ^ n51684;
  assign n55131 = n55129 & ~n55130;
  assign n55132 = n55131 ^ n51684;
  assign n55133 = n55132 ^ n55074;
  assign n55134 = n55075 & n55133;
  assign n55135 = n55134 ^ n52336;
  assign n55136 = n55135 ^ n52394;
  assign n55137 = n55029 ^ n54900;
  assign n55138 = n55137 ^ n55135;
  assign n55139 = n55136 & ~n55138;
  assign n55140 = n55139 ^ n52394;
  assign n55141 = n55140 ^ n55072;
  assign n55142 = ~n55073 & ~n55141;
  assign n55143 = n55142 ^ n52452;
  assign n55144 = n55143 ^ n55070;
  assign n55145 = n55071 & n55144;
  assign n55146 = n55145 ^ n52465;
  assign n55147 = n55146 ^ n55068;
  assign n55148 = ~n55069 & n55147;
  assign n55149 = n55148 ^ n52505;
  assign n55150 = n55149 ^ n55066;
  assign n55151 = ~n55067 & ~n55150;
  assign n55152 = n55151 ^ n52520;
  assign n55153 = n55152 ^ n55064;
  assign n55154 = ~n55065 & n55153;
  assign n55155 = n55154 ^ n52534;
  assign n55156 = n55155 ^ n55061;
  assign n55157 = ~n55062 & ~n55156;
  assign n55158 = n55157 ^ n52548;
  assign n55159 = n55158 ^ n55059;
  assign n55160 = ~n55060 & n55159;
  assign n55161 = n55160 ^ n52562;
  assign n55212 = n55170 ^ n55161;
  assign n55213 = n55211 & n55212;
  assign n55214 = n55213 ^ n52577;
  assign n55223 = n55222 ^ n55214;
  assign n55226 = n55222 ^ n52728;
  assign n55227 = n55223 & ~n55226;
  assign n55228 = n55227 ^ n52728;
  assign n55241 = n55237 ^ n55228;
  assign n55242 = ~n55238 & n55241;
  assign n55243 = n55242 ^ n52774;
  assign n55252 = n55251 ^ n55243;
  assign n55439 = n55251 ^ n52798;
  assign n55440 = ~n55252 & ~n55439;
  assign n55441 = n55440 ^ n52798;
  assign n55527 = n55450 ^ n55441;
  assign n55528 = ~n55451 & n55527;
  assign n55529 = n55528 ^ n52873;
  assign n55550 = n55538 ^ n55529;
  assign n55551 = ~n55539 & n55550;
  assign n55552 = n55551 ^ n52117;
  assign n55575 = n55559 ^ n55552;
  assign n55576 = ~n55560 & ~n55575;
  assign n55577 = n55576 ^ n52122;
  assign n55593 = n55584 ^ n55577;
  assign n55594 = n55585 & n55593;
  assign n55595 = n55594 ^ n52111;
  assign n55603 = n55602 ^ n55595;
  assign n55613 = n55602 ^ n52132;
  assign n55614 = n55603 & n55613;
  assign n55615 = n55614 ^ n52132;
  assign n55624 = n55623 ^ n55615;
  assign n55635 = n55623 ^ n52106;
  assign n55636 = n55624 & ~n55635;
  assign n55637 = n55636 ^ n52106;
  assign n55646 = n55645 ^ n55637;
  assign n55625 = n55624 ^ n52106;
  assign n55586 = n55585 ^ n55577;
  assign n55561 = n55560 ^ n55552;
  assign n55540 = n55539 ^ n55529;
  assign n55452 = n55451 ^ n55441;
  assign n55162 = n55161 ^ n52577;
  assign n55171 = n55170 ^ n55162;
  assign n55172 = n55146 ^ n55069;
  assign n55173 = n55140 ^ n55073;
  assign n55174 = n55137 ^ n52394;
  assign n55175 = n55174 ^ n55135;
  assign n55194 = n55192 & ~n55193;
  assign n55195 = n55132 ^ n55075;
  assign n55196 = n55194 & n55195;
  assign n55197 = ~n55175 & n55196;
  assign n55198 = n55173 & n55197;
  assign n55199 = n55143 ^ n55071;
  assign n55200 = ~n55198 & ~n55199;
  assign n55201 = ~n55172 & n55200;
  assign n55202 = n55149 ^ n55067;
  assign n55203 = ~n55201 & n55202;
  assign n55204 = n55152 ^ n55065;
  assign n55205 = ~n55203 & n55204;
  assign n55206 = n55155 ^ n55062;
  assign n55207 = ~n55205 & ~n55206;
  assign n55208 = n55158 ^ n55060;
  assign n55209 = n55207 & n55208;
  assign n55210 = ~n55171 & n55209;
  assign n55224 = n55223 ^ n52728;
  assign n55225 = ~n55210 & n55224;
  assign n55239 = n55238 ^ n55228;
  assign n55240 = n55225 & n55239;
  assign n55253 = n55252 ^ n52798;
  assign n55453 = ~n55240 & ~n55253;
  assign n55541 = n55452 & n55453;
  assign n55562 = ~n55540 & ~n55541;
  assign n55587 = n55561 & ~n55562;
  assign n55592 = ~n55586 & ~n55587;
  assign n55604 = n55603 ^ n52132;
  assign n55626 = ~n55592 & ~n55604;
  assign n55647 = ~n55625 & n55626;
  assign n55669 = ~n55646 & ~n55647;
  assign n55673 = n55672 ^ n55669;
  assign n55663 = n54250 ^ n52910;
  assign n55664 = n55663 ^ n52993;
  assign n55662 = n54843 ^ n54639;
  assign n55665 = n55664 ^ n55662;
  assign n55659 = n55643 ^ n55470;
  assign n55660 = n55641 & n55659;
  assign n55661 = n55660 ^ n55643;
  assign n55666 = n55665 ^ n55661;
  assign n55667 = n55666 ^ n52147;
  assign n55656 = n55644 ^ n55637;
  assign n55657 = n55645 & ~n55656;
  assign n55658 = n55657 ^ n52139;
  assign n55668 = n55667 ^ n55658;
  assign n55674 = n55673 ^ n55668;
  assign n55648 = n55647 ^ n55646;
  assign n55627 = n55626 ^ n55625;
  assign n55605 = n55604 ^ n55592;
  assign n55571 = n53492 ^ n45856;
  assign n55572 = n55571 ^ n49862;
  assign n55573 = n55572 ^ n44260;
  assign n55563 = n55562 ^ n55561;
  assign n55542 = n55541 ^ n55540;
  assign n55455 = n53331 ^ n45668;
  assign n55456 = n55455 ^ n49877;
  assign n55457 = n55456 ^ n44266;
  assign n55454 = n55453 ^ n55452;
  assign n55458 = n55457 ^ n55454;
  assign n55254 = n55253 ^ n55240;
  assign n54872 = n53336 ^ n45662;
  assign n54873 = n54872 ^ n49882;
  assign n54874 = n54873 ^ n44271;
  assign n55255 = n55254 ^ n54874;
  assign n55257 = n53341 ^ n45481;
  assign n55258 = n55257 ^ n49887;
  assign n55259 = n55258 ^ n44276;
  assign n55256 = n55239 ^ n55225;
  assign n55260 = n55259 ^ n55256;
  assign n55262 = n53346 ^ n45637;
  assign n55263 = n55262 ^ n49892;
  assign n55264 = n55263 ^ n44280;
  assign n55261 = n55224 ^ n55210;
  assign n55265 = n55264 ^ n55261;
  assign n55267 = n53350 ^ n45486;
  assign n55268 = n55267 ^ n49896;
  assign n55269 = n55268 ^ n44425;
  assign n55266 = n55209 ^ n55171;
  assign n55270 = n55269 ^ n55266;
  assign n55272 = n53356 ^ n45491;
  assign n55273 = n55272 ^ n49902;
  assign n55274 = n55273 ^ n44285;
  assign n55271 = n55208 ^ n55207;
  assign n55275 = n55274 ^ n55271;
  assign n55277 = n53361 ^ n45495;
  assign n55278 = n55277 ^ n49907;
  assign n55279 = n55278 ^ n44291;
  assign n55276 = n55206 ^ n55205;
  assign n55280 = n55279 ^ n55276;
  assign n55282 = n53366 ^ n45501;
  assign n55283 = n55282 ^ n49912;
  assign n55284 = n55283 ^ n44296;
  assign n55281 = n55204 ^ n55203;
  assign n55285 = n55284 ^ n55281;
  assign n55287 = n53371 ^ n45615;
  assign n55288 = n55287 ^ n49917;
  assign n55289 = n55288 ^ n44301;
  assign n55286 = n55202 ^ n55201;
  assign n55290 = n55289 ^ n55286;
  assign n55292 = n53453 ^ n45506;
  assign n55293 = n55292 ^ n49926;
  assign n55294 = n55293 ^ n44306;
  assign n55291 = n55200 ^ n55172;
  assign n55295 = n55294 ^ n55291;
  assign n55297 = n53376 ^ n45604;
  assign n55298 = n55297 ^ n49627;
  assign n55299 = n55298 ^ n2216;
  assign n55296 = n55199 ^ n55198;
  assign n55300 = n55299 ^ n55296;
  assign n55302 = n53380 ^ n45511;
  assign n55303 = n55302 ^ n2066;
  assign n55304 = n55303 ^ n44313;
  assign n55301 = n55197 ^ n55173;
  assign n55305 = n55304 ^ n55301;
  assign n55307 = n53385 ^ n49518;
  assign n55308 = n55307 ^ n45515;
  assign n55309 = n55308 ^ n2055;
  assign n55306 = n55196 ^ n55175;
  assign n55310 = n55309 ^ n55306;
  assign n55314 = n55195 ^ n55194;
  assign n55311 = n53390 ^ n1892;
  assign n55312 = n55311 ^ n49598;
  assign n55313 = n55312 ^ n44320;
  assign n55315 = n55314 ^ n55313;
  assign n55397 = n55396 ^ n55316;
  assign n55398 = ~n55320 & n55397;
  assign n55399 = n55398 ^ n55319;
  assign n55400 = n55399 ^ n55313;
  assign n55401 = n55315 & ~n55400;
  assign n55402 = n55401 ^ n55314;
  assign n55403 = n55402 ^ n55306;
  assign n55404 = ~n55310 & n55403;
  assign n55405 = n55404 ^ n55309;
  assign n55406 = n55405 ^ n55301;
  assign n55407 = n55305 & ~n55406;
  assign n55408 = n55407 ^ n55304;
  assign n55409 = n55408 ^ n55296;
  assign n55410 = ~n55300 & n55409;
  assign n55411 = n55410 ^ n55299;
  assign n55412 = n55411 ^ n55291;
  assign n55413 = n55295 & ~n55412;
  assign n55414 = n55413 ^ n55294;
  assign n55415 = n55414 ^ n55286;
  assign n55416 = ~n55290 & n55415;
  assign n55417 = n55416 ^ n55289;
  assign n55418 = n55417 ^ n55281;
  assign n55419 = n55285 & ~n55418;
  assign n55420 = n55419 ^ n55284;
  assign n55421 = n55420 ^ n55276;
  assign n55422 = n55280 & ~n55421;
  assign n55423 = n55422 ^ n55279;
  assign n55424 = n55423 ^ n55271;
  assign n55425 = n55275 & ~n55424;
  assign n55426 = n55425 ^ n55274;
  assign n55427 = n55426 ^ n55266;
  assign n55428 = ~n55270 & n55427;
  assign n55429 = n55428 ^ n55269;
  assign n55430 = n55429 ^ n55261;
  assign n55431 = n55265 & ~n55430;
  assign n55432 = n55431 ^ n55264;
  assign n55433 = n55432 ^ n55256;
  assign n55434 = ~n55260 & n55433;
  assign n55435 = n55434 ^ n55259;
  assign n55436 = n55435 ^ n54874;
  assign n55437 = n55255 & ~n55436;
  assign n55438 = n55437 ^ n55254;
  assign n55524 = n55454 ^ n55438;
  assign n55525 = n55458 & ~n55524;
  assign n55526 = n55525 ^ n55457;
  assign n55543 = n55542 ^ n55526;
  assign n55544 = n53325 ^ n45866;
  assign n55545 = n55544 ^ n49871;
  assign n55546 = n55545 ^ n941;
  assign n55547 = n55546 ^ n55542;
  assign n55548 = n55543 & ~n55547;
  assign n55549 = n55548 ^ n55546;
  assign n55564 = n55563 ^ n55549;
  assign n55565 = n53321 ^ n45860;
  assign n55566 = n55565 ^ n49867;
  assign n55567 = n55566 ^ n44448;
  assign n55568 = n55567 ^ n55563;
  assign n55569 = n55564 & ~n55568;
  assign n55570 = n55569 ^ n55567;
  assign n55574 = n55573 ^ n55570;
  assign n55588 = n55587 ^ n55586;
  assign n55589 = n55588 ^ n55570;
  assign n55590 = n55574 & n55589;
  assign n55591 = n55590 ^ n55573;
  assign n55606 = n55605 ^ n55591;
  assign n55607 = n53316 ^ n45850;
  assign n55608 = n55607 ^ n49670;
  assign n55609 = n55608 ^ n44255;
  assign n55610 = n55609 ^ n55605;
  assign n55611 = ~n55606 & n55610;
  assign n55612 = n55611 ^ n55609;
  assign n55628 = n55627 ^ n55612;
  assign n55629 = n53311 ^ n45845;
  assign n55630 = n55629 ^ n49989;
  assign n55631 = n55630 ^ n44251;
  assign n55632 = n55631 ^ n55627;
  assign n55633 = n55628 & ~n55632;
  assign n55634 = n55633 ^ n55631;
  assign n55649 = n55648 ^ n55634;
  assign n55650 = n53306 ^ n45840;
  assign n55651 = n55650 ^ n50019;
  assign n55652 = n55651 ^ n43760;
  assign n55653 = n55652 ^ n55648;
  assign n55654 = n55649 & ~n55653;
  assign n55655 = n55654 ^ n55652;
  assign n55675 = n55674 ^ n55655;
  assign n55522 = n54909 ^ n54301;
  assign n55523 = n55522 ^ n53639;
  assign n55676 = n55675 ^ n55523;
  assign n55696 = n55652 ^ n55649;
  assign n55689 = n55631 ^ n55628;
  assign n55679 = n55588 ^ n55573;
  assign n55680 = n55679 ^ n55570;
  assign n55681 = n54928 ^ n53853;
  assign n55682 = n55681 ^ n52904;
  assign n55683 = ~n55680 & n55682;
  assign n55677 = n53848 ^ n52898;
  assign n55678 = n55677 ^ n54924;
  assign n55684 = n55683 ^ n55678;
  assign n55685 = n55609 ^ n55606;
  assign n55686 = n55685 ^ n55678;
  assign n55687 = ~n55684 & n55686;
  assign n55688 = n55687 ^ n55683;
  assign n55690 = n55689 ^ n55688;
  assign n55691 = n54919 ^ n52892;
  assign n55692 = n55691 ^ n53845;
  assign n55693 = n55692 ^ n55689;
  assign n55694 = n55690 & ~n55693;
  assign n55695 = n55694 ^ n55692;
  assign n55697 = n55696 ^ n55695;
  assign n55698 = n53841 ^ n53577;
  assign n55699 = n55698 ^ n54914;
  assign n55700 = n55699 ^ n55696;
  assign n55701 = n55697 & n55700;
  assign n55702 = n55701 ^ n55699;
  assign n55703 = n55702 ^ n55675;
  assign n55704 = n55676 & ~n55703;
  assign n55705 = n55704 ^ n55523;
  assign n55707 = n55706 ^ n55705;
  assign n55708 = n54905 ^ n54308;
  assign n55709 = n55708 ^ n53672;
  assign n55710 = n55709 ^ n55706;
  assign n55711 = n55707 & n55710;
  assign n55712 = n55711 ^ n55709;
  assign n55715 = n55714 ^ n55712;
  assign n55716 = n54901 ^ n53686;
  assign n55717 = n55716 ^ n54316;
  assign n55718 = n55717 ^ n55714;
  assign n55719 = n55715 & ~n55718;
  assign n55720 = n55719 ^ n55717;
  assign n55722 = n55721 ^ n55720;
  assign n55723 = n53832 ^ n53809;
  assign n55724 = n55723 ^ n54899;
  assign n55725 = n55724 ^ n55721;
  assign n55726 = n55722 & n55725;
  assign n55727 = n55726 ^ n55724;
  assign n55729 = n55728 ^ n55727;
  assign n55730 = n54892 ^ n53838;
  assign n55731 = n55730 ^ n53826;
  assign n55732 = n55731 ^ n55728;
  assign n55733 = n55729 & n55732;
  assign n55734 = n55733 ^ n55731;
  assign n55735 = n55734 ^ n55518;
  assign n55736 = ~n55521 & ~n55735;
  assign n55737 = n55736 ^ n55520;
  assign n55740 = n55739 ^ n55737;
  assign n55741 = n55376 ^ n55340;
  assign n55742 = n55741 ^ n55737;
  assign n55743 = n55740 & ~n55742;
  assign n55744 = n55743 ^ n55739;
  assign n55746 = n55745 ^ n55744;
  assign n55747 = n54879 ^ n53819;
  assign n55748 = n55747 ^ n53893;
  assign n55749 = n55748 ^ n55745;
  assign n55750 = ~n55746 & ~n55749;
  assign n55751 = n55750 ^ n55748;
  assign n55753 = n55752 ^ n55751;
  assign n55754 = n54875 ^ n53817;
  assign n55755 = n55754 ^ n53833;
  assign n55756 = n55755 ^ n55752;
  assign n55757 = ~n55753 & ~n55756;
  assign n55758 = n55757 ^ n55755;
  assign n55759 = n55758 ^ n55514;
  assign n55760 = n55517 & n55759;
  assign n55761 = n55760 ^ n55516;
  assign n55762 = n55761 ^ n55510;
  assign n55763 = ~n55513 & n55762;
  assign n55764 = n55763 ^ n55512;
  assign n55766 = n55765 ^ n55764;
  assign n55767 = n55168 ^ n54480;
  assign n55768 = n55767 ^ n53880;
  assign n55769 = n55768 ^ n55765;
  assign n55770 = n55766 & n55769;
  assign n55771 = n55770 ^ n55768;
  assign n55506 = n55221 ^ n54489;
  assign n55507 = n55506 ^ n53936;
  assign n55505 = n55399 ^ n55315;
  assign n55508 = n55507 ^ n55505;
  assign n55853 = n55771 ^ n55508;
  assign n55854 = n55853 ^ n52939;
  assign n55855 = n55768 ^ n55766;
  assign n55856 = n55855 ^ n52941;
  assign n55857 = n55761 ^ n55513;
  assign n55858 = n55857 ^ n52946;
  assign n55859 = n55758 ^ n55516;
  assign n55860 = n55859 ^ n55514;
  assign n55861 = n55860 ^ n52952;
  assign n55862 = n55755 ^ n55753;
  assign n55863 = n55862 ^ n52955;
  assign n55864 = n55748 ^ n55746;
  assign n55865 = n55864 ^ n52959;
  assign n55914 = n55741 ^ n55739;
  assign n55915 = n55914 ^ n55737;
  assign n55866 = n55734 ^ n55521;
  assign n55867 = n55866 ^ n52965;
  assign n55868 = n55731 ^ n55729;
  assign n55869 = n55868 ^ n52329;
  assign n55870 = n55724 ^ n55722;
  assign n55871 = n55870 ^ n52894;
  assign n55872 = n55717 ^ n55715;
  assign n55873 = n55872 ^ n52899;
  assign n55897 = n55709 ^ n55707;
  assign n55874 = n55702 ^ n55523;
  assign n55875 = n55874 ^ n55675;
  assign n55876 = n55875 ^ n52912;
  assign n55877 = n55699 ^ n55697;
  assign n55878 = n55877 ^ n52917;
  assign n55879 = n55692 ^ n55690;
  assign n55880 = n55879 ^ n52982;
  assign n55881 = n55682 ^ n55680;
  assign n55882 = n52988 & ~n55881;
  assign n55883 = n55882 ^ n53012;
  assign n55884 = n55685 ^ n55684;
  assign n55885 = n55884 ^ n55882;
  assign n55886 = n55883 & n55885;
  assign n55887 = n55886 ^ n53012;
  assign n55888 = n55887 ^ n55879;
  assign n55889 = n55880 & n55888;
  assign n55890 = n55889 ^ n52982;
  assign n55891 = n55890 ^ n55877;
  assign n55892 = n55878 & n55891;
  assign n55893 = n55892 ^ n52917;
  assign n55894 = n55893 ^ n55875;
  assign n55895 = n55876 & n55894;
  assign n55896 = n55895 ^ n52912;
  assign n55898 = n55897 ^ n55896;
  assign n55899 = n55897 ^ n52906;
  assign n55900 = ~n55898 & ~n55899;
  assign n55901 = n55900 ^ n52906;
  assign n55902 = n55901 ^ n55872;
  assign n55903 = ~n55873 & n55902;
  assign n55904 = n55903 ^ n52899;
  assign n55905 = n55904 ^ n55870;
  assign n55906 = n55871 & ~n55905;
  assign n55907 = n55906 ^ n52894;
  assign n55908 = n55907 ^ n55868;
  assign n55909 = ~n55869 & n55908;
  assign n55910 = n55909 ^ n52329;
  assign n55911 = n55910 ^ n55866;
  assign n55912 = n55867 & n55911;
  assign n55913 = n55912 ^ n52965;
  assign n55916 = n55915 ^ n55913;
  assign n55917 = n55915 ^ n52964;
  assign n55918 = ~n55916 & ~n55917;
  assign n55919 = n55918 ^ n52964;
  assign n55920 = n55919 ^ n55864;
  assign n55921 = ~n55865 & ~n55920;
  assign n55922 = n55921 ^ n52959;
  assign n55923 = n55922 ^ n55862;
  assign n55924 = n55863 & ~n55923;
  assign n55925 = n55924 ^ n52955;
  assign n55926 = n55925 ^ n55860;
  assign n55927 = ~n55861 & ~n55926;
  assign n55928 = n55927 ^ n52952;
  assign n55929 = n55928 ^ n55857;
  assign n55930 = ~n55858 & n55929;
  assign n55931 = n55930 ^ n52946;
  assign n55932 = n55931 ^ n55855;
  assign n55933 = ~n55856 & ~n55932;
  assign n55934 = n55933 ^ n52941;
  assign n55935 = n55934 ^ n55853;
  assign n55936 = ~n55854 & ~n55935;
  assign n55937 = n55936 ^ n52939;
  assign n55938 = n55937 ^ n52935;
  assign n55772 = n55771 ^ n55505;
  assign n55773 = n55508 & n55772;
  assign n55774 = n55773 ^ n55507;
  assign n55503 = n55402 ^ n55310;
  assign n55501 = n55233 ^ n53940;
  assign n55502 = n55501 ^ n54552;
  assign n55504 = n55503 ^ n55502;
  assign n55939 = n55774 ^ n55504;
  assign n55940 = n55939 ^ n55937;
  assign n55941 = n55938 & n55940;
  assign n55942 = n55941 ^ n52935;
  assign n55775 = n55774 ^ n55502;
  assign n55776 = ~n55504 & ~n55775;
  assign n55777 = n55776 ^ n55503;
  assign n55498 = n54574 ^ n53948;
  assign n55499 = n55498 ^ n55249;
  assign n55497 = n55405 ^ n55305;
  assign n55500 = n55499 ^ n55497;
  assign n55851 = n55777 ^ n55500;
  assign n55852 = n55851 ^ n53076;
  assign n56026 = n55942 ^ n55852;
  assign n55987 = n55916 ^ n52964;
  assign n55988 = n55890 ^ n52917;
  assign n55989 = n55988 ^ n55877;
  assign n55990 = n55884 ^ n55883;
  assign n55991 = n55887 ^ n55880;
  assign n55992 = n55990 & ~n55991;
  assign n55993 = ~n55989 & ~n55992;
  assign n55994 = n55893 ^ n52912;
  assign n55995 = n55994 ^ n55875;
  assign n55996 = ~n55993 & ~n55995;
  assign n55997 = n55898 ^ n52906;
  assign n55998 = ~n55996 & n55997;
  assign n55999 = n55901 ^ n52899;
  assign n56000 = n55999 ^ n55872;
  assign n56001 = ~n55998 & n56000;
  assign n56002 = n55904 ^ n55871;
  assign n56003 = n56001 & ~n56002;
  assign n56004 = n55907 ^ n52329;
  assign n56005 = n56004 ^ n55868;
  assign n56006 = n56003 & n56005;
  assign n56007 = n55910 ^ n55867;
  assign n56008 = ~n56006 & n56007;
  assign n56009 = n55987 & n56008;
  assign n56010 = n55919 ^ n55865;
  assign n56011 = n56009 & ~n56010;
  assign n56012 = n55922 ^ n52955;
  assign n56013 = n56012 ^ n55862;
  assign n56014 = n56011 & ~n56013;
  assign n56015 = n55925 ^ n55861;
  assign n56016 = n56014 & n56015;
  assign n56017 = n55928 ^ n55858;
  assign n56018 = ~n56016 & n56017;
  assign n56019 = n55931 ^ n55856;
  assign n56020 = n56018 & n56019;
  assign n56021 = n55934 ^ n55854;
  assign n56022 = ~n56020 & n56021;
  assign n56023 = n55939 ^ n52935;
  assign n56024 = n56023 ^ n55937;
  assign n56025 = ~n56022 & n56024;
  assign n56232 = n56026 ^ n56025;
  assign n56095 = n56024 ^ n56022;
  assign n56092 = n54164 ^ n45076;
  assign n56093 = n56092 ^ n50432;
  assign n56094 = n56093 ^ n46242;
  assign n56096 = n56095 ^ n56094;
  assign n56098 = n54151 ^ n46120;
  assign n56099 = n56098 ^ n50437;
  assign n56100 = n56099 ^ n45081;
  assign n56097 = n56021 ^ n56020;
  assign n56101 = n56100 ^ n56097;
  assign n56105 = n56019 ^ n56018;
  assign n56102 = n46124 ^ n2264;
  assign n56103 = n56102 ^ n50442;
  assign n56104 = n56103 ^ n45086;
  assign n56106 = n56105 ^ n56104;
  assign n56108 = n53696 ^ n46130;
  assign n56109 = n56108 ^ n50447;
  assign n56110 = n56109 ^ n45091;
  assign n56107 = n56017 ^ n56016;
  assign n56111 = n56110 ^ n56107;
  assign n56212 = n56015 ^ n56014;
  assign n56113 = n53701 ^ n46137;
  assign n56114 = n56113 ^ n50542;
  assign n56115 = n56114 ^ n44743;
  assign n56112 = n56013 ^ n56011;
  assign n56116 = n56115 ^ n56112;
  assign n56118 = n53705 ^ n46142;
  assign n56119 = n56118 ^ n50457;
  assign n56120 = n56119 ^ n44645;
  assign n56117 = n56010 ^ n56009;
  assign n56121 = n56120 ^ n56117;
  assign n56125 = n56008 ^ n55987;
  assign n56122 = n53711 ^ n46146;
  assign n56123 = n56122 ^ n50531;
  assign n56124 = n56123 ^ n44719;
  assign n56126 = n56125 ^ n56124;
  assign n56128 = n53716 ^ n46151;
  assign n56129 = n56128 ^ n50462;
  assign n56130 = n56129 ^ n44650;
  assign n56127 = n56007 ^ n56006;
  assign n56131 = n56130 ^ n56127;
  assign n56133 = n53720 ^ n46156;
  assign n56134 = n56133 ^ n50518;
  assign n56135 = n56134 ^ n44708;
  assign n56132 = n56005 ^ n56003;
  assign n56136 = n56135 ^ n56132;
  assign n56138 = n53725 ^ n46162;
  assign n56139 = n56138 ^ n50467;
  assign n56140 = n56139 ^ n44654;
  assign n56137 = n56002 ^ n56001;
  assign n56141 = n56140 ^ n56137;
  assign n56143 = n53768 ^ n50507;
  assign n56144 = n56143 ^ n46166;
  assign n56145 = n56144 ^ n44697;
  assign n56142 = n56000 ^ n55998;
  assign n56146 = n56145 ^ n56142;
  assign n56148 = n53758 ^ n46201;
  assign n56149 = n56148 ^ n50499;
  assign n56150 = n56149 ^ n44660;
  assign n56147 = n55997 ^ n55996;
  assign n56151 = n56150 ^ n56147;
  assign n56153 = n53750 ^ n46193;
  assign n56154 = n56153 ^ n50472;
  assign n56155 = n56154 ^ n44665;
  assign n56152 = n55995 ^ n55993;
  assign n56156 = n56155 ^ n56152;
  assign n56177 = n55992 ^ n55989;
  assign n56169 = n53735 ^ n46181;
  assign n56170 = n56169 ^ n50481;
  assign n56171 = n56170 ^ n44679;
  assign n56162 = n53730 ^ n46176;
  assign n56163 = n56162 ^ n50484;
  assign n56164 = n56163 ^ n44674;
  assign n56157 = n54246 ^ n46613;
  assign n56158 = n56157 ^ n50864;
  assign n56159 = n56158 ^ n45247;
  assign n56160 = n55881 ^ n52988;
  assign n56161 = n56159 & ~n56160;
  assign n56165 = n56164 ^ n56161;
  assign n56166 = n56161 ^ n55990;
  assign n56167 = n56165 & ~n56166;
  assign n56168 = n56167 ^ n56164;
  assign n56172 = n56171 ^ n56168;
  assign n56173 = n55991 ^ n55990;
  assign n56174 = n56173 ^ n56168;
  assign n56175 = n56172 & ~n56174;
  assign n56176 = n56175 ^ n56171;
  assign n56178 = n56177 ^ n56176;
  assign n56179 = n53742 ^ n46172;
  assign n56180 = n56179 ^ n50477;
  assign n56181 = n56180 ^ n44669;
  assign n56182 = n56181 ^ n56177;
  assign n56183 = ~n56178 & n56182;
  assign n56184 = n56183 ^ n56181;
  assign n56185 = n56184 ^ n56152;
  assign n56186 = ~n56156 & n56185;
  assign n56187 = n56186 ^ n56155;
  assign n56188 = n56187 ^ n56147;
  assign n56189 = ~n56151 & n56188;
  assign n56190 = n56189 ^ n56150;
  assign n56191 = n56190 ^ n56142;
  assign n56192 = n56146 & ~n56191;
  assign n56193 = n56192 ^ n56145;
  assign n56194 = n56193 ^ n56137;
  assign n56195 = n56141 & ~n56194;
  assign n56196 = n56195 ^ n56140;
  assign n56197 = n56196 ^ n56132;
  assign n56198 = ~n56136 & n56197;
  assign n56199 = n56198 ^ n56135;
  assign n56200 = n56199 ^ n56127;
  assign n56201 = ~n56131 & n56200;
  assign n56202 = n56201 ^ n56130;
  assign n56203 = n56202 ^ n56124;
  assign n56204 = n56126 & ~n56203;
  assign n56205 = n56204 ^ n56125;
  assign n56206 = n56205 ^ n56117;
  assign n56207 = ~n56121 & n56206;
  assign n56208 = n56207 ^ n56120;
  assign n56209 = n56208 ^ n56112;
  assign n56210 = ~n56116 & n56209;
  assign n56211 = n56210 ^ n56115;
  assign n56213 = n56212 ^ n56211;
  assign n56214 = n53794 ^ n2148;
  assign n56215 = n56214 ^ n50452;
  assign n56216 = n56215 ^ n45096;
  assign n56217 = n56216 ^ n56212;
  assign n56218 = ~n56213 & n56217;
  assign n56219 = n56218 ^ n56216;
  assign n56220 = n56219 ^ n56107;
  assign n56221 = n56111 & ~n56220;
  assign n56222 = n56221 ^ n56110;
  assign n56223 = n56222 ^ n56104;
  assign n56224 = ~n56106 & ~n56223;
  assign n56225 = n56224 ^ n56105;
  assign n56226 = n56225 ^ n56097;
  assign n56227 = ~n56101 & ~n56226;
  assign n56228 = n56227 ^ n56100;
  assign n56229 = n56228 ^ n56094;
  assign n56230 = n56096 & ~n56229;
  assign n56231 = n56230 ^ n56095;
  assign n56233 = n56232 ^ n56231;
  assign n56312 = n56236 ^ n56233;
  assign n56313 = n56160 ^ n56159;
  assign n56314 = n56164 ^ n55990;
  assign n56315 = n56314 ^ n56161;
  assign n56316 = ~n56313 & n56315;
  assign n56317 = n56173 ^ n56171;
  assign n56318 = n56317 ^ n56168;
  assign n56319 = n56316 & n56318;
  assign n56320 = n56181 ^ n56178;
  assign n56321 = n56319 & n56320;
  assign n56322 = n56184 ^ n56155;
  assign n56323 = n56322 ^ n56152;
  assign n56324 = n56321 & ~n56323;
  assign n56325 = n56187 ^ n56151;
  assign n56326 = n56324 & ~n56325;
  assign n56327 = n56190 ^ n56146;
  assign n56328 = n56326 & n56327;
  assign n56329 = n56193 ^ n56140;
  assign n56330 = n56329 ^ n56137;
  assign n56331 = n56328 & n56330;
  assign n56332 = n56196 ^ n56136;
  assign n56333 = ~n56331 & n56332;
  assign n56334 = n56199 ^ n56131;
  assign n56335 = n56333 & n56334;
  assign n56336 = n56202 ^ n56126;
  assign n56337 = ~n56335 & n56336;
  assign n56338 = n56205 ^ n56121;
  assign n56339 = n56337 & ~n56338;
  assign n56340 = n56208 ^ n56116;
  assign n56341 = n56339 & ~n56340;
  assign n56342 = n56216 ^ n56213;
  assign n56343 = ~n56341 & ~n56342;
  assign n56344 = n56219 ^ n56111;
  assign n56345 = ~n56343 & n56344;
  assign n56346 = n56222 ^ n56106;
  assign n56347 = n56345 & ~n56346;
  assign n56348 = n56225 ^ n56101;
  assign n56349 = ~n56347 & ~n56348;
  assign n56350 = n56228 ^ n56096;
  assign n56351 = ~n56349 & n56350;
  assign n56352 = n56312 & ~n56351;
  assign n56237 = n56236 ^ n56232;
  assign n56238 = n56233 & ~n56237;
  assign n56239 = n56238 ^ n56236;
  assign n55943 = n55942 ^ n55851;
  assign n55944 = n55852 & n55943;
  assign n55945 = n55944 ^ n53076;
  assign n55778 = n55777 ^ n55497;
  assign n55779 = n55500 & n55778;
  assign n55780 = n55779 ^ n55499;
  assign n55494 = n55446 ^ n54585;
  assign n55495 = n55494 ^ n53874;
  assign n55492 = n55408 ^ n55299;
  assign n55493 = n55492 ^ n55296;
  assign n55496 = n55495 ^ n55493;
  assign n55849 = n55780 ^ n55496;
  assign n55850 = n55849 ^ n52929;
  assign n56028 = n55945 ^ n55850;
  assign n56027 = ~n56025 & n56026;
  assign n56090 = n56028 ^ n56027;
  assign n56087 = n54141 ^ n46269;
  assign n56088 = n56087 ^ n50427;
  assign n56089 = n56088 ^ n45128;
  assign n56091 = n56090 ^ n56089;
  assign n56353 = n56239 ^ n56091;
  assign n56354 = ~n56352 & ~n56353;
  assign n56240 = n56239 ^ n56089;
  assign n56241 = ~n56091 & ~n56240;
  assign n56242 = n56241 ^ n56090;
  assign n55946 = n55945 ^ n55849;
  assign n55947 = n55850 & n55946;
  assign n55948 = n55947 ^ n52929;
  assign n55786 = n55531 ^ n53869;
  assign n55787 = n55786 ^ n54599;
  assign n55784 = n55411 ^ n55295;
  assign n55781 = n55780 ^ n55493;
  assign n55782 = n55496 & n55781;
  assign n55783 = n55782 ^ n55495;
  assign n55785 = n55784 ^ n55783;
  assign n55847 = n55787 ^ n55785;
  assign n55848 = n55847 ^ n52925;
  assign n56030 = n55948 ^ n55848;
  assign n56029 = n56027 & ~n56028;
  assign n56085 = n56030 ^ n56029;
  assign n56082 = n54137 ^ n46532;
  assign n56083 = n56082 ^ n50576;
  assign n56084 = n56083 ^ n45136;
  assign n56086 = n56085 ^ n56084;
  assign n56355 = n56242 ^ n56086;
  assign n56356 = n56354 & ~n56355;
  assign n56243 = n56242 ^ n56084;
  assign n56244 = n56086 & n56243;
  assign n56245 = n56244 ^ n56085;
  assign n56078 = n54132 ^ n46545;
  assign n56079 = n56078 ^ n50422;
  assign n56080 = n56079 ^ n45071;
  assign n56357 = n56245 ^ n56080;
  assign n56031 = n56029 & n56030;
  assign n55949 = n55948 ^ n55847;
  assign n55950 = n55848 & n55949;
  assign n55951 = n55950 ^ n52925;
  assign n55788 = n55787 ^ n55784;
  assign n55789 = n55785 & n55788;
  assign n55790 = n55789 ^ n55787;
  assign n55490 = n55414 ^ n55290;
  assign n55488 = n55487 ^ n53866;
  assign n55489 = n55488 ^ n54618;
  assign n55491 = n55490 ^ n55489;
  assign n55845 = n55790 ^ n55491;
  assign n55846 = n55845 ^ n52921;
  assign n55986 = n55951 ^ n55846;
  assign n56077 = n56031 ^ n55986;
  assign n56358 = n56357 ^ n56077;
  assign n56359 = n56356 & n56358;
  assign n56251 = n54184 ^ n46528;
  assign n56252 = n56251 ^ n50417;
  assign n56253 = n56252 ^ n45066;
  assign n55952 = n55951 ^ n55845;
  assign n55953 = n55846 & n55952;
  assign n55954 = n55953 ^ n52921;
  assign n55791 = n55790 ^ n55489;
  assign n55792 = n55491 & n55791;
  assign n55793 = n55792 ^ n55490;
  assign n55484 = n55483 ^ n53967;
  assign n55485 = n55484 ^ n54863;
  assign n55481 = n55417 ^ n55284;
  assign n55482 = n55481 ^ n55281;
  assign n55486 = n55485 ^ n55482;
  assign n55843 = n55793 ^ n55486;
  assign n55844 = n55843 ^ n53095;
  assign n56033 = n55954 ^ n55844;
  assign n56032 = n55986 & ~n56031;
  assign n56249 = n56033 ^ n56032;
  assign n56081 = n56080 ^ n56077;
  assign n56246 = n56245 ^ n56077;
  assign n56247 = n56081 & ~n56246;
  assign n56248 = n56247 ^ n56080;
  assign n56250 = n56249 ^ n56248;
  assign n56360 = n56253 ^ n56250;
  assign n56361 = ~n56359 & n56360;
  assign n56259 = n54190 ^ n46522;
  assign n56260 = n56259 ^ n50590;
  assign n56261 = n56260 ^ n45150;
  assign n56034 = n56032 & n56033;
  assign n55794 = n55793 ^ n55482;
  assign n55795 = ~n55486 & n55794;
  assign n55796 = n55795 ^ n55485;
  assign n55478 = n55477 ^ n54057;
  assign n55479 = n55478 ^ n54942;
  assign n55475 = n55420 ^ n55279;
  assign n55476 = n55475 ^ n55276;
  assign n55480 = n55479 ^ n55476;
  assign n55958 = n55796 ^ n55480;
  assign n55955 = n55954 ^ n55843;
  assign n55956 = ~n55844 & ~n55955;
  assign n55957 = n55956 ^ n53095;
  assign n55959 = n55958 ^ n55957;
  assign n55985 = n55959 ^ n53234;
  assign n56257 = n56034 ^ n55985;
  assign n56254 = n56253 ^ n56249;
  assign n56255 = n56250 & ~n56254;
  assign n56256 = n56255 ^ n56253;
  assign n56258 = n56257 ^ n56256;
  assign n56362 = n56261 ^ n56258;
  assign n56363 = ~n56361 & ~n56362;
  assign n56262 = n56261 ^ n56257;
  assign n56263 = n56258 & ~n56262;
  assign n56264 = n56263 ^ n56261;
  assign n56073 = n54127 ^ n46518;
  assign n56074 = n56073 ^ n50412;
  assign n56075 = n56074 ^ n45061;
  assign n55960 = n55958 ^ n53234;
  assign n55961 = ~n55959 & ~n55960;
  assign n55962 = n55961 ^ n53234;
  assign n55802 = n55619 ^ n54234;
  assign n55803 = n55802 ^ n54968;
  assign n55800 = n55423 ^ n55275;
  assign n55797 = n55796 ^ n55476;
  assign n55798 = n55480 & n55797;
  assign n55799 = n55798 ^ n55479;
  assign n55801 = n55800 ^ n55799;
  assign n55841 = n55803 ^ n55801;
  assign n55842 = n55841 ^ n53517;
  assign n56036 = n55962 ^ n55842;
  assign n56035 = n55985 & ~n56034;
  assign n56072 = n56036 ^ n56035;
  assign n56076 = n56075 ^ n56072;
  assign n56364 = n56264 ^ n56076;
  assign n56365 = ~n56363 & n56364;
  assign n56265 = n56264 ^ n56072;
  assign n56266 = ~n56076 & n56265;
  assign n56267 = n56266 ^ n56075;
  assign n56068 = n54203 ^ n46513;
  assign n56069 = n56068 ^ n50407;
  assign n56070 = n56069 ^ n45161;
  assign n56366 = n56267 ^ n56070;
  assign n55804 = n55803 ^ n55800;
  assign n55805 = ~n55801 & n55804;
  assign n55806 = n55805 ^ n55803;
  assign n55472 = n55426 ^ n55269;
  assign n55473 = n55472 ^ n55266;
  assign n55469 = n54265 ^ n53544;
  assign n55471 = n55470 ^ n55469;
  assign n55474 = n55473 ^ n55471;
  assign n55966 = n55806 ^ n55474;
  assign n55963 = n55962 ^ n55841;
  assign n55964 = ~n55842 & ~n55963;
  assign n55965 = n55964 ^ n53517;
  assign n55967 = n55966 ^ n55965;
  assign n56038 = n55967 ^ n52741;
  assign n56037 = n56035 & ~n56036;
  assign n56067 = n56038 ^ n56037;
  assign n56367 = n56366 ^ n56067;
  assign n56368 = n56365 & ~n56367;
  assign n56071 = n56070 ^ n56067;
  assign n56268 = n56267 ^ n56067;
  assign n56269 = n56071 & ~n56268;
  assign n56270 = n56269 ^ n56070;
  assign n56063 = n54211 ^ n1022;
  assign n56064 = n56063 ^ n50402;
  assign n56065 = n56064 ^ n45056;
  assign n56369 = n56270 ^ n56065;
  assign n55968 = n55966 ^ n52741;
  assign n55969 = ~n55967 & n55968;
  assign n55970 = n55969 ^ n52741;
  assign n55813 = n55662 ^ n53549;
  assign n55814 = n55813 ^ n54258;
  assign n55810 = n55429 ^ n55264;
  assign n55811 = n55810 ^ n55261;
  assign n55807 = n55806 ^ n55471;
  assign n55808 = ~n55474 & ~n55807;
  assign n55809 = n55808 ^ n55473;
  assign n55812 = n55811 ^ n55809;
  assign n55839 = n55814 ^ n55812;
  assign n55840 = n55839 ^ n52735;
  assign n56040 = n55970 ^ n55840;
  assign n56039 = ~n56037 & n56038;
  assign n56062 = n56040 ^ n56039;
  assign n56370 = n56369 ^ n56062;
  assign n56371 = n56368 & n56370;
  assign n56066 = n56065 ^ n56062;
  assign n56271 = n56270 ^ n56062;
  assign n56272 = ~n56066 & n56271;
  assign n56273 = n56272 ^ n56065;
  assign n55971 = n55970 ^ n55839;
  assign n55972 = ~n55840 & ~n55971;
  assign n55973 = n55972 ^ n52735;
  assign n55815 = n55814 ^ n55811;
  assign n55816 = n55812 & n55815;
  assign n55817 = n55816 ^ n55814;
  assign n55466 = n54273 ^ n53538;
  assign n55467 = n55466 ^ n54984;
  assign n55465 = n55432 ^ n55260;
  assign n55468 = n55467 ^ n55465;
  assign n55837 = n55817 ^ n55468;
  assign n55838 = n55837 ^ n52780;
  assign n56042 = n55973 ^ n55838;
  assign n56041 = ~n56039 & n56040;
  assign n56060 = n56042 ^ n56041;
  assign n56057 = n54122 ^ n46506;
  assign n56058 = n56057 ^ n50621;
  assign n56059 = n56058 ^ n1188;
  assign n56061 = n56060 ^ n56059;
  assign n56372 = n56273 ^ n56061;
  assign n56373 = ~n56371 & n56372;
  assign n56274 = n56273 ^ n56059;
  assign n56275 = n56061 & ~n56274;
  assign n56276 = n56275 ^ n56060;
  assign n56053 = n54117 ^ n46501;
  assign n56054 = n56053 ^ n1199;
  assign n56055 = n56054 ^ n45175;
  assign n55974 = n55973 ^ n55837;
  assign n55975 = ~n55838 & n55974;
  assign n55976 = n55975 ^ n52780;
  assign n55818 = n55817 ^ n55465;
  assign n55819 = ~n55468 & n55818;
  assign n55820 = n55819 ^ n55467;
  assign n55462 = n54254 ^ n53535;
  assign n55463 = n55462 ^ n54989;
  assign n55461 = n55435 ^ n55255;
  assign n55464 = n55463 ^ n55461;
  assign n55835 = n55820 ^ n55464;
  assign n55836 = n55835 ^ n52811;
  assign n56044 = n55976 ^ n55836;
  assign n56043 = ~n56041 & n56042;
  assign n56052 = n56044 ^ n56043;
  assign n56056 = n56055 ^ n56052;
  assign n56374 = n56276 ^ n56056;
  assign n56375 = n56373 & n56374;
  assign n56282 = n54112 ^ n46495;
  assign n56283 = n56282 ^ n50679;
  assign n56284 = n56283 ^ n1361;
  assign n56045 = ~n56043 & ~n56044;
  assign n55977 = n55976 ^ n55835;
  assign n55978 = ~n55836 & ~n55977;
  assign n55979 = n55978 ^ n52811;
  assign n55821 = n55820 ^ n55461;
  assign n55822 = n55464 & ~n55821;
  assign n55823 = n55822 ^ n55463;
  assign n55459 = n55458 ^ n55438;
  assign n54870 = n54869 ^ n54250;
  assign n54871 = n54870 ^ n53528;
  assign n55460 = n55459 ^ n54871;
  assign n55833 = n55823 ^ n55460;
  assign n55834 = n55833 ^ n52883;
  assign n55984 = n55979 ^ n55834;
  assign n56280 = n56045 ^ n55984;
  assign n56277 = n56276 ^ n56052;
  assign n56278 = n56056 & ~n56277;
  assign n56279 = n56278 ^ n56055;
  assign n56281 = n56280 ^ n56279;
  assign n56376 = n56284 ^ n56281;
  assign n56377 = ~n56375 & n56376;
  assign n56285 = n56284 ^ n56280;
  assign n56286 = n56281 & ~n56285;
  assign n56287 = n56286 ^ n56284;
  assign n56048 = n54106 ^ n46491;
  assign n56049 = n56048 ^ n50722;
  assign n56050 = n56049 ^ n44800;
  assign n56378 = n56287 ^ n56050;
  assign n56046 = ~n55984 & n56045;
  assign n55980 = n55979 ^ n55833;
  assign n55981 = n55834 & ~n55980;
  assign n55982 = n55981 ^ n52883;
  assign n55828 = n55002 ^ n52916;
  assign n55829 = n55828 ^ n53862;
  assign n55827 = n55546 ^ n55543;
  assign n55830 = n55829 ^ n55827;
  assign n55824 = n55823 ^ n54871;
  assign n55825 = ~n55460 & n55824;
  assign n55826 = n55825 ^ n55459;
  assign n55831 = n55830 ^ n55826;
  assign n55832 = n55831 ^ n52995;
  assign n55983 = n55982 ^ n55832;
  assign n56047 = n56046 ^ n55983;
  assign n56379 = n56378 ^ n56047;
  assign n56380 = n56377 & n56379;
  assign n56307 = n54102 ^ n46594;
  assign n56308 = n56307 ^ n50743;
  assign n56309 = n56308 ^ n44797;
  assign n56300 = n54977 ^ n53858;
  assign n56301 = n56300 ^ n52910;
  assign n56299 = n55567 ^ n55564;
  assign n56302 = n56301 ^ n56299;
  assign n56296 = n55829 ^ n55826;
  assign n56297 = ~n55830 & ~n56296;
  assign n56298 = n56297 ^ n55826;
  assign n56303 = n56302 ^ n56298;
  assign n56292 = n55982 ^ n52995;
  assign n56293 = n55982 ^ n55831;
  assign n56294 = n56292 & n56293;
  assign n56295 = n56294 ^ n52995;
  assign n56304 = n56303 ^ n56295;
  assign n56305 = n56304 ^ n52993;
  assign n56291 = ~n55983 & ~n56046;
  assign n56306 = n56305 ^ n56291;
  assign n56310 = n56309 ^ n56306;
  assign n56051 = n56050 ^ n56047;
  assign n56288 = n56287 ^ n56047;
  assign n56289 = ~n56051 & n56288;
  assign n56290 = n56289 ^ n56050;
  assign n56311 = n56310 ^ n56290;
  assign n56381 = n56380 ^ n56311;
  assign n56382 = n56379 ^ n56377;
  assign n56383 = n56376 ^ n56375;
  assign n56384 = n56374 ^ n56373;
  assign n56385 = n56372 ^ n56371;
  assign n56386 = n56370 ^ n56368;
  assign n56387 = n56367 ^ n56365;
  assign n56388 = n56364 ^ n56363;
  assign n56389 = n56362 ^ n56361;
  assign n56390 = n56360 ^ n56359;
  assign n56391 = n56358 ^ n56356;
  assign n56392 = n56355 ^ n56354;
  assign n56393 = n56353 ^ n56352;
  assign n56394 = n56351 ^ n56312;
  assign n56395 = n56350 ^ n56349;
  assign n56396 = n56348 ^ n56347;
  assign n56397 = n56346 ^ n56345;
  assign n56398 = n56344 ^ n56343;
  assign n56399 = n56342 ^ n56341;
  assign n56400 = n56340 ^ n56339;
  assign n56401 = n56338 ^ n56337;
  assign n56402 = n56336 ^ n56335;
  assign n56403 = n56334 ^ n56333;
  assign n56404 = n56332 ^ n56331;
  assign n56405 = n56330 ^ n56328;
  assign n56406 = n56327 ^ n56326;
  assign n56407 = n56325 ^ n56324;
  assign n56408 = n56323 ^ n56321;
  assign n56409 = n56320 ^ n56319;
  assign n56410 = n56318 ^ n56316;
  assign n56411 = n56315 ^ n56313;
  assign n56412 = n55706 & ~n55714;
  assign n56413 = ~n55721 & n56412;
  assign n56414 = ~n55728 & ~n56413;
  assign n56415 = n55518 & ~n56414;
  assign n56416 = ~n55741 & n56415;
  assign n56417 = ~n55745 & n56416;
  assign n56418 = ~n55752 & ~n56417;
  assign n56419 = ~n55514 & n56418;
  assign n56420 = n55510 & n56419;
  assign n56421 = ~n55765 & ~n56420;
  assign n56422 = ~n55505 & ~n56421;
  assign n56423 = ~n55503 & ~n56422;
  assign n56424 = ~n55497 & ~n56423;
  assign n56425 = ~n55493 & ~n56424;
  assign n56426 = ~n55784 & ~n56425;
  assign n56427 = n55490 & n56426;
  assign n56428 = n55482 & ~n56427;
  assign n56429 = ~n55476 & ~n56428;
  assign n56430 = ~n55800 & n56429;
  assign n56431 = ~n55473 & ~n56430;
  assign n56432 = n55811 & n56431;
  assign n56433 = n55465 & ~n56432;
  assign n56434 = ~n55461 & n56433;
  assign n56435 = ~n55459 & n56434;
  assign n56436 = n55827 & n56435;
  assign n56437 = n56299 & n56436;
  assign n56438 = n55680 & n56437;
  assign n56439 = n55685 & ~n56438;
  assign n56440 = n55689 & ~n56439;
  assign n56441 = n55696 & n56440;
  assign n56442 = n56441 ^ n55675;
  assign n56443 = n56440 ^ n55696;
  assign n56444 = n56439 ^ n55689;
  assign n56445 = n56438 ^ n55685;
  assign n56446 = n56437 ^ n55680;
  assign n56447 = n56436 ^ n56299;
  assign n56448 = n56435 ^ n55827;
  assign n56449 = n56434 ^ n55459;
  assign n56450 = n56433 ^ n55461;
  assign n56451 = n56432 ^ n55465;
  assign n56452 = n56431 ^ n55811;
  assign n56453 = n56430 ^ n55473;
  assign n56454 = n56429 ^ n55800;
  assign n56455 = n56428 ^ n55476;
  assign n56456 = n56427 ^ n55482;
  assign n56457 = n56426 ^ n55490;
  assign n56458 = n56425 ^ n55784;
  assign n56459 = n56424 ^ n55493;
  assign n56460 = n56423 ^ n55497;
  assign n56461 = n56422 ^ n55503;
  assign n56462 = n56421 ^ n55505;
  assign n56463 = n56420 ^ n55765;
  assign n56464 = n56419 ^ n55510;
  assign n56465 = n56418 ^ n55514;
  assign n56466 = n56417 ^ n55752;
  assign n56467 = n56416 ^ n55745;
  assign n56468 = n56415 ^ n55741;
  assign n56469 = n56414 ^ n55518;
  assign n56470 = n56413 ^ n55728;
  assign n56471 = n56412 ^ n55721;
  assign n56472 = n55714 ^ n55706;
  assign n56473 = n54909 & ~n54914;
  assign n56474 = ~n54905 & n56473;
  assign n56475 = n54901 & n56474;
  assign n56476 = ~n54899 & n56475;
  assign n56477 = n54892 & n56476;
  assign n56478 = n54890 & n56477;
  assign n56479 = ~n54886 & ~n56478;
  assign n56480 = ~n54879 & n56479;
  assign n56481 = ~n54875 & ~n56480;
  assign n56482 = ~n55048 & n56481;
  assign n56483 = n55057 & n56482;
  assign n56484 = ~n55168 & ~n56483;
  assign n56485 = ~n55221 & ~n56484;
  assign n56486 = n55233 & n56485;
  assign n56487 = ~n55249 & ~n56486;
  assign n56488 = n55446 & ~n56487;
  assign n56489 = n55531 & ~n56488;
  assign n56490 = ~n55487 & ~n56489;
  assign n56491 = n55483 & n56490;
  assign n56492 = n55477 & n56491;
  assign n56493 = n55619 & ~n56492;
  assign n56494 = n55470 & ~n56493;
  assign n56495 = n55662 & ~n56494;
  assign n56496 = n54984 & n56495;
  assign n56497 = n54989 & n56496;
  assign n56498 = n54869 & ~n56497;
  assign n56499 = ~n55002 & n56498;
  assign n56500 = n54977 & ~n56499;
  assign n56501 = ~n54928 & n56500;
  assign n56502 = n56501 ^ n54924;
  assign n56503 = n56500 ^ n54928;
  assign n56504 = n56499 ^ n54977;
  assign n56505 = n56498 ^ n55002;
  assign n56506 = n56497 ^ n54869;
  assign n56507 = n56496 ^ n54989;
  assign n56508 = n56495 ^ n54984;
  assign n56509 = n56494 ^ n55662;
  assign n56510 = n56493 ^ n55470;
  assign n56511 = n56492 ^ n55619;
  assign n56512 = n56491 ^ n55477;
  assign n56513 = n56490 ^ n55483;
  assign n56514 = n56489 ^ n55487;
  assign n56515 = n56488 ^ n55531;
  assign n56516 = n56487 ^ n55446;
  assign n56517 = n56486 ^ n55249;
  assign n56518 = n56485 ^ n55233;
  assign n56519 = n56484 ^ n55221;
  assign n56520 = n56483 ^ n55168;
  assign n56521 = n56482 ^ n55057;
  assign n56522 = n56481 ^ n55048;
  assign n56523 = n56480 ^ n54875;
  assign n56524 = n56479 ^ n54879;
  assign n56525 = n56478 ^ n54886;
  assign n56526 = n56477 ^ n54890;
  assign n56527 = n56476 ^ n54892;
  assign n56528 = n56475 ^ n54899;
  assign n56529 = n56474 ^ n54901;
  assign n56530 = n56473 ^ n54905;
  assign n56531 = n54914 ^ n54909;
  assign n56532 = ~n53845 & n53848;
  assign n56533 = n53841 & ~n56532;
  assign n56534 = ~n54301 & ~n56533;
  assign n56535 = ~n54308 & n56534;
  assign n56536 = ~n54316 & n56535;
  assign n56537 = ~n53832 & ~n56536;
  assign n56538 = ~n53826 & n56537;
  assign n56539 = n53824 & n56538;
  assign n56540 = ~n54332 & ~n56539;
  assign n56541 = ~n53819 & ~n56540;
  assign n56542 = ~n53817 & ~n56541;
  assign n56543 = ~n54354 & ~n56542;
  assign n56544 = n54469 & ~n56543;
  assign n56545 = ~n54480 & ~n56544;
  assign n56546 = n54489 & n56545;
  assign n56547 = ~n54552 & ~n56546;
  assign n56548 = n54574 & ~n56547;
  assign n56549 = ~n54585 & n56548;
  assign n56550 = n54599 & ~n56549;
  assign n56551 = n54618 & n56550;
  assign n56552 = ~n54863 & ~n56551;
  assign n56553 = n54942 & n56552;
  assign n56554 = ~n54968 & n56553;
  assign n56555 = ~n54265 & n56554;
  assign n56556 = ~n54258 & n56555;
  assign n56557 = ~n54273 & n56556;
  assign n56558 = n54254 & ~n56557;
  assign n56559 = n54250 & ~n56558;
  assign n56560 = n53862 & n56559;
  assign n56561 = n56560 ^ n53858;
  assign n56562 = n56559 ^ n53862;
  assign n56563 = n56558 ^ n54250;
  assign n56564 = n56557 ^ n54254;
  assign n56565 = n56556 ^ n54273;
  assign n56566 = n56555 ^ n54258;
  assign n56567 = n56554 ^ n54265;
  assign n56568 = n56553 ^ n54968;
  assign n56569 = n56552 ^ n54942;
  assign n56570 = n56551 ^ n54863;
  assign n56571 = n56550 ^ n54618;
  assign n56572 = n56549 ^ n54599;
  assign n56573 = n56548 ^ n54585;
  assign n56574 = n56547 ^ n54574;
  assign n56575 = n56546 ^ n54552;
  assign n56576 = n56545 ^ n54489;
  assign n56577 = n56544 ^ n54480;
  assign n56578 = n56543 ^ n54469;
  assign n56579 = n56542 ^ n54354;
  assign n56580 = n56541 ^ n53817;
  assign n56581 = n56540 ^ n53819;
  assign n56582 = n56539 ^ n54332;
  assign n56583 = n56538 ^ n53824;
  assign n56584 = n56537 ^ n53826;
  assign n56585 = n56536 ^ n53832;
  assign n56586 = n56535 ^ n54316;
  assign n56587 = n56534 ^ n54308;
  assign n56588 = n56533 ^ n54301;
  assign n56589 = n56532 ^ n53841;
  assign n56590 = n53848 ^ n53845;
  assign n56591 = ~n53639 & ~n53672;
  assign n56592 = n53686 & n56591;
  assign n56593 = ~n53809 & n56592;
  assign n56594 = ~n53838 & n56593;
  assign n56595 = n53901 & ~n56594;
  assign n56596 = n53896 & n56595;
  assign n56597 = n53893 & n56596;
  assign n56598 = ~n53833 & n56597;
  assign n56599 = n53828 & ~n56598;
  assign n56600 = ~n53821 & n56599;
  assign n56601 = n53880 & n56600;
  assign n56602 = n53936 & ~n56601;
  assign n56603 = n53940 & ~n56602;
  assign n56604 = ~n53948 & ~n56603;
  assign n56605 = ~n53874 & n56604;
  assign n56606 = n53869 & ~n56605;
  assign n56607 = n53866 & ~n56606;
  assign n56608 = n53967 & ~n56607;
  assign n56609 = n54057 & n56608;
  assign n56610 = n54234 & n56609;
  assign n56611 = ~n53544 & n56610;
  assign n56612 = ~n53549 & ~n56611;
  assign n56613 = ~n53538 & n56612;
  assign n56614 = ~n53535 & n56613;
  assign n56615 = n53528 & n56614;
  assign n56616 = n52916 & ~n56615;
  assign n56617 = n56616 ^ n52910;
  assign n56618 = n56615 ^ n52916;
  assign n56619 = n56614 ^ n53528;
  assign n56620 = n56613 ^ n53535;
  assign n56621 = n56612 ^ n53538;
  assign n56622 = n56611 ^ n53549;
  assign n56623 = n56610 ^ n53544;
  assign n56624 = n56609 ^ n54234;
  assign n56625 = n56608 ^ n54057;
  assign n56626 = n56607 ^ n53967;
  assign n56627 = n56606 ^ n53866;
  assign n56628 = n56605 ^ n53869;
  assign n56629 = n56604 ^ n53874;
  assign n56630 = n56603 ^ n53948;
  assign n56631 = n56602 ^ n53940;
  assign n56632 = n56601 ^ n53936;
  assign n56633 = n56600 ^ n53880;
  assign n56634 = n56599 ^ n53821;
  assign n56635 = n56598 ^ n53828;
  assign n56636 = n56597 ^ n53833;
  assign n56637 = n56596 ^ n53893;
  assign n56638 = n56595 ^ n53896;
  assign n56639 = n56594 ^ n53901;
  assign n56640 = n56593 ^ n53838;
  assign n56641 = n56592 ^ n53809;
  assign n56642 = n56591 ^ n53686;
  assign n56643 = n53672 ^ n53639;
  assign y0 = ~n56381;
  assign y1 = ~n56382;
  assign y2 = n56383;
  assign y3 = n56384;
  assign y4 = ~n56385;
  assign y5 = ~n56386;
  assign y6 = n56387;
  assign y7 = n56388;
  assign y8 = n56389;
  assign y9 = n56390;
  assign y10 = n56391;
  assign y11 = ~n56392;
  assign y12 = n56393;
  assign y13 = n56394;
  assign y14 = ~n56395;
  assign y15 = ~n56396;
  assign y16 = ~n56397;
  assign y17 = ~n56398;
  assign y18 = ~n56399;
  assign y19 = ~n56400;
  assign y20 = ~n56401;
  assign y21 = ~n56402;
  assign y22 = ~n56403;
  assign y23 = n56404;
  assign y24 = n56405;
  assign y25 = n56406;
  assign y26 = ~n56407;
  assign y27 = ~n56408;
  assign y28 = n56409;
  assign y29 = n56410;
  assign y30 = ~n56411;
  assign y31 = n56313;
  assign y32 = ~n56442;
  assign y33 = ~n56443;
  assign y34 = n56444;
  assign y35 = ~n56445;
  assign y36 = ~n56446;
  assign y37 = ~n56447;
  assign y38 = ~n56448;
  assign y39 = n56449;
  assign y40 = n56450;
  assign y41 = n56451;
  assign y42 = n56452;
  assign y43 = n56453;
  assign y44 = n56454;
  assign y45 = ~n56455;
  assign y46 = ~n56456;
  assign y47 = ~n56457;
  assign y48 = ~n56458;
  assign y49 = n56459;
  assign y50 = ~n56460;
  assign y51 = n56461;
  assign y52 = ~n56462;
  assign y53 = n56463;
  assign y54 = ~n56464;
  assign y55 = n56465;
  assign y56 = ~n56466;
  assign y57 = ~n56467;
  assign y58 = ~n56468;
  assign y59 = ~n56469;
  assign y60 = ~n56470;
  assign y61 = ~n56471;
  assign y62 = ~n56472;
  assign y63 = ~n55706;
  assign y64 = ~n56502;
  assign y65 = ~n56503;
  assign y66 = ~n56504;
  assign y67 = n56505;
  assign y68 = n56506;
  assign y69 = n56507;
  assign y70 = n56508;
  assign y71 = ~n56509;
  assign y72 = n56510;
  assign y73 = ~n56511;
  assign y74 = ~n56512;
  assign y75 = ~n56513;
  assign y76 = ~n56514;
  assign y77 = ~n56515;
  assign y78 = n56516;
  assign y79 = n56517;
  assign y80 = ~n56518;
  assign y81 = ~n56519;
  assign y82 = n56520;
  assign y83 = ~n56521;
  assign y84 = n56522;
  assign y85 = ~n56523;
  assign y86 = ~n56524;
  assign y87 = n56525;
  assign y88 = ~n56526;
  assign y89 = ~n56527;
  assign y90 = n56528;
  assign y91 = ~n56529;
  assign y92 = n56530;
  assign y93 = n56531;
  assign y94 = ~n54914;
  assign y95 = ~n54919;
  assign y96 = n56561;
  assign y97 = n56562;
  assign y98 = ~n56563;
  assign y99 = n56564;
  assign y100 = ~n56565;
  assign y101 = ~n56566;
  assign y102 = ~n56567;
  assign y103 = ~n56568;
  assign y104 = n56569;
  assign y105 = n56570;
  assign y106 = ~n56571;
  assign y107 = n56572;
  assign y108 = ~n56573;
  assign y109 = ~n56574;
  assign y110 = ~n56575;
  assign y111 = n56576;
  assign y112 = n56577;
  assign y113 = n56578;
  assign y114 = n56579;
  assign y115 = ~n56580;
  assign y116 = n56581;
  assign y117 = ~n56582;
  assign y118 = n56583;
  assign y119 = ~n56584;
  assign y120 = n56585;
  assign y121 = n56586;
  assign y122 = n56587;
  assign y123 = ~n56588;
  assign y124 = ~n56589;
  assign y125 = n56590;
  assign y126 = n53848;
  assign y127 = n53853;
  assign y128 = ~n56617;
  assign y129 = n56618;
  assign y130 = n56619;
  assign y131 = ~n56620;
  assign y132 = ~n56621;
  assign y133 = n56622;
  assign y134 = n56623;
  assign y135 = ~n56624;
  assign y136 = ~n56625;
  assign y137 = n56626;
  assign y138 = ~n56627;
  assign y139 = n56628;
  assign y140 = ~n56629;
  assign y141 = n56630;
  assign y142 = n56631;
  assign y143 = ~n56632;
  assign y144 = ~n56633;
  assign y145 = n56634;
  assign y146 = n56635;
  assign y147 = ~n56636;
  assign y148 = n56637;
  assign y149 = n56638;
  assign y150 = ~n56639;
  assign y151 = n56640;
  assign y152 = n56641;
  assign y153 = ~n56642;
  assign y154 = ~n56643;
  assign y155 = ~n53639;
  assign y156 = ~n53577;
  assign y157 = ~n52892;
  assign y158 = n52898;
  assign y159 = ~n52904;
endmodule
