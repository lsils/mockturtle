module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 ;
  wire n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 ;
  assign n36 = x1 & x11 ;
  assign n37 = ( x0 & x10 ) | ( x0 & n36 ) | ( x10 & n36 ) ;
  assign n38 = ~x0 & n37 ;
  assign n39 = ( x1 & x9 ) | ( x1 & ~n38 ) | ( x9 & ~n38 ) ;
  assign n40 = x3 & n39 ;
  assign n41 = ( x3 & n38 ) | ( x3 & ~n40 ) | ( n38 & ~n40 ) ;
  assign n27 = ~x17 & x18 ;
  assign n42 = x16 & ~n27 ;
  assign n43 = ( x14 & ~n41 ) | ( x14 & n42 ) | ( ~n41 & n42 ) ;
  assign n44 = n41 & n43 ;
  assign n45 = ~x0 & x2 ;
  assign n46 = x1 & n45 ;
  assign n47 = x3 & n46 ;
  assign n48 = ( x5 & x18 ) | ( x5 & n47 ) | ( x18 & n47 ) ;
  assign n49 = ~x18 & n48 ;
  assign n50 = ( x2 & x5 ) | ( x2 & ~n49 ) | ( x5 & ~n49 ) ;
  assign n51 = n44 & n50 ;
  assign n52 = ( n44 & n49 ) | ( n44 & ~n51 ) | ( n49 & ~n51 ) ;
  assign n79 = ~x15 & n52 ;
  assign n53 = x1 & x3 ;
  assign n54 = ( x0 & x2 ) | ( x0 & n53 ) | ( x2 & n53 ) ;
  assign n55 = ~x0 & n54 ;
  assign n56 = x17 | x18 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = ( x5 & x15 ) | ( x5 & n57 ) | ( x15 & n57 ) ;
  assign n59 = ~x15 & n58 ;
  assign n60 = x14 & x16 ;
  assign n69 = x5 | x18 ;
  assign n70 = x9 | n69 ;
  assign n71 = ~x2 & x3 ;
  assign n72 = ( x1 & ~n70 ) | ( x1 & n71 ) | ( ~n70 & n71 ) ;
  assign n73 = ~x1 & n72 ;
  assign n61 = x10 & ~x18 ;
  assign n62 = x11 & n61 ;
  assign n63 = x3 & x17 ;
  assign n64 = ( ~x2 & x5 ) | ( ~x2 & n63 ) | ( x5 & n63 ) ;
  assign n65 = x2 & n64 ;
  assign n66 = ( x2 & x5 ) | ( x2 & ~n65 ) | ( x5 & ~n65 ) ;
  assign n67 = n62 & n66 ;
  assign n68 = ( n62 & n65 ) | ( n62 & ~n67 ) | ( n65 & ~n67 ) ;
  assign n74 = ( ~x0 & n68 ) | ( ~x0 & n73 ) | ( n68 & n73 ) ;
  assign n75 = x1 & ~n74 ;
  assign n76 = ( x1 & n73 ) | ( x1 & ~n75 ) | ( n73 & ~n75 ) ;
  assign n77 = ~x15 & n76 ;
  assign n78 = ( ~n60 & n76 ) | ( ~n60 & n77 ) | ( n76 & n77 ) ;
  assign n80 = n59 | n78 ;
  assign n81 = ( n52 & ~n79 ) | ( n52 & n80 ) | ( ~n79 & n80 ) ;
  assign n82 = x4 & n81 ;
  assign n28 = x1 & x5 ;
  assign n29 = ( x2 & n27 ) | ( x2 & n28 ) | ( n27 & n28 ) ;
  assign n30 = ~n27 & n29 ;
  assign n33 = ( x0 & x7 ) | ( x0 & n30 ) | ( x7 & n30 ) ;
  assign n31 = x1 | x9 ;
  assign n32 = x2 | n31 ;
  assign n34 = x7 & ~n32 ;
  assign n35 = ( ~x0 & n33 ) | ( ~x0 & n34 ) | ( n33 & n34 ) ;
  assign n83 = n35 | n82 ;
  assign n84 = ( x3 & n82 ) | ( x3 & n83 ) | ( n82 & n83 ) ;
  assign n85 = x13 & ~n84 ;
  assign n25 = ~x20 & x22 ;
  assign n26 = x21 & n25 ;
  assign n86 = ~x19 & n26 ;
  assign n87 = x13 | n86 ;
  assign n88 = ~n85 & n87 ;
  assign n92 = ~x3 & x14 ;
  assign n139 = x14 & ~x18 ;
  assign n140 = x3 & n139 ;
  assign n141 = ( x3 & n92 ) | ( x3 & ~n140 ) | ( n92 & ~n140 ) ;
  assign n142 = x16 & ~n141 ;
  assign n143 = x15 & n142 ;
  assign n103 = x15 & x16 ;
  assign n104 = ( x14 & x16 ) | ( x14 & n103 ) | ( x16 & n103 ) ;
  assign n136 = x14 & x15 ;
  assign n137 = ~x3 & n104 ;
  assign n138 = ( n104 & n136 ) | ( n104 & n137 ) | ( n136 & n137 ) ;
  assign n144 = ( x17 & n138 ) | ( x17 & ~n143 ) | ( n138 & ~n143 ) ;
  assign n145 = ~x18 & n144 ;
  assign n146 = ( x18 & ~n143 ) | ( x18 & n145 ) | ( ~n143 & n145 ) ;
  assign n153 = ( x4 & x5 ) | ( x4 & n146 ) | ( x5 & n146 ) ;
  assign n147 = x3 & ~x7 ;
  assign n148 = ~x3 & x6 ;
  assign n149 = ( x3 & ~n147 ) | ( x3 & n148 ) | ( ~n147 & n148 ) ;
  assign n150 = ( x17 & ~x18 ) | ( x17 & n149 ) | ( ~x18 & n149 ) ;
  assign n151 = ( x15 & ~x17 ) | ( x15 & n149 ) | ( ~x17 & n149 ) ;
  assign n152 = n150 & n151 ;
  assign n154 = x5 & n152 ;
  assign n155 = ( ~n146 & n153 ) | ( ~n146 & n154 ) | ( n153 & n154 ) ;
  assign n156 = x2 & ~n155 ;
  assign n127 = ( x16 & x17 ) | ( x16 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n128 = x14 & ~n127 ;
  assign n129 = ( ~x14 & x18 ) | ( ~x14 & n128 ) | ( x18 & n128 ) ;
  assign n130 = ( ~x11 & x15 ) | ( ~x11 & n129 ) | ( x15 & n129 ) ;
  assign n131 = ( x11 & x15 ) | ( x11 & ~x18 ) | ( x15 & ~x18 ) ;
  assign n132 = ~n130 & n131 ;
  assign n133 = x4 & x10 ;
  assign n134 = ( x5 & n132 ) | ( x5 & n133 ) | ( n132 & n133 ) ;
  assign n135 = ~x5 & n134 ;
  assign n157 = ~x2 & n135 ;
  assign n158 = ( x2 & ~n156 ) | ( x2 & n157 ) | ( ~n156 & n157 ) ;
  assign n159 = x1 & ~n158 ;
  assign n122 = ( x15 & x16 ) | ( x15 & ~n27 ) | ( x16 & ~n27 ) ;
  assign n123 = ( n27 & n60 ) | ( n27 & n122 ) | ( n60 & n122 ) ;
  assign n124 = ~x5 & x10 ;
  assign n125 = ( x4 & n123 ) | ( x4 & n124 ) | ( n123 & n124 ) ;
  assign n126 = ~n123 & n125 ;
  assign n160 = x2 & n126 ;
  assign n161 = x1 | n160 ;
  assign n162 = ~n159 & n161 ;
  assign n163 = ~x0 & n162 ;
  assign n97 = x3 & ~x9 ;
  assign n98 = ( ~x18 & n60 ) | ( ~x18 & n97 ) | ( n60 & n97 ) ;
  assign n99 = ~n60 & n98 ;
  assign n93 = x14 & ~n92 ;
  assign n94 = ~x9 & n93 ;
  assign n95 = ( x0 & ~n92 ) | ( x0 & n93 ) | ( ~n92 & n93 ) ;
  assign n96 = ( ~x3 & n94 ) | ( ~x3 & n95 ) | ( n94 & n95 ) ;
  assign n100 = ( ~n27 & n96 ) | ( ~n27 & n99 ) | ( n96 & n99 ) ;
  assign n101 = x16 & ~n100 ;
  assign n102 = ( x16 & n99 ) | ( x16 & ~n101 ) | ( n99 & ~n101 ) ;
  assign n111 = ( x5 & ~x15 ) | ( x5 & n102 ) | ( ~x15 & n102 ) ;
  assign n105 = x0 & ~n104 ;
  assign n106 = ~x3 & n105 ;
  assign n107 = x3 & ~x15 ;
  assign n108 = ( x9 & ~x18 ) | ( x9 & n107 ) | ( ~x18 & n107 ) ;
  assign n109 = ~x9 & n108 ;
  assign n110 = n106 | n109 ;
  assign n112 = ~x5 & n110 ;
  assign n113 = ( n102 & ~n111 ) | ( n102 & n112 ) | ( ~n111 & n112 ) ;
  assign n119 = ( x2 & ~x4 ) | ( x2 & n113 ) | ( ~x4 & n113 ) ;
  assign n114 = ~x6 & x9 ;
  assign n115 = x0 & ~x3 ;
  assign n116 = ( x6 & n114 ) | ( x6 & n115 ) | ( n114 & n115 ) ;
  assign n117 = x7 & n97 ;
  assign n118 = n116 | n117 ;
  assign n120 = ~x2 & n118 ;
  assign n121 = ( n113 & ~n119 ) | ( n113 & n120 ) | ( ~n119 & n120 ) ;
  assign n164 = n121 | n163 ;
  assign n165 = ( ~x1 & n163 ) | ( ~x1 & n164 ) | ( n163 & n164 ) ;
  assign n166 = x13 & n165 ;
  assign n89 = ( ~x19 & x20 ) | ( ~x19 & x22 ) | ( x20 & x22 ) ;
  assign n90 = ( ~x19 & x20 ) | ( ~x19 & x21 ) | ( x20 & x21 ) ;
  assign n91 = n89 & ~n90 ;
  assign n167 = x13 | n91 ;
  assign n168 = ( ~x13 & n166 ) | ( ~x13 & n167 ) | ( n166 & n167 ) ;
  assign n211 = ~x20 & n90 ;
  assign n212 = ( x21 & x22 ) | ( x21 & ~n211 ) | ( x22 & ~n211 ) ;
  assign n213 = ( n90 & n211 ) | ( n90 & ~n212 ) | ( n211 & ~n212 ) ;
  assign n214 = ~x13 & n213 ;
  assign n169 = x15 | x18 ;
  assign n170 = ( x18 & n60 ) | ( x18 & n169 ) | ( n60 & n169 ) ;
  assign n171 = ( x3 & ~x9 ) | ( x3 & n106 ) | ( ~x9 & n106 ) ;
  assign n172 = n170 | n171 ;
  assign n173 = ( n106 & ~n170 ) | ( n106 & n172 ) | ( ~n170 & n172 ) ;
  assign n174 = x4 & n173 ;
  assign n175 = ~x5 & n174 ;
  assign n176 = n118 & ~n175 ;
  assign n177 = x1 | x2 ;
  assign n178 = ( n175 & n176 ) | ( n175 & ~n177 ) | ( n176 & ~n177 ) ;
  assign n188 = ( ~x3 & x14 ) | ( ~x3 & x15 ) | ( x14 & x15 ) ;
  assign n189 = x16 & n188 ;
  assign n193 = ( x5 & x17 ) | ( x5 & n189 ) | ( x17 & n189 ) ;
  assign n190 = x3 & ~x17 ;
  assign n191 = ( ~x18 & n136 ) | ( ~x18 & n190 ) | ( n136 & n190 ) ;
  assign n192 = ~n136 & n191 ;
  assign n194 = x5 & n192 ;
  assign n195 = ( ~n189 & n193 ) | ( ~n189 & n194 ) | ( n193 & n194 ) ;
  assign n196 = x1 & n195 ;
  assign n183 = ~x1 & x5 ;
  assign n184 = x5 & ~n183 ;
  assign n185 = ~n56 & n184 ;
  assign n186 = ( x10 & ~n183 ) | ( x10 & n184 ) | ( ~n183 & n184 ) ;
  assign n187 = ( ~x1 & n185 ) | ( ~x1 & n186 ) | ( n185 & n186 ) ;
  assign n197 = n187 | n196 ;
  assign n198 = ( ~n104 & n196 ) | ( ~n104 & n197 ) | ( n196 & n197 ) ;
  assign n199 = x4 & n198 ;
  assign n179 = ~x15 & x17 ;
  assign n180 = ( x17 & n27 ) | ( x17 & ~n179 ) | ( n27 & ~n179 ) ;
  assign n181 = x5 & n149 ;
  assign n182 = ~n180 & n181 ;
  assign n200 = n182 | n199 ;
  assign n201 = ( x1 & n199 ) | ( x1 & n200 ) | ( n199 & n200 ) ;
  assign n208 = ( x0 & ~x2 ) | ( x0 & n201 ) | ( ~x2 & n201 ) ;
  assign n202 = x11 & ~n170 ;
  assign n203 = ( x5 & x10 ) | ( x5 & n202 ) | ( x10 & n202 ) ;
  assign n204 = ~x5 & n203 ;
  assign n205 = x1 & x4 ;
  assign n206 = ( x2 & n204 ) | ( x2 & n205 ) | ( n204 & n205 ) ;
  assign n207 = ~x2 & n206 ;
  assign n209 = ~x0 & n207 ;
  assign n210 = ( n201 & ~n208 ) | ( n201 & n209 ) | ( ~n208 & n209 ) ;
  assign n215 = n178 | n210 ;
  assign n216 = x13 & n215 ;
  assign n217 = n214 | n216 ;
  assign n238 = ( x20 & x21 ) | ( x20 & x22 ) | ( x21 & x22 ) ;
  assign n239 = ~n89 & n238 ;
  assign n240 = x13 | n239 ;
  assign n218 = x3 & x11 ;
  assign n219 = x8 & n218 ;
  assign n233 = x0 & x1 ;
  assign n234 = x0 & ~n233 ;
  assign n235 = n219 & n234 ;
  assign n230 = ( x5 & n27 ) | ( x5 & n149 ) | ( n27 & n149 ) ;
  assign n221 = x3 | x14 ;
  assign n222 = x15 | n27 ;
  assign n223 = ( ~x3 & n221 ) | ( ~x3 & n222 ) | ( n221 & n222 ) ;
  assign n224 = ( ~x3 & x14 ) | ( ~x3 & n223 ) | ( x14 & n223 ) ;
  assign n225 = ~n56 & n224 ;
  assign n226 = ( n56 & n223 ) | ( n56 & n225 ) | ( n223 & n225 ) ;
  assign n220 = x16 | n180 ;
  assign n227 = ( x4 & n143 ) | ( x4 & ~n220 ) | ( n143 & ~n220 ) ;
  assign n228 = n226 & n227 ;
  assign n229 = ( x4 & ~n226 ) | ( x4 & n228 ) | ( ~n226 & n228 ) ;
  assign n231 = x5 & n229 ;
  assign n232 = ( ~n27 & n230 ) | ( ~n27 & n231 ) | ( n230 & n231 ) ;
  assign n236 = ( n232 & ~n233 ) | ( n232 & n234 ) | ( ~n233 & n234 ) ;
  assign n237 = ( x1 & n235 ) | ( x1 & n236 ) | ( n235 & n236 ) ;
  assign n241 = x2 & n237 ;
  assign n242 = x13 & ~n241 ;
  assign n243 = n240 & ~n242 ;
  assign n244 = ( x15 & x16 ) | ( x15 & x17 ) | ( x16 & x17 ) ;
  assign n245 = ( ~x17 & n60 ) | ( ~x17 & n244 ) | ( n60 & n244 ) ;
  assign n246 = ~x1 & x10 ;
  assign n247 = ( x2 & n245 ) | ( x2 & n246 ) | ( n245 & n246 ) ;
  assign n248 = ~n245 & n247 ;
  assign n261 = ( x0 & x13 ) | ( x0 & n248 ) | ( x13 & n248 ) ;
  assign n256 = ( x15 & ~x18 ) | ( x15 & n41 ) | ( ~x18 & n41 ) ;
  assign n252 = ~x14 & x16 ;
  assign n253 = ( x16 & x18 ) | ( x16 & ~n252 ) | ( x18 & ~n252 ) ;
  assign n254 = ( ~x16 & x17 ) | ( ~x16 & n252 ) | ( x17 & n252 ) ;
  assign n255 = ( ~x17 & n253 ) | ( ~x17 & n254 ) | ( n253 & n254 ) ;
  assign n257 = ( x15 & ~n41 ) | ( x15 & n255 ) | ( ~n41 & n255 ) ;
  assign n258 = n256 & ~n257 ;
  assign n249 = x0 & ~x1 ;
  assign n250 = ( ~x3 & n245 ) | ( ~x3 & n249 ) | ( n245 & n249 ) ;
  assign n251 = ~n245 & n250 ;
  assign n259 = ~x2 & n251 ;
  assign n260 = ( ~x2 & n258 ) | ( ~x2 & n259 ) | ( n258 & n259 ) ;
  assign n262 = x13 & n260 ;
  assign n263 = ( ~x0 & n261 ) | ( ~x0 & n262 ) | ( n261 & n262 ) ;
  assign n264 = x12 & x18 ;
  assign n265 = ( x4 & ~x5 ) | ( x4 & n264 ) | ( ~x5 & n264 ) ;
  assign n266 = n263 & ~n265 ;
  assign n267 = ( n263 & n264 ) | ( n263 & ~n266 ) | ( n264 & ~n266 ) ;
  assign n269 = x16 | x18 ;
  assign n270 = ( x16 & ~x17 ) | ( x16 & n269 ) | ( ~x17 & n269 ) ;
  assign n271 = ( x3 & ~n252 ) | ( x3 & n270 ) | ( ~n252 & n270 ) ;
  assign n268 = ( x14 & x18 ) | ( x14 & n27 ) | ( x18 & n27 ) ;
  assign n272 = ( ~x3 & n268 ) | ( ~x3 & n270 ) | ( n268 & n270 ) ;
  assign n273 = n271 & n272 ;
  assign n274 = ( x2 & n28 ) | ( x2 & n273 ) | ( n28 & n273 ) ;
  assign n275 = ~n273 & n274 ;
  assign n301 = ( x0 & x15 ) | ( x0 & n275 ) | ( x15 & n275 ) ;
  assign n281 = ~x2 & n96 ;
  assign n282 = ~x1 & n281 ;
  assign n276 = ~x1 & x2 ;
  assign n277 = x1 & x14 ;
  assign n278 = ~x2 & x11 ;
  assign n279 = x14 & ~n278 ;
  assign n280 = ( n276 & n277 ) | ( n276 & ~n279 ) | ( n277 & ~n279 ) ;
  assign n283 = ( ~x0 & n280 ) | ( ~x0 & n282 ) | ( n280 & n282 ) ;
  assign n284 = x10 & ~n283 ;
  assign n285 = ( x10 & n282 ) | ( x10 & ~n284 ) | ( n282 & ~n284 ) ;
  assign n286 = ~n27 & n285 ;
  assign n298 = ( x5 & ~x16 ) | ( x5 & n286 ) | ( ~x16 & n286 ) ;
  assign n287 = ( x1 & ~x16 ) | ( x1 & n115 ) | ( ~x16 & n115 ) ;
  assign n288 = ~x1 & n287 ;
  assign n289 = ~x18 & n41 ;
  assign n290 = ~n60 & n289 ;
  assign n291 = x2 & ~x16 ;
  assign n292 = x10 & n291 ;
  assign n293 = ~x0 & n292 ;
  assign n294 = ~x1 & n293 ;
  assign n295 = ( ~n288 & n290 ) | ( ~n288 & n294 ) | ( n290 & n294 ) ;
  assign n296 = x2 & ~n294 ;
  assign n297 = ( n288 & n295 ) | ( n288 & ~n296 ) | ( n295 & ~n296 ) ;
  assign n299 = ~x5 & n297 ;
  assign n300 = ( n286 & ~n298 ) | ( n286 & n299 ) | ( ~n298 & n299 ) ;
  assign n302 = x15 & n300 ;
  assign n303 = ( ~x0 & n301 ) | ( ~x0 & n302 ) | ( n301 & n302 ) ;
  assign n304 = ( x4 & n264 ) | ( x4 & n303 ) | ( n264 & n303 ) ;
  assign n305 = x13 & ~n304 ;
  assign n306 = ( x13 & n264 ) | ( x13 & ~n305 ) | ( n264 & ~n305 ) ;
  assign n307 = ( ~x3 & x6 ) | ( ~x3 & x8 ) | ( x6 & x8 ) ;
  assign n308 = ~x9 & n307 ;
  assign n309 = ( ~x3 & x9 ) | ( ~x3 & n308 ) | ( x9 & n308 ) ;
  assign n310 = x0 | n117 ;
  assign n311 = ( n117 & n309 ) | ( n117 & n310 ) | ( n309 & n310 ) ;
  assign n312 = ~x1 & x13 ;
  assign n313 = ( x2 & n311 ) | ( x2 & ~n312 ) | ( n311 & ~n312 ) ;
  assign n314 = n311 & ~n313 ;
  assign n326 = ( x16 & n56 ) | ( x16 & n60 ) | ( n56 & n60 ) ;
  assign n315 = ( x16 & x17 ) | ( x16 & x18 ) | ( x17 & x18 ) ;
  assign n316 = x14 & ~n315 ;
  assign n317 = ( x14 & x18 ) | ( x14 & ~n316 ) | ( x18 & ~n316 ) ;
  assign n327 = x9 | n317 ;
  assign n328 = ( x2 & x3 ) | ( x2 & ~n327 ) | ( x3 & ~n327 ) ;
  assign n329 = ~x2 & n328 ;
  assign n321 = x0 & x2 ;
  assign n322 = x2 & ~n321 ;
  assign n323 = x10 & n322 ;
  assign n324 = ( x3 & n321 ) | ( x3 & ~n322 ) | ( n321 & ~n322 ) ;
  assign n325 = ( x0 & n323 ) | ( x0 & ~n324 ) | ( n323 & ~n324 ) ;
  assign n330 = n325 | n329 ;
  assign n331 = ( ~n326 & n329 ) | ( ~n326 & n330 ) | ( n329 & n330 ) ;
  assign n332 = x1 | n331 ;
  assign n318 = x11 & ~n317 ;
  assign n319 = ( x2 & x10 ) | ( x2 & n318 ) | ( x10 & n318 ) ;
  assign n320 = ~x2 & n319 ;
  assign n333 = ~x0 & n320 ;
  assign n334 = x1 & ~n333 ;
  assign n335 = n332 & ~n334 ;
  assign n336 = ~x5 & x15 ;
  assign n337 = ( x13 & ~n335 ) | ( x13 & n336 ) | ( ~n335 & n336 ) ;
  assign n338 = n335 & n337 ;
  assign n339 = n264 | n338 ;
  assign n340 = ( x4 & n264 ) | ( x4 & n339 ) | ( n264 & n339 ) ;
  assign n343 = ( x5 & ~x6 ) | ( x5 & n104 ) | ( ~x6 & n104 ) ;
  assign n344 = x4 & n343 ;
  assign n345 = ( x4 & x6 ) | ( x4 & ~n344 ) | ( x6 & ~n344 ) ;
  assign n346 = ( x1 & ~x2 ) | ( x1 & n345 ) | ( ~x2 & n345 ) ;
  assign n347 = ~x2 & x8 ;
  assign n348 = ( ~x1 & n346 ) | ( ~x1 & n347 ) | ( n346 & n347 ) ;
  assign n349 = x0 & n348 ;
  assign n341 = x6 & ~n56 ;
  assign n342 = x5 & n341 ;
  assign n350 = n342 | n349 ;
  assign n351 = ( n46 & n349 ) | ( n46 & n350 ) | ( n349 & n350 ) ;
  assign n390 = ( x3 & ~x13 ) | ( x3 & n351 ) | ( ~x13 & n351 ) ;
  assign n363 = x5 & ~n56 ;
  assign n364 = n46 & n363 ;
  assign n365 = ~x15 & n60 ;
  assign n366 = x5 | x9 ;
  assign n367 = ( n60 & ~n365 ) | ( n60 & n366 ) | ( ~n365 & n366 ) ;
  assign n368 = x5 & ~n136 ;
  assign n369 = ~x17 & n368 ;
  assign n370 = x2 & n369 ;
  assign n371 = ( x0 & x1 ) | ( x0 & n370 ) | ( x1 & n370 ) ;
  assign n372 = ~x0 & n371 ;
  assign n373 = ( x1 & x2 ) | ( x1 & ~n372 ) | ( x2 & ~n372 ) ;
  assign n374 = ~n367 & n373 ;
  assign n375 = ( n367 & ~n372 ) | ( n367 & n374 ) | ( ~n372 & n374 ) ;
  assign n381 = ( x4 & ~x18 ) | ( x4 & n375 ) | ( ~x18 & n375 ) ;
  assign n376 = x23 & ~n136 ;
  assign n377 = x5 & n376 ;
  assign n378 = x2 & n377 ;
  assign n379 = ( x0 & x1 ) | ( x0 & n378 ) | ( x1 & n378 ) ;
  assign n380 = ~x0 & n379 ;
  assign n382 = ~x18 & n380 ;
  assign n383 = ( ~n375 & n381 ) | ( ~n375 & n382 ) | ( n381 & n382 ) ;
  assign n384 = ( n32 & n364 ) | ( n32 & ~n383 ) | ( n364 & ~n383 ) ;
  assign n385 = x7 | n383 ;
  assign n386 = ( n364 & ~n384 ) | ( n364 & n385 ) | ( ~n384 & n385 ) ;
  assign n387 = x3 & n386 ;
  assign n355 = ( x1 & x4 ) | ( x1 & n124 ) | ( x4 & n124 ) ;
  assign n356 = ~x1 & n355 ;
  assign n352 = ( x4 & x17 ) | ( x4 & ~x18 ) | ( x17 & ~x18 ) ;
  assign n353 = ~x18 & x23 ;
  assign n354 = ( ~x17 & n352 ) | ( ~x17 & n353 ) | ( n352 & n353 ) ;
  assign n357 = ( x1 & n354 ) | ( x1 & n356 ) | ( n354 & n356 ) ;
  assign n358 = x5 & ~n357 ;
  assign n359 = ( x5 & n356 ) | ( x5 & ~n358 ) | ( n356 & ~n358 ) ;
  assign n360 = ( ~n104 & n207 ) | ( ~n104 & n359 ) | ( n207 & n359 ) ;
  assign n361 = x2 & ~n360 ;
  assign n362 = ( x2 & n207 ) | ( x2 & ~n361 ) | ( n207 & ~n361 ) ;
  assign n388 = n362 | n387 ;
  assign n389 = ( ~x0 & n387 ) | ( ~x0 & n388 ) | ( n387 & n388 ) ;
  assign n391 = x13 & n389 ;
  assign n392 = ( n351 & ~n390 ) | ( n351 & n391 ) | ( ~n390 & n391 ) ;
  assign n404 = ( x3 & x14 ) | ( x3 & x17 ) | ( x14 & x17 ) ;
  assign n405 = ~x16 & x17 ;
  assign n406 = ( ~x14 & n404 ) | ( ~x14 & n405 ) | ( n404 & n405 ) ;
  assign n407 = ( x2 & n28 ) | ( x2 & ~n406 ) | ( n28 & ~n406 ) ;
  assign n408 = n406 & n407 ;
  assign n416 = ( x0 & x4 ) | ( x0 & n408 ) | ( x4 & n408 ) ;
  assign n413 = ( x5 & x16 ) | ( x5 & n286 ) | ( x16 & n286 ) ;
  assign n409 = x5 & ~n141 ;
  assign n410 = x2 & n409 ;
  assign n411 = ( x0 & x1 ) | ( x0 & n410 ) | ( x1 & n410 ) ;
  assign n412 = ~x0 & n411 ;
  assign n414 = x16 & n412 ;
  assign n415 = ( ~x5 & n413 ) | ( ~x5 & n414 ) | ( n413 & n414 ) ;
  assign n417 = x4 & n415 ;
  assign n418 = ( ~x0 & n416 ) | ( ~x0 & n417 ) | ( n416 & n417 ) ;
  assign n398 = ( x3 & ~x7 ) | ( x3 & x17 ) | ( ~x7 & x17 ) ;
  assign n397 = n60 & n353 ;
  assign n399 = x3 & n397 ;
  assign n400 = ( x7 & n398 ) | ( x7 & n399 ) | ( n398 & n399 ) ;
  assign n394 = ( x3 & x6 ) | ( x3 & ~x17 ) | ( x6 & ~x17 ) ;
  assign n393 = n252 & n353 ;
  assign n395 = ~x3 & n393 ;
  assign n396 = ( x6 & ~n394 ) | ( x6 & n395 ) | ( ~n394 & n395 ) ;
  assign n401 = n396 & ~n400 ;
  assign n402 = x2 & x5 ;
  assign n403 = ( n400 & n401 ) | ( n400 & n402 ) | ( n401 & n402 ) ;
  assign n419 = ( ~x0 & n403 ) | ( ~x0 & n418 ) | ( n403 & n418 ) ;
  assign n420 = x1 & ~n419 ;
  assign n421 = ( x1 & n418 ) | ( x1 & ~n420 ) | ( n418 & ~n420 ) ;
  assign n433 = ( x13 & x15 ) | ( x13 & ~n421 ) | ( x15 & ~n421 ) ;
  assign n422 = x4 & ~n60 ;
  assign n423 = x6 | n422 ;
  assign n424 = ( ~x3 & n422 ) | ( ~x3 & n423 ) | ( n422 & n423 ) ;
  assign n425 = ( ~x4 & x7 ) | ( ~x4 & n424 ) | ( x7 & n424 ) ;
  assign n426 = x3 | n424 ;
  assign n427 = ( x4 & n425 ) | ( x4 & n426 ) | ( n425 & n426 ) ;
  assign n428 = ( x5 & n179 ) | ( x5 & ~n427 ) | ( n179 & ~n427 ) ;
  assign n429 = n427 & n428 ;
  assign n430 = x2 & n429 ;
  assign n431 = ( x0 & x1 ) | ( x0 & n430 ) | ( x1 & n430 ) ;
  assign n432 = ~x0 & n431 ;
  assign n434 = x13 & n432 ;
  assign n435 = ( n421 & n433 ) | ( n421 & n434 ) | ( n433 & n434 ) ;
  assign n443 = ( ~x18 & n60 ) | ( ~x18 & n278 ) | ( n60 & n278 ) ;
  assign n444 = ~n60 & n443 ;
  assign n446 = ( x1 & x15 ) | ( x1 & ~n444 ) | ( x15 & ~n444 ) ;
  assign n445 = n42 & n280 ;
  assign n447 = x15 & n445 ;
  assign n448 = ( n444 & n446 ) | ( n444 & n447 ) | ( n446 & n447 ) ;
  assign n436 = x11 & ~x15 ;
  assign n437 = ~x18 & n436 ;
  assign n438 = x1 & x2 ;
  assign n439 = x1 & ~n438 ;
  assign n440 = n437 & n439 ;
  assign n441 = ( n104 & n438 ) | ( n104 & ~n439 ) | ( n438 & ~n439 ) ;
  assign n442 = ( x2 & n440 ) | ( x2 & ~n441 ) | ( n440 & ~n441 ) ;
  assign n449 = n442 & ~n448 ;
  assign n450 = x10 & x13 ;
  assign n451 = ( n448 & n449 ) | ( n448 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ~x5 & n451 ;
  assign n453 = ( x0 & x4 ) | ( x0 & n452 ) | ( x4 & n452 ) ;
  assign n454 = ~x0 & n453 ;
  assign n455 = x0 & ~x2 ;
  assign n456 = ( x1 & ~x3 ) | ( x1 & n455 ) | ( ~x3 & n455 ) ;
  assign n457 = ~x1 & n456 ;
  assign n458 = x13 & n457 ;
  assign n459 = x9 & n458 ;
  assign n460 = ( x1 & x2 ) | ( x1 & ~x13 ) | ( x2 & ~x13 ) ;
  assign n461 = ( x2 & ~x3 ) | ( x2 & x13 ) | ( ~x3 & x13 ) ;
  assign n462 = ~n460 & n461 ;
  assign n463 = x8 & n462 ;
  assign n464 = x0 & n463 ;
  assign n465 = x15 & ~x17 ;
  assign n466 = ( x5 & ~x18 ) | ( x5 & n465 ) | ( ~x18 & n465 ) ;
  assign n467 = ~x5 & n466 ;
  assign y0 = n88 ;
  assign y1 = n168 ;
  assign y2 = n217 ;
  assign y3 = n243 ;
  assign y4 = n267 ;
  assign y5 = n306 ;
  assign y6 = n314 ;
  assign y7 = n340 ;
  assign y8 = n392 ;
  assign y9 = n435 ;
  assign y10 = n454 ;
  assign y11 = n459 ;
  assign y12 = n464 ;
  assign y13 = n467 ;
endmodule
