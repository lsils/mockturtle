module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 ;
  wire n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 ;
  assign n95 = ~x87 & x89 ;
  assign n96 = ( x85 & x86 ) | ( x85 & n95 ) | ( x86 & n95 ) ;
  assign n97 = ~x86 & n96 ;
  assign n98 = ( x28 & ~x91 ) | ( x28 & n97 ) | ( ~x91 & n97 ) ;
  assign n99 = x4 | x88 ;
  assign n100 = ( ~x28 & x91 ) | ( ~x28 & n99 ) | ( x91 & n99 ) ;
  assign n101 = n98 & n100 ;
  assign n102 = ( x29 & ~x50 ) | ( x29 & n101 ) | ( ~x50 & n101 ) ;
  assign n103 = x50 & ~x86 ;
  assign n104 = ( x85 & ~n99 ) | ( x85 & n103 ) | ( ~n99 & n103 ) ;
  assign n105 = n99 & n104 ;
  assign n106 = ( x87 & ~x89 ) | ( x87 & x90 ) | ( ~x89 & x90 ) ;
  assign n107 = n105 & n106 ;
  assign n108 = ( x90 & ~n105 ) | ( x90 & n107 ) | ( ~n105 & n107 ) ;
  assign n109 = ~x29 & n108 ;
  assign n110 = ( n101 & ~n102 ) | ( n101 & n109 ) | ( ~n102 & n109 ) ;
  assign n111 = ~x3 & x28 ;
  assign n112 = ( x2 & ~x4 ) | ( x2 & n111 ) | ( ~x4 & n111 ) ;
  assign n113 = ~x2 & n112 ;
  assign n114 = x27 & ~x58 ;
  assign n115 = ( x27 & n113 ) | ( x27 & n114 ) | ( n113 & n114 ) ;
  assign n116 = ( x48 & ~x93 ) | ( x48 & n115 ) | ( ~x93 & n115 ) ;
  assign n117 = x30 | x93 ;
  assign n118 = ( x26 & x30 ) | ( x26 & n117 ) | ( x30 & n117 ) ;
  assign n119 = ~x48 & n118 ;
  assign n120 = ( n115 & ~n116 ) | ( n115 & n119 ) | ( ~n116 & n119 ) ;
  assign n121 = x87 | x89 ;
  assign n122 = ( ~x86 & x88 ) | ( ~x86 & n121 ) | ( x88 & n121 ) ;
  assign n123 = x86 | n122 ;
  assign n124 = x85 & ~n123 ;
  assign n125 = x50 & n124 ;
  assign n126 = x31 & ~x48 ;
  assign n127 = ( ~x48 & n125 ) | ( ~x48 & n126 ) | ( n125 & n126 ) ;
  assign n128 = x93 & n115 ;
  assign n129 = ( x27 & x29 ) | ( x27 & ~x93 ) | ( x29 & ~x93 ) ;
  assign n130 = x29 | x32 ;
  assign n131 = ( ~x27 & n129 ) | ( ~x27 & n130 ) | ( n129 & n130 ) ;
  assign n132 = n128 | n131 ;
  assign n133 = x50 & ~x88 ;
  assign n134 = ( x87 & ~x89 ) | ( x87 & n133 ) | ( ~x89 & n133 ) ;
  assign n135 = ~x87 & n134 ;
  assign n136 = ( x33 & x85 ) | ( x33 & ~x86 ) | ( x85 & ~x86 ) ;
  assign n137 = n135 & ~n136 ;
  assign n138 = ( x33 & n135 ) | ( x33 & ~n137 ) | ( n135 & ~n137 ) ;
  assign n139 = ~x48 & n138 ;
  assign n140 = ~x29 & n139 ;
  assign n141 = ~x29 & x34 ;
  assign n142 = ~x48 & n141 ;
  assign n143 = ~x29 & x35 ;
  assign n144 = ~x48 & n143 ;
  assign n145 = ~x29 & x36 ;
  assign n146 = ~x48 & n145 ;
  assign n147 = ~x29 & x37 ;
  assign n148 = ~x48 & n147 ;
  assign n149 = ~x29 & x38 ;
  assign n150 = ~x48 & n149 ;
  assign n151 = ~x29 & x39 ;
  assign n152 = ~x48 & n151 ;
  assign n153 = x1 & ~x29 ;
  assign n154 = x0 & ~x29 ;
  assign n155 = ~x29 & x41 ;
  assign n156 = ~x29 & x42 ;
  assign n157 = ~x29 & x43 ;
  assign n158 = ~x29 & x44 ;
  assign n159 = ~x29 & x45 ;
  assign n160 = ~x29 & x46 ;
  assign n161 = x26 & ~x93 ;
  assign n162 = ~x86 & x89 ;
  assign n163 = ( x87 & n99 ) | ( x87 & ~n162 ) | ( n99 & ~n162 ) ;
  assign n164 = n99 & ~n163 ;
  assign n165 = ( x50 & n128 ) | ( x50 & n164 ) | ( n128 & n164 ) ;
  assign n166 = x85 & ~n165 ;
  assign n167 = ( x85 & n128 ) | ( x85 & ~n166 ) | ( n128 & ~n166 ) ;
  assign n168 = x29 | n167 ;
  assign n169 = ( x26 & ~n161 ) | ( x26 & n168 ) | ( ~n161 & n168 ) ;
  assign n170 = ~x27 & x29 ;
  assign n171 = ( ~x58 & n113 ) | ( ~x58 & n170 ) | ( n113 & n170 ) ;
  assign n172 = ~n113 & n171 ;
  assign n173 = x93 & n172 ;
  assign n174 = x83 & x84 ;
  assign n175 = ~x49 & x82 ;
  assign n176 = ( x49 & n174 ) | ( x49 & ~n175 ) | ( n174 & ~n175 ) ;
  assign n177 = ~x48 & x50 ;
  assign n178 = ( ~x48 & n176 ) | ( ~x48 & n177 ) | ( n176 & n177 ) ;
  assign n179 = ~x85 & x86 ;
  assign n180 = n135 & n179 ;
  assign n181 = x51 & ~n180 ;
  assign n182 = x86 & ~x88 ;
  assign n183 = ( x87 & ~x89 ) | ( x87 & n182 ) | ( ~x89 & n182 ) ;
  assign n184 = ~x87 & n183 ;
  assign n185 = ~x85 & n184 ;
  assign n186 = ( x34 & x50 ) | ( x34 & n185 ) | ( x50 & n185 ) ;
  assign n187 = ~x34 & n186 ;
  assign n188 = x48 | n187 ;
  assign n189 = ( n180 & n181 ) | ( n180 & ~n188 ) | ( n181 & ~n188 ) ;
  assign n190 = x52 & ~n180 ;
  assign n191 = ( x35 & x50 ) | ( x35 & n185 ) | ( x50 & n185 ) ;
  assign n192 = ~x35 & n191 ;
  assign n193 = x48 | n192 ;
  assign n194 = ( n180 & n190 ) | ( n180 & ~n193 ) | ( n190 & ~n193 ) ;
  assign n195 = x53 & ~n180 ;
  assign n196 = ( x36 & x50 ) | ( x36 & n185 ) | ( x50 & n185 ) ;
  assign n197 = ~x36 & n196 ;
  assign n198 = x48 | n197 ;
  assign n199 = ( n180 & n195 ) | ( n180 & ~n198 ) | ( n195 & ~n198 ) ;
  assign n200 = x54 & ~n180 ;
  assign n201 = ( x37 & x50 ) | ( x37 & n185 ) | ( x50 & n185 ) ;
  assign n202 = ~x37 & n201 ;
  assign n203 = x48 | n202 ;
  assign n204 = ( n180 & n200 ) | ( n180 & ~n203 ) | ( n200 & ~n203 ) ;
  assign n205 = x55 & ~n180 ;
  assign n206 = ( x38 & x50 ) | ( x38 & n185 ) | ( x50 & n185 ) ;
  assign n207 = ~x38 & n206 ;
  assign n208 = x48 | n207 ;
  assign n209 = ( n180 & n205 ) | ( n180 & ~n208 ) | ( n205 & ~n208 ) ;
  assign n210 = x56 & ~n180 ;
  assign n211 = ( x39 & x50 ) | ( x39 & n185 ) | ( x50 & n185 ) ;
  assign n212 = ~x39 & n211 ;
  assign n213 = x48 | n212 ;
  assign n214 = ( n180 & n210 ) | ( n180 & ~n213 ) | ( n210 & ~n213 ) ;
  assign n215 = ~x48 & x57 ;
  assign n216 = ( ~x48 & n125 ) | ( ~x48 & n215 ) | ( n125 & n215 ) ;
  assign n217 = ~x3 & n174 ;
  assign n218 = ( x2 & ~x82 ) | ( x2 & n217 ) | ( ~x82 & n217 ) ;
  assign n219 = ~x2 & n218 ;
  assign n220 = x29 | x93 ;
  assign n221 = ( x27 & x29 ) | ( x27 & n220 ) | ( x29 & n220 ) ;
  assign n222 = x58 & ~n221 ;
  assign n223 = ( n219 & ~n221 ) | ( n219 & n222 ) | ( ~n221 & n222 ) ;
  assign n224 = ( x2 & x3 ) | ( x2 & x58 ) | ( x3 & x58 ) ;
  assign n225 = x28 & n224 ;
  assign n226 = ( ~x28 & x58 ) | ( ~x28 & n225 ) | ( x58 & n225 ) ;
  assign n227 = x93 & n226 ;
  assign n228 = x27 & n227 ;
  assign n229 = ~x32 & x50 ;
  assign n230 = ( ~x60 & n228 ) | ( ~x60 & n229 ) | ( n228 & n229 ) ;
  assign n231 = ~n228 & n230 ;
  assign n232 = ~x2 & x28 ;
  assign n233 = ~x3 & n232 ;
  assign n234 = x27 & x93 ;
  assign n235 = ( x58 & n233 ) | ( x58 & n234 ) | ( n233 & n234 ) ;
  assign n236 = ~n233 & n235 ;
  assign n237 = x59 & ~n236 ;
  assign n238 = ~n229 & n237 ;
  assign n239 = ( ~x4 & x58 ) | ( ~x4 & n234 ) | ( x58 & n234 ) ;
  assign n240 = x4 & n239 ;
  assign n241 = ( ~x29 & n238 ) | ( ~x29 & n240 ) | ( n238 & n240 ) ;
  assign n242 = ~n231 & n241 ;
  assign n243 = ( ~x29 & n231 ) | ( ~x29 & n242 ) | ( n231 & n242 ) ;
  assign n244 = ( x29 & x60 ) | ( x29 & ~n229 ) | ( x60 & ~n229 ) ;
  assign n245 = ( x29 & ~x61 ) | ( x29 & n229 ) | ( ~x61 & n229 ) ;
  assign n246 = n244 | n245 ;
  assign n247 = x27 & ~n113 ;
  assign n248 = ( x58 & n246 ) | ( x58 & n247 ) | ( n246 & n247 ) ;
  assign n249 = x93 & ~n248 ;
  assign n250 = ( x93 & n246 ) | ( x93 & ~n249 ) | ( n246 & ~n249 ) ;
  assign n251 = ( x58 & n229 ) | ( x58 & n247 ) | ( n229 & n247 ) ;
  assign n252 = x93 & ~n251 ;
  assign n253 = ( x93 & n229 ) | ( x93 & ~n252 ) | ( n229 & ~n252 ) ;
  assign n254 = ( ~x29 & x61 ) | ( ~x29 & n253 ) | ( x61 & n253 ) ;
  assign n255 = ( x58 & n113 ) | ( x58 & n234 ) | ( n113 & n234 ) ;
  assign n256 = ~n113 & n255 ;
  assign n257 = ~x32 & x62 ;
  assign n258 = ( x50 & n256 ) | ( x50 & n257 ) | ( n256 & n257 ) ;
  assign n259 = ~n256 & n258 ;
  assign n260 = ~x29 & n259 ;
  assign n261 = ( ~n253 & n254 ) | ( ~n253 & n260 ) | ( n254 & n260 ) ;
  assign n262 = ~x29 & x93 ;
  assign n263 = x58 & n262 ;
  assign n264 = ( n247 & n261 ) | ( n247 & n263 ) | ( n261 & n263 ) ;
  assign n265 = x5 & ~n264 ;
  assign n266 = ( x5 & n261 ) | ( x5 & ~n265 ) | ( n261 & ~n265 ) ;
  assign n267 = ( ~x29 & x62 ) | ( ~x29 & n253 ) | ( x62 & n253 ) ;
  assign n268 = ~x32 & x63 ;
  assign n269 = ( x50 & n256 ) | ( x50 & n268 ) | ( n256 & n268 ) ;
  assign n270 = ~n256 & n269 ;
  assign n271 = ~x29 & n270 ;
  assign n272 = ( ~n253 & n267 ) | ( ~n253 & n271 ) | ( n267 & n271 ) ;
  assign n273 = ( n247 & n263 ) | ( n247 & n272 ) | ( n263 & n272 ) ;
  assign n274 = x6 & ~n273 ;
  assign n275 = ( x6 & n272 ) | ( x6 & ~n274 ) | ( n272 & ~n274 ) ;
  assign n276 = ( ~x29 & x63 ) | ( ~x29 & n253 ) | ( x63 & n253 ) ;
  assign n277 = ~x32 & x64 ;
  assign n278 = ( x50 & n256 ) | ( x50 & n277 ) | ( n256 & n277 ) ;
  assign n279 = ~n256 & n278 ;
  assign n280 = ~x29 & n279 ;
  assign n281 = ( ~n253 & n276 ) | ( ~n253 & n280 ) | ( n276 & n280 ) ;
  assign n282 = ( n247 & n263 ) | ( n247 & n281 ) | ( n263 & n281 ) ;
  assign n283 = x7 & ~n282 ;
  assign n284 = ( x7 & n281 ) | ( x7 & ~n283 ) | ( n281 & ~n283 ) ;
  assign n285 = ( ~x29 & x64 ) | ( ~x29 & n253 ) | ( x64 & n253 ) ;
  assign n286 = ~x32 & x65 ;
  assign n287 = ( x50 & n256 ) | ( x50 & n286 ) | ( n256 & n286 ) ;
  assign n288 = ~n256 & n287 ;
  assign n289 = ~x29 & n288 ;
  assign n290 = ( ~n253 & n285 ) | ( ~n253 & n289 ) | ( n285 & n289 ) ;
  assign n291 = ( n247 & n263 ) | ( n247 & n290 ) | ( n263 & n290 ) ;
  assign n292 = x8 & ~n291 ;
  assign n293 = ( x8 & n290 ) | ( x8 & ~n292 ) | ( n290 & ~n292 ) ;
  assign n294 = ( ~x29 & x65 ) | ( ~x29 & n253 ) | ( x65 & n253 ) ;
  assign n295 = ~x32 & x66 ;
  assign n296 = ( x50 & n256 ) | ( x50 & n295 ) | ( n256 & n295 ) ;
  assign n297 = ~n256 & n296 ;
  assign n298 = ~x29 & n297 ;
  assign n299 = ( ~n253 & n294 ) | ( ~n253 & n298 ) | ( n294 & n298 ) ;
  assign n300 = ( n247 & n263 ) | ( n247 & n299 ) | ( n263 & n299 ) ;
  assign n301 = x9 & ~n300 ;
  assign n302 = ( x9 & n299 ) | ( x9 & ~n301 ) | ( n299 & ~n301 ) ;
  assign n303 = ( ~x29 & x66 ) | ( ~x29 & n253 ) | ( x66 & n253 ) ;
  assign n304 = ~x32 & x67 ;
  assign n305 = ( x50 & n256 ) | ( x50 & n304 ) | ( n256 & n304 ) ;
  assign n306 = ~n256 & n305 ;
  assign n307 = ~x29 & n306 ;
  assign n308 = ( ~n253 & n303 ) | ( ~n253 & n307 ) | ( n303 & n307 ) ;
  assign n309 = ( n247 & n263 ) | ( n247 & n308 ) | ( n263 & n308 ) ;
  assign n310 = x10 & ~n309 ;
  assign n311 = ( x10 & n308 ) | ( x10 & ~n310 ) | ( n308 & ~n310 ) ;
  assign n312 = ( ~x29 & x67 ) | ( ~x29 & n253 ) | ( x67 & n253 ) ;
  assign n313 = ~x32 & x68 ;
  assign n314 = ( x50 & n256 ) | ( x50 & n313 ) | ( n256 & n313 ) ;
  assign n315 = ~n256 & n314 ;
  assign n316 = ~x29 & n315 ;
  assign n317 = ( ~n253 & n312 ) | ( ~n253 & n316 ) | ( n312 & n316 ) ;
  assign n318 = ( n247 & n263 ) | ( n247 & n317 ) | ( n263 & n317 ) ;
  assign n319 = x11 & ~n318 ;
  assign n320 = ( x11 & n317 ) | ( x11 & ~n319 ) | ( n317 & ~n319 ) ;
  assign n321 = ( ~x29 & x68 ) | ( ~x29 & n253 ) | ( x68 & n253 ) ;
  assign n322 = ~x32 & x69 ;
  assign n323 = ( x50 & n256 ) | ( x50 & n322 ) | ( n256 & n322 ) ;
  assign n324 = ~n256 & n323 ;
  assign n325 = ~x29 & n324 ;
  assign n326 = ( ~n253 & n321 ) | ( ~n253 & n325 ) | ( n321 & n325 ) ;
  assign n327 = ( n247 & n263 ) | ( n247 & n326 ) | ( n263 & n326 ) ;
  assign n328 = x12 & ~n327 ;
  assign n329 = ( x12 & n326 ) | ( x12 & ~n328 ) | ( n326 & ~n328 ) ;
  assign n330 = ( ~x29 & x69 ) | ( ~x29 & n253 ) | ( x69 & n253 ) ;
  assign n331 = ~x32 & x70 ;
  assign n332 = ( x50 & n256 ) | ( x50 & n331 ) | ( n256 & n331 ) ;
  assign n333 = ~n256 & n332 ;
  assign n334 = ~x29 & n333 ;
  assign n335 = ( ~n253 & n330 ) | ( ~n253 & n334 ) | ( n330 & n334 ) ;
  assign n336 = ( n247 & n263 ) | ( n247 & n335 ) | ( n263 & n335 ) ;
  assign n337 = x13 & ~n336 ;
  assign n338 = ( x13 & n335 ) | ( x13 & ~n337 ) | ( n335 & ~n337 ) ;
  assign n339 = ( ~x29 & x70 ) | ( ~x29 & n253 ) | ( x70 & n253 ) ;
  assign n340 = ~x32 & x71 ;
  assign n341 = ( x50 & n256 ) | ( x50 & n340 ) | ( n256 & n340 ) ;
  assign n342 = ~n256 & n341 ;
  assign n343 = ~x29 & n342 ;
  assign n344 = ( ~n253 & n339 ) | ( ~n253 & n343 ) | ( n339 & n343 ) ;
  assign n345 = ( n247 & n263 ) | ( n247 & n344 ) | ( n263 & n344 ) ;
  assign n346 = x14 & ~n345 ;
  assign n347 = ( x14 & n344 ) | ( x14 & ~n346 ) | ( n344 & ~n346 ) ;
  assign n348 = ( ~x29 & x71 ) | ( ~x29 & n253 ) | ( x71 & n253 ) ;
  assign n349 = ~x32 & x72 ;
  assign n350 = ( x50 & n256 ) | ( x50 & n349 ) | ( n256 & n349 ) ;
  assign n351 = ~n256 & n350 ;
  assign n352 = ~x29 & n351 ;
  assign n353 = ( ~n253 & n348 ) | ( ~n253 & n352 ) | ( n348 & n352 ) ;
  assign n354 = ( n247 & n263 ) | ( n247 & n353 ) | ( n263 & n353 ) ;
  assign n355 = x15 & ~n354 ;
  assign n356 = ( x15 & n353 ) | ( x15 & ~n355 ) | ( n353 & ~n355 ) ;
  assign n357 = ( ~x29 & x72 ) | ( ~x29 & n253 ) | ( x72 & n253 ) ;
  assign n358 = ~x32 & x73 ;
  assign n359 = ( x50 & n256 ) | ( x50 & n358 ) | ( n256 & n358 ) ;
  assign n360 = ~n256 & n359 ;
  assign n361 = ~x29 & n360 ;
  assign n362 = ( ~n253 & n357 ) | ( ~n253 & n361 ) | ( n357 & n361 ) ;
  assign n363 = ( n247 & n263 ) | ( n247 & n362 ) | ( n263 & n362 ) ;
  assign n364 = x16 & ~n363 ;
  assign n365 = ( x16 & n362 ) | ( x16 & ~n364 ) | ( n362 & ~n364 ) ;
  assign n366 = ( ~x29 & x73 ) | ( ~x29 & n253 ) | ( x73 & n253 ) ;
  assign n367 = ~x32 & x74 ;
  assign n368 = ( x50 & n256 ) | ( x50 & n367 ) | ( n256 & n367 ) ;
  assign n369 = ~n256 & n368 ;
  assign n370 = ~x29 & n369 ;
  assign n371 = ( ~n253 & n366 ) | ( ~n253 & n370 ) | ( n366 & n370 ) ;
  assign n372 = ( n247 & n263 ) | ( n247 & n371 ) | ( n263 & n371 ) ;
  assign n373 = x17 & ~n372 ;
  assign n374 = ( x17 & n371 ) | ( x17 & ~n373 ) | ( n371 & ~n373 ) ;
  assign n375 = ( ~x29 & x74 ) | ( ~x29 & n253 ) | ( x74 & n253 ) ;
  assign n376 = ~x32 & x75 ;
  assign n377 = ( x50 & n256 ) | ( x50 & n376 ) | ( n256 & n376 ) ;
  assign n378 = ~n256 & n377 ;
  assign n379 = ~x29 & n378 ;
  assign n380 = ( ~n253 & n375 ) | ( ~n253 & n379 ) | ( n375 & n379 ) ;
  assign n381 = ( n247 & n263 ) | ( n247 & n380 ) | ( n263 & n380 ) ;
  assign n382 = x18 & ~n381 ;
  assign n383 = ( x18 & n380 ) | ( x18 & ~n382 ) | ( n380 & ~n382 ) ;
  assign n384 = ( ~x29 & x75 ) | ( ~x29 & n253 ) | ( x75 & n253 ) ;
  assign n385 = ~x32 & x76 ;
  assign n386 = ( x50 & n256 ) | ( x50 & n385 ) | ( n256 & n385 ) ;
  assign n387 = ~n256 & n386 ;
  assign n388 = ~x29 & n387 ;
  assign n389 = ( ~n253 & n384 ) | ( ~n253 & n388 ) | ( n384 & n388 ) ;
  assign n390 = ( n247 & n263 ) | ( n247 & n389 ) | ( n263 & n389 ) ;
  assign n391 = x19 & ~n390 ;
  assign n392 = ( x19 & n389 ) | ( x19 & ~n391 ) | ( n389 & ~n391 ) ;
  assign n393 = ( ~x29 & x76 ) | ( ~x29 & n253 ) | ( x76 & n253 ) ;
  assign n394 = ~x32 & x77 ;
  assign n395 = ( x50 & n256 ) | ( x50 & n394 ) | ( n256 & n394 ) ;
  assign n396 = ~n256 & n395 ;
  assign n397 = ~x29 & n396 ;
  assign n398 = ( ~n253 & n393 ) | ( ~n253 & n397 ) | ( n393 & n397 ) ;
  assign n399 = ( n247 & n263 ) | ( n247 & n398 ) | ( n263 & n398 ) ;
  assign n400 = x20 & ~n399 ;
  assign n401 = ( x20 & n398 ) | ( x20 & ~n400 ) | ( n398 & ~n400 ) ;
  assign n402 = ( ~x29 & x77 ) | ( ~x29 & n253 ) | ( x77 & n253 ) ;
  assign n403 = ~x32 & x78 ;
  assign n404 = ( x50 & n256 ) | ( x50 & n403 ) | ( n256 & n403 ) ;
  assign n405 = ~n256 & n404 ;
  assign n406 = ~x29 & n405 ;
  assign n407 = ( ~n253 & n402 ) | ( ~n253 & n406 ) | ( n402 & n406 ) ;
  assign n408 = ( n247 & n263 ) | ( n247 & n407 ) | ( n263 & n407 ) ;
  assign n409 = x21 & ~n408 ;
  assign n410 = ( x21 & n407 ) | ( x21 & ~n409 ) | ( n407 & ~n409 ) ;
  assign n411 = ( ~x29 & x78 ) | ( ~x29 & n253 ) | ( x78 & n253 ) ;
  assign n412 = ~x32 & x79 ;
  assign n413 = ( x50 & n256 ) | ( x50 & n412 ) | ( n256 & n412 ) ;
  assign n414 = ~n256 & n413 ;
  assign n415 = ~x29 & n414 ;
  assign n416 = ( ~n253 & n411 ) | ( ~n253 & n415 ) | ( n411 & n415 ) ;
  assign n417 = ( n247 & n263 ) | ( n247 & n416 ) | ( n263 & n416 ) ;
  assign n418 = x22 & ~n417 ;
  assign n419 = ( x22 & n416 ) | ( x22 & ~n418 ) | ( n416 & ~n418 ) ;
  assign n420 = ( ~x29 & x79 ) | ( ~x29 & n253 ) | ( x79 & n253 ) ;
  assign n421 = ~x32 & x80 ;
  assign n422 = ( x50 & n256 ) | ( x50 & n421 ) | ( n256 & n421 ) ;
  assign n423 = ~n256 & n422 ;
  assign n424 = ~x29 & n423 ;
  assign n425 = ( ~n253 & n420 ) | ( ~n253 & n424 ) | ( n420 & n424 ) ;
  assign n426 = ( n247 & n263 ) | ( n247 & n425 ) | ( n263 & n425 ) ;
  assign n427 = x23 & ~n426 ;
  assign n428 = ( x23 & n425 ) | ( x23 & ~n427 ) | ( n425 & ~n427 ) ;
  assign n429 = ( ~x29 & x80 ) | ( ~x29 & n253 ) | ( x80 & n253 ) ;
  assign n430 = ~x32 & x81 ;
  assign n431 = ( x50 & n256 ) | ( x50 & n430 ) | ( n256 & n430 ) ;
  assign n432 = ~n256 & n431 ;
  assign n433 = ~x29 & n432 ;
  assign n434 = ( ~n253 & n429 ) | ( ~n253 & n433 ) | ( n429 & n433 ) ;
  assign n435 = ( n247 & n263 ) | ( n247 & n434 ) | ( n263 & n434 ) ;
  assign n436 = x24 & ~n435 ;
  assign n437 = ( x24 & n434 ) | ( x24 & ~n436 ) | ( n434 & ~n436 ) ;
  assign n438 = x27 & n263 ;
  assign n439 = ( x25 & n113 ) | ( x25 & n438 ) | ( n113 & n438 ) ;
  assign n440 = ~n113 & n439 ;
  assign n441 = ( x29 & n253 ) | ( x29 & ~n440 ) | ( n253 & ~n440 ) ;
  assign n442 = x81 & n441 ;
  assign n443 = ( x81 & n440 ) | ( x81 & ~n442 ) | ( n440 & ~n442 ) ;
  assign n444 = x1 & ~x40 ;
  assign n445 = ( ~x48 & x92 ) | ( ~x48 & n444 ) | ( x92 & n444 ) ;
  assign n446 = x82 & ~n445 ;
  assign n447 = ( x48 & ~x82 ) | ( x48 & n445 ) | ( ~x82 & n445 ) ;
  assign n448 = ( ~x48 & n446 ) | ( ~x48 & n447 ) | ( n446 & n447 ) ;
  assign n449 = x92 | n444 ;
  assign n450 = ( ~x48 & x83 ) | ( ~x48 & x84 ) | ( x83 & x84 ) ;
  assign n451 = ~x48 & x82 ;
  assign n452 = ( ~x84 & n450 ) | ( ~x84 & n451 ) | ( n450 & n451 ) ;
  assign n453 = ( x83 & n449 ) | ( x83 & n452 ) | ( n449 & n452 ) ;
  assign n454 = ( x82 & n449 ) | ( x82 & ~n452 ) | ( n449 & ~n452 ) ;
  assign n455 = n453 & ~n454 ;
  assign n456 = ( ~x83 & n453 ) | ( ~x83 & n455 ) | ( n453 & n455 ) ;
  assign n457 = ( x48 & ~x82 ) | ( x48 & x83 ) | ( ~x82 & x83 ) ;
  assign n458 = n450 & ~n457 ;
  assign n459 = ( x84 & n449 ) | ( x84 & n458 ) | ( n449 & n458 ) ;
  assign n460 = ( x83 & n449 ) | ( x83 & ~n458 ) | ( n449 & ~n458 ) ;
  assign n461 = n459 & ~n460 ;
  assign n462 = ( ~x84 & n459 ) | ( ~x84 & n461 ) | ( n459 & n461 ) ;
  assign n463 = ( ~x48 & x50 ) | ( ~x48 & n176 ) | ( x50 & n176 ) ;
  assign n464 = x85 & ~n463 ;
  assign n465 = ( x48 & ~x85 ) | ( x48 & n463 ) | ( ~x85 & n463 ) ;
  assign n466 = ( ~x48 & n464 ) | ( ~x48 & n465 ) | ( n464 & n465 ) ;
  assign n467 = x82 & n174 ;
  assign n468 = x49 | x50 ;
  assign n469 = ( n174 & ~n467 ) | ( n174 & n468 ) | ( ~n467 & n468 ) ;
  assign n470 = x85 & n469 ;
  assign n471 = x86 & ~n470 ;
  assign n472 = x50 | n176 ;
  assign n473 = ~x86 & n472 ;
  assign n474 = n471 | n473 ;
  assign n475 = ~x48 & n474 ;
  assign n476 = ( x85 & n179 ) | ( x85 & n475 ) | ( n179 & n475 ) ;
  assign n477 = x85 & x86 ;
  assign n478 = x87 & ~n477 ;
  assign n479 = x86 & n469 ;
  assign n480 = x85 & n479 ;
  assign n481 = x87 & ~n480 ;
  assign n482 = ~x87 & n472 ;
  assign n483 = n481 | n482 ;
  assign n484 = ~x48 & n483 ;
  assign n485 = ( n477 & n478 ) | ( n477 & n484 ) | ( n478 & n484 ) ;
  assign n486 = ( x86 & x87 ) | ( x86 & x88 ) | ( x87 & x88 ) ;
  assign n487 = x85 & ~n486 ;
  assign n488 = ( x85 & x88 ) | ( x85 & ~n487 ) | ( x88 & ~n487 ) ;
  assign n489 = x88 & n477 ;
  assign n490 = ( x87 & ~n469 ) | ( x87 & n489 ) | ( ~n469 & n489 ) ;
  assign n491 = n469 & n490 ;
  assign n492 = ( x50 & x88 ) | ( x50 & ~n491 ) | ( x88 & ~n491 ) ;
  assign n493 = ~n176 & n492 ;
  assign n494 = ( n176 & ~n491 ) | ( n176 & n493 ) | ( ~n491 & n493 ) ;
  assign n495 = n488 & n494 ;
  assign n496 = ~x48 & n495 ;
  assign n497 = x87 & x89 ;
  assign n498 = ( x88 & ~n469 ) | ( x88 & n497 ) | ( ~n469 & n497 ) ;
  assign n499 = n469 & n498 ;
  assign n500 = ~n477 & n499 ;
  assign n501 = ( ~x50 & x89 ) | ( ~x50 & n176 ) | ( x89 & n176 ) ;
  assign n502 = x87 & n489 ;
  assign n503 = x89 | n502 ;
  assign n504 = ( x50 & n501 ) | ( x50 & n503 ) | ( n501 & n503 ) ;
  assign n505 = ~x48 & n504 ;
  assign n506 = ( ~n499 & n500 ) | ( ~n499 & n505 ) | ( n500 & n505 ) ;
  assign n507 = ( ~x29 & x47 ) | ( ~x29 & n229 ) | ( x47 & n229 ) ;
  assign n508 = ( x29 & ~x59 ) | ( x29 & n229 ) | ( ~x59 & n229 ) ;
  assign n509 = n507 & ~n508 ;
  assign n510 = ( x48 & x57 ) | ( x48 & x90 ) | ( x57 & x90 ) ;
  assign n511 = ~x91 & n510 ;
  assign n512 = ( x48 & x91 ) | ( x48 & ~n510 ) | ( x91 & ~n510 ) ;
  assign n513 = ( ~x48 & n511 ) | ( ~x48 & n512 ) | ( n511 & n512 ) ;
  assign n514 = n174 & ~n444 ;
  assign n515 = ~x82 & n514 ;
  assign n516 = ~x29 & n449 ;
  assign n517 = ~n515 & n516 ;
  assign n518 = ( x26 & x93 ) | ( x26 & ~n221 ) | ( x93 & ~n221 ) ;
  assign n519 = x89 & n99 ;
  assign n520 = ~x86 & n519 ;
  assign n521 = x50 & n520 ;
  assign n522 = ( x85 & x87 ) | ( x85 & n521 ) | ( x87 & n521 ) ;
  assign n523 = ~x87 & n522 ;
  assign n524 = ~n221 & n523 ;
  assign n525 = ( ~x26 & n518 ) | ( ~x26 & n524 ) | ( n518 & n524 ) ;
  assign y0 = ~x51 ;
  assign y1 = ~x52 ;
  assign y2 = ~x53 ;
  assign y3 = ~x54 ;
  assign y4 = ~x55 ;
  assign y5 = ~x56 ;
  assign y6 = n110 ;
  assign y7 = n120 ;
  assign y8 = n127 ;
  assign y9 = n132 ;
  assign y10 = n140 ;
  assign y11 = n142 ;
  assign y12 = n144 ;
  assign y13 = n146 ;
  assign y14 = n148 ;
  assign y15 = n150 ;
  assign y16 = n152 ;
  assign y17 = n153 ;
  assign y18 = n154 ;
  assign y19 = n155 ;
  assign y20 = n156 ;
  assign y21 = n157 ;
  assign y22 = n158 ;
  assign y23 = n159 ;
  assign y24 = n160 ;
  assign y25 = n169 ;
  assign y26 = n173 ;
  assign y27 = n178 ;
  assign y28 = n189 ;
  assign y29 = n194 ;
  assign y30 = n199 ;
  assign y31 = n204 ;
  assign y32 = n209 ;
  assign y33 = n214 ;
  assign y34 = n216 ;
  assign y35 = n223 ;
  assign y36 = n243 ;
  assign y37 = n250 ;
  assign y38 = n266 ;
  assign y39 = n275 ;
  assign y40 = n284 ;
  assign y41 = n293 ;
  assign y42 = n302 ;
  assign y43 = n311 ;
  assign y44 = n320 ;
  assign y45 = n329 ;
  assign y46 = n338 ;
  assign y47 = n347 ;
  assign y48 = n356 ;
  assign y49 = n365 ;
  assign y50 = n374 ;
  assign y51 = n383 ;
  assign y52 = n392 ;
  assign y53 = n401 ;
  assign y54 = n410 ;
  assign y55 = n419 ;
  assign y56 = n428 ;
  assign y57 = n437 ;
  assign y58 = n443 ;
  assign y59 = n448 ;
  assign y60 = n456 ;
  assign y61 = n462 ;
  assign y62 = n466 ;
  assign y63 = n476 ;
  assign y64 = n485 ;
  assign y65 = n496 ;
  assign y66 = n506 ;
  assign y67 = n509 ;
  assign y68 = n513 ;
  assign y69 = n517 ;
  assign y70 = n525 ;
endmodule
