module top( N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 , N223 , N329 , N370 , N421 , N430 , N431 , N432 );
  input N1 , N102 , N105 , N108 , N11 , N112 , N115 , N14 , N17 , N21 , N24 , N27 , N30 , N34 , N37 , N4 , N40 , N43 , N47 , N50 , N53 , N56 , N60 , N63 , N66 , N69 , N73 , N76 , N79 , N8 , N82 , N86 , N89 , N92 , N95 , N99 ;
  output N223 , N329 , N370 , N421 , N430 , N431 , N432 ;
  wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 ;
  assign n37 = ~N24 & N30 ;
  assign n38 = ~N102 & N108 ;
  assign n39 = n37 | n38 ;
  assign n40 = ~N1 & N4 ;
  assign n41 = ~N89 & N95 ;
  assign n42 = ~N76 & N82 ;
  assign n43 = n41 | n42 ;
  assign n44 = n40 | n43 ;
  assign n45 = ~N63 & N69 ;
  assign n46 = ~N37 & N43 ;
  assign n47 = n45 | n46 ;
  assign n48 = ~N50 & N56 ;
  assign n49 = ~N11 & N17 ;
  assign n50 = n48 | n49 ;
  assign n51 = n47 | n50 ;
  assign n52 = n44 | n51 ;
  assign n53 = n39 | n52 ;
  assign n54 = N102 & n53 ;
  assign n55 = N108 & ~n54 ;
  assign n56 = ~N112 & n55 ;
  assign n57 = N76 & n53 ;
  assign n58 = N82 & ~n57 ;
  assign n59 = ~N86 & n58 ;
  assign n60 = n56 | n59 ;
  assign n61 = N30 & ~n53 ;
  assign n62 = n37 | n61 ;
  assign n63 = ~N34 & n62 ;
  assign n64 = N11 & n53 ;
  assign n65 = N17 & ~n64 ;
  assign n66 = ~N21 & n65 ;
  assign n67 = n63 | n66 ;
  assign n68 = n60 | n67 ;
  assign n69 = N1 & n53 ;
  assign n70 = N4 & ~n69 ;
  assign n71 = ~N8 & n70 ;
  assign n72 = N89 & n53 ;
  assign n73 = N95 & ~n72 ;
  assign n74 = ~N99 & n73 ;
  assign n75 = n71 | n74 ;
  assign n76 = N50 & n53 ;
  assign n77 = N56 & ~n76 ;
  assign n78 = ~N60 & n77 ;
  assign n79 = N69 & ~n53 ;
  assign n80 = n45 | n79 ;
  assign n81 = ~N73 & n80 ;
  assign n82 = N37 & n53 ;
  assign n83 = N43 & ~n82 ;
  assign n84 = ~N47 & n83 ;
  assign n85 = n81 | n84 ;
  assign n86 = n78 | n85 ;
  assign n87 = n75 | n86 ;
  assign n88 = n68 | n87 ;
  assign n89 = N34 & n88 ;
  assign n90 = n62 & ~n89 ;
  assign n91 = ~N40 & n90 ;
  assign n92 = N99 & n88 ;
  assign n93 = n73 & ~n92 ;
  assign n94 = ~N105 & n93 ;
  assign n95 = N21 & n88 ;
  assign n96 = n65 & ~n95 ;
  assign n97 = ~N27 & n96 ;
  assign n98 = n94 | n97 ;
  assign n99 = n91 | n98 ;
  assign n100 = N8 & n88 ;
  assign n101 = n70 & ~n100 ;
  assign n102 = ~N14 & n101 ;
  assign n103 = N86 & n88 ;
  assign n104 = n58 & ~n103 ;
  assign n105 = ~N92 & n104 ;
  assign n106 = n102 | n105 ;
  assign n107 = N73 & n88 ;
  assign n108 = n80 & ~n107 ;
  assign n109 = ~N79 & n108 ;
  assign n110 = N60 & n88 ;
  assign n111 = n77 & ~n110 ;
  assign n112 = ~N66 & n111 ;
  assign n113 = n109 | n112 ;
  assign n114 = N47 & n88 ;
  assign n115 = n83 & ~n114 ;
  assign n116 = ~N53 & n115 ;
  assign n117 = N112 & n88 ;
  assign n118 = n55 & ~n117 ;
  assign n119 = ~N115 & n118 ;
  assign n120 = n116 | n119 ;
  assign n121 = n113 | n120 ;
  assign n122 = n106 | n121 ;
  assign n123 = n99 | n122 ;
  assign n124 = N40 & n123 ;
  assign n125 = n90 & ~n124 ;
  assign n126 = N27 & n123 ;
  assign n127 = n96 & ~n126 ;
  assign n128 = n125 | n127 ;
  assign n129 = N53 & n123 ;
  assign n130 = n115 & ~n129 ;
  assign n131 = n111 & ~n123 ;
  assign n132 = n112 | n131 ;
  assign n133 = n130 | n132 ;
  assign n134 = n128 | n133 ;
  assign n135 = N92 & n123 ;
  assign n136 = n104 & ~n135 ;
  assign n137 = N79 & n123 ;
  assign n138 = n108 & ~n137 ;
  assign n139 = n136 | n138 ;
  assign n140 = N105 & n123 ;
  assign n141 = n93 & ~n140 ;
  assign n142 = N115 & n123 ;
  assign n143 = n118 & ~n142 ;
  assign n144 = n141 | n143 ;
  assign n145 = n139 | n144 ;
  assign n146 = n134 | n145 ;
  assign n147 = N14 & n123 ;
  assign n148 = n101 & ~n147 ;
  assign n149 = n146 & ~n148 ;
  assign n150 = ~n133 & n139 ;
  assign n151 = n128 | n150 ;
  assign n152 = ~n133 & n138 ;
  assign n153 = ~n136 & n141 ;
  assign n154 = n130 | n153 ;
  assign n155 = n152 | n154 ;
  assign n156 = ~n125 & n155 ;
  assign n157 = n127 | n156 ;
  assign N223 = n53 ;
  assign N329 = n88 ;
  assign N370 = n123 ;
  assign N421 = n149 ;
  assign N430 = n134 ;
  assign N431 = n151 ;
  assign N432 = n157 ;
endmodule
