module top(x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476;
  assign n129 = x64 ^ x0;
  assign n131 = x65 ^ x1;
  assign n130 = x0 & x64;
  assign n132 = n131 ^ n130;
  assign n133 = n130 ^ x65;
  assign n134 = n131 & ~n133;
  assign n135 = n134 ^ x1;
  assign n136 = n135 ^ x2;
  assign n137 = n136 ^ x66;
  assign n138 = x66 ^ x2;
  assign n139 = n135 ^ x66;
  assign n140 = n138 & ~n139;
  assign n141 = n140 ^ x2;
  assign n142 = n141 ^ x67;
  assign n143 = n142 ^ x3;
  assign n144 = x67 ^ x3;
  assign n145 = ~n142 & n144;
  assign n146 = n145 ^ x3;
  assign n147 = n146 ^ x4;
  assign n148 = n147 ^ x68;
  assign n149 = x68 ^ x4;
  assign n150 = n146 ^ x68;
  assign n151 = n149 & ~n150;
  assign n152 = n151 ^ x4;
  assign n153 = n152 ^ x5;
  assign n154 = n153 ^ x69;
  assign n155 = x69 ^ x5;
  assign n156 = n152 ^ x69;
  assign n157 = n155 & ~n156;
  assign n158 = n157 ^ x5;
  assign n159 = n158 ^ x6;
  assign n160 = n159 ^ x70;
  assign n161 = x70 ^ x6;
  assign n162 = n158 ^ x70;
  assign n163 = n161 & ~n162;
  assign n164 = n163 ^ x6;
  assign n165 = n164 ^ x7;
  assign n166 = n165 ^ x71;
  assign n167 = x71 ^ x7;
  assign n168 = n164 ^ x71;
  assign n169 = n167 & ~n168;
  assign n170 = n169 ^ x7;
  assign n171 = n170 ^ x8;
  assign n172 = n171 ^ x72;
  assign n173 = x72 ^ x8;
  assign n174 = n170 ^ x72;
  assign n175 = n173 & ~n174;
  assign n176 = n175 ^ x8;
  assign n177 = n176 ^ x9;
  assign n178 = n177 ^ x73;
  assign n179 = x73 ^ x9;
  assign n180 = n176 ^ x73;
  assign n181 = n179 & ~n180;
  assign n182 = n181 ^ x9;
  assign n183 = n182 ^ x10;
  assign n184 = n183 ^ x74;
  assign n185 = x74 ^ x10;
  assign n186 = n182 ^ x74;
  assign n187 = n185 & ~n186;
  assign n188 = n187 ^ x10;
  assign n189 = n188 ^ x11;
  assign n190 = n189 ^ x75;
  assign n191 = x75 ^ x11;
  assign n192 = n188 ^ x75;
  assign n193 = n191 & ~n192;
  assign n194 = n193 ^ x11;
  assign n195 = n194 ^ x12;
  assign n196 = n195 ^ x76;
  assign n197 = x76 ^ x12;
  assign n198 = n194 ^ x76;
  assign n199 = n197 & ~n198;
  assign n200 = n199 ^ x12;
  assign n201 = n200 ^ x13;
  assign n202 = n201 ^ x77;
  assign n203 = x77 ^ x13;
  assign n204 = n200 ^ x77;
  assign n205 = n203 & ~n204;
  assign n206 = n205 ^ x13;
  assign n207 = n206 ^ x14;
  assign n208 = n207 ^ x78;
  assign n209 = x78 ^ x14;
  assign n210 = n206 ^ x78;
  assign n211 = n209 & ~n210;
  assign n212 = n211 ^ x14;
  assign n213 = n212 ^ x15;
  assign n214 = n213 ^ x79;
  assign n215 = x79 ^ x15;
  assign n216 = n212 ^ x79;
  assign n217 = n215 & ~n216;
  assign n218 = n217 ^ x15;
  assign n219 = n218 ^ x80;
  assign n220 = n219 ^ x16;
  assign n221 = x80 ^ x16;
  assign n222 = ~n219 & n221;
  assign n223 = n222 ^ x16;
  assign n224 = n223 ^ x17;
  assign n225 = n224 ^ x81;
  assign n226 = x81 ^ x17;
  assign n227 = n223 ^ x81;
  assign n228 = n226 & ~n227;
  assign n229 = n228 ^ x17;
  assign n230 = n229 ^ x82;
  assign n231 = n230 ^ x18;
  assign n232 = x82 ^ x18;
  assign n233 = ~n230 & n232;
  assign n234 = n233 ^ x18;
  assign n235 = n234 ^ x19;
  assign n236 = n235 ^ x83;
  assign n237 = x83 ^ x19;
  assign n238 = n234 ^ x83;
  assign n239 = n237 & ~n238;
  assign n240 = n239 ^ x19;
  assign n241 = n240 ^ x20;
  assign n242 = n241 ^ x84;
  assign n243 = x84 ^ x20;
  assign n244 = n240 ^ x84;
  assign n245 = n243 & ~n244;
  assign n246 = n245 ^ x20;
  assign n247 = n246 ^ x21;
  assign n248 = n247 ^ x85;
  assign n249 = x85 ^ x21;
  assign n250 = n246 ^ x85;
  assign n251 = n249 & ~n250;
  assign n252 = n251 ^ x21;
  assign n253 = n252 ^ x22;
  assign n254 = n253 ^ x86;
  assign n255 = x86 ^ x22;
  assign n256 = n252 ^ x86;
  assign n257 = n255 & ~n256;
  assign n258 = n257 ^ x22;
  assign n259 = n258 ^ x87;
  assign n260 = n259 ^ x23;
  assign n261 = x87 ^ x23;
  assign n262 = ~n259 & n261;
  assign n263 = n262 ^ x23;
  assign n264 = n263 ^ x88;
  assign n265 = n264 ^ x24;
  assign n266 = x88 ^ x24;
  assign n267 = ~n264 & n266;
  assign n268 = n267 ^ x24;
  assign n269 = n268 ^ x25;
  assign n270 = n269 ^ x89;
  assign n271 = x89 ^ x25;
  assign n272 = n268 ^ x89;
  assign n273 = n271 & ~n272;
  assign n274 = n273 ^ x25;
  assign n275 = n274 ^ x26;
  assign n276 = n275 ^ x90;
  assign n277 = x90 ^ x26;
  assign n278 = n274 ^ x90;
  assign n279 = n277 & ~n278;
  assign n280 = n279 ^ x26;
  assign n281 = n280 ^ x27;
  assign n282 = n281 ^ x91;
  assign n283 = x91 ^ x27;
  assign n284 = n280 ^ x91;
  assign n285 = n283 & ~n284;
  assign n286 = n285 ^ x27;
  assign n287 = n286 ^ x28;
  assign n288 = n287 ^ x92;
  assign n289 = x92 ^ x28;
  assign n290 = n286 ^ x92;
  assign n291 = n289 & ~n290;
  assign n292 = n291 ^ x28;
  assign n293 = n292 ^ x93;
  assign n294 = n293 ^ x29;
  assign n295 = x93 ^ x29;
  assign n296 = ~n293 & n295;
  assign n297 = n296 ^ x29;
  assign n298 = n297 ^ x30;
  assign n299 = n298 ^ x94;
  assign n300 = x94 ^ x30;
  assign n301 = n297 ^ x94;
  assign n302 = n300 & ~n301;
  assign n303 = n302 ^ x30;
  assign n304 = n303 ^ x31;
  assign n305 = n304 ^ x95;
  assign n310 = x96 ^ x32;
  assign n306 = x95 ^ x31;
  assign n307 = n303 ^ x95;
  assign n308 = n306 & ~n307;
  assign n309 = n308 ^ x31;
  assign n311 = n310 ^ n309;
  assign n312 = n309 ^ x96;
  assign n313 = n310 & ~n312;
  assign n314 = n313 ^ x32;
  assign n315 = n314 ^ x97;
  assign n316 = n315 ^ x33;
  assign n320 = x98 ^ x34;
  assign n317 = x97 ^ x33;
  assign n318 = ~n315 & n317;
  assign n319 = n318 ^ x33;
  assign n321 = n320 ^ n319;
  assign n323 = n319 ^ x98;
  assign n324 = n320 & ~n323;
  assign n325 = n324 ^ x34;
  assign n322 = x99 ^ x35;
  assign n326 = n325 ^ n322;
  assign n327 = n325 ^ x99;
  assign n328 = n322 & ~n327;
  assign n329 = n328 ^ x35;
  assign n330 = n329 ^ x100;
  assign n331 = n330 ^ x36;
  assign n335 = x101 ^ x37;
  assign n332 = x100 ^ x36;
  assign n333 = ~n330 & n332;
  assign n334 = n333 ^ x36;
  assign n336 = n335 ^ n334;
  assign n337 = n334 ^ x101;
  assign n338 = n335 & ~n337;
  assign n339 = n338 ^ x37;
  assign n340 = n339 ^ x38;
  assign n341 = n340 ^ x102;
  assign n342 = x102 ^ x38;
  assign n343 = n339 ^ x102;
  assign n344 = n342 & ~n343;
  assign n345 = n344 ^ x38;
  assign n346 = n345 ^ x39;
  assign n347 = n346 ^ x103;
  assign n348 = x103 ^ x39;
  assign n349 = n345 ^ x103;
  assign n350 = n348 & ~n349;
  assign n351 = n350 ^ x39;
  assign n352 = n351 ^ x104;
  assign n353 = n352 ^ x40;
  assign n354 = x104 ^ x40;
  assign n355 = ~n352 & n354;
  assign n356 = n355 ^ x40;
  assign n357 = n356 ^ x41;
  assign n358 = n357 ^ x105;
  assign n359 = x105 ^ x41;
  assign n360 = n356 ^ x105;
  assign n361 = n359 & ~n360;
  assign n362 = n361 ^ x41;
  assign n363 = n362 ^ x106;
  assign n364 = n363 ^ x42;
  assign n365 = x106 ^ x42;
  assign n366 = ~n363 & n365;
  assign n367 = n366 ^ x42;
  assign n368 = n367 ^ x43;
  assign n369 = n368 ^ x107;
  assign n370 = x107 ^ x43;
  assign n371 = n367 ^ x107;
  assign n372 = n370 & ~n371;
  assign n373 = n372 ^ x43;
  assign n374 = n373 ^ x108;
  assign n375 = n374 ^ x44;
  assign n376 = x108 ^ x44;
  assign n377 = ~n374 & n376;
  assign n378 = n377 ^ x44;
  assign n379 = n378 ^ x109;
  assign n380 = n379 ^ x45;
  assign n381 = x109 ^ x45;
  assign n382 = ~n379 & n381;
  assign n383 = n382 ^ x45;
  assign n384 = n383 ^ x46;
  assign n385 = n384 ^ x110;
  assign n386 = x110 ^ x46;
  assign n387 = n383 ^ x110;
  assign n388 = n386 & ~n387;
  assign n389 = n388 ^ x46;
  assign n390 = n389 ^ x47;
  assign n391 = n390 ^ x111;
  assign n393 = x111 ^ x47;
  assign n394 = n389 ^ x111;
  assign n395 = n393 & ~n394;
  assign n396 = n395 ^ x47;
  assign n392 = x112 ^ x48;
  assign n397 = n396 ^ n392;
  assign n399 = n396 ^ x112;
  assign n400 = n392 & ~n399;
  assign n401 = n400 ^ x48;
  assign n398 = x113 ^ x49;
  assign n402 = n401 ^ n398;
  assign n404 = n401 ^ x113;
  assign n405 = n398 & ~n404;
  assign n406 = n405 ^ x49;
  assign n403 = x114 ^ x50;
  assign n407 = n406 ^ n403;
  assign n411 = x115 ^ x51;
  assign n408 = n406 ^ x114;
  assign n409 = n403 & ~n408;
  assign n410 = n409 ^ x50;
  assign n412 = n411 ^ n410;
  assign n414 = n410 ^ x115;
  assign n415 = n411 & ~n414;
  assign n416 = n415 ^ x51;
  assign n413 = x116 ^ x52;
  assign n417 = n416 ^ n413;
  assign n419 = n416 ^ x116;
  assign n420 = n413 & ~n419;
  assign n421 = n420 ^ x52;
  assign n418 = x117 ^ x53;
  assign n422 = n421 ^ n418;
  assign n424 = n421 ^ x117;
  assign n425 = n418 & ~n424;
  assign n426 = n425 ^ x53;
  assign n423 = x118 ^ x54;
  assign n427 = n426 ^ n423;
  assign n431 = x119 ^ x55;
  assign n428 = n426 ^ x118;
  assign n429 = n423 & ~n428;
  assign n430 = n429 ^ x54;
  assign n432 = n431 ^ n430;
  assign n434 = n430 ^ x119;
  assign n435 = n431 & ~n434;
  assign n436 = n435 ^ x55;
  assign n433 = x120 ^ x56;
  assign n437 = n436 ^ n433;
  assign n438 = n436 ^ x120;
  assign n439 = n433 & ~n438;
  assign n440 = n439 ^ x56;
  assign n441 = n440 ^ x57;
  assign n442 = n441 ^ x121;
  assign n444 = x121 ^ x57;
  assign n445 = n440 ^ x121;
  assign n446 = n444 & ~n445;
  assign n447 = n446 ^ x57;
  assign n443 = x122 ^ x58;
  assign n448 = n447 ^ n443;
  assign n452 = x123 ^ x59;
  assign n449 = n447 ^ x122;
  assign n450 = n443 & ~n449;
  assign n451 = n450 ^ x58;
  assign n453 = n452 ^ n451;
  assign n455 = n451 ^ x123;
  assign n456 = n452 & ~n455;
  assign n457 = n456 ^ x59;
  assign n454 = x124 ^ x60;
  assign n458 = n457 ^ n454;
  assign n460 = n457 ^ x124;
  assign n461 = n454 & ~n460;
  assign n462 = n461 ^ x60;
  assign n459 = x125 ^ x61;
  assign n463 = n462 ^ n459;
  assign n465 = n462 ^ x125;
  assign n466 = n459 & ~n465;
  assign n467 = n466 ^ x61;
  assign n464 = x126 ^ x62;
  assign n468 = n467 ^ n464;
  assign n470 = n467 ^ x126;
  assign n471 = n464 & ~n470;
  assign n472 = n471 ^ x62;
  assign n469 = x127 ^ x63;
  assign n473 = n472 ^ n469;
  assign n474 = n472 ^ x127;
  assign n475 = n469 & ~n474;
  assign n476 = n475 ^ x63;
  assign y0 = n129;
  assign y1 = n132;
  assign y2 = n137;
  assign y3 = n143;
  assign y4 = n148;
  assign y5 = n154;
  assign y6 = n160;
  assign y7 = n166;
  assign y8 = n172;
  assign y9 = n178;
  assign y10 = n184;
  assign y11 = n190;
  assign y12 = n196;
  assign y13 = n202;
  assign y14 = n208;
  assign y15 = n214;
  assign y16 = n220;
  assign y17 = n225;
  assign y18 = n231;
  assign y19 = n236;
  assign y20 = n242;
  assign y21 = n248;
  assign y22 = n254;
  assign y23 = n260;
  assign y24 = n265;
  assign y25 = n270;
  assign y26 = n276;
  assign y27 = n282;
  assign y28 = n288;
  assign y29 = n294;
  assign y30 = n299;
  assign y31 = n305;
  assign y32 = n311;
  assign y33 = n316;
  assign y34 = n321;
  assign y35 = n326;
  assign y36 = n331;
  assign y37 = n336;
  assign y38 = n341;
  assign y39 = n347;
  assign y40 = n353;
  assign y41 = n358;
  assign y42 = n364;
  assign y43 = n369;
  assign y44 = n375;
  assign y45 = n380;
  assign y46 = n385;
  assign y47 = n391;
  assign y48 = n397;
  assign y49 = n402;
  assign y50 = n407;
  assign y51 = n412;
  assign y52 = n417;
  assign y53 = n422;
  assign y54 = n427;
  assign y55 = n432;
  assign y56 = n437;
  assign y57 = n442;
  assign y58 = n448;
  assign y59 = n453;
  assign y60 = n458;
  assign y61 = n463;
  assign y62 = n468;
  assign y63 = n473;
  assign y64 = n476;
endmodule
