module top(x0, x1, x2, x3, x4, x5, x6, x7, y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239, y240, y241, y242, y243, y244, y245, y246, y247, y248, y249, y250, y251, y252, y253, y254, y255);
  input x0, x1, x2, x3, x4, x5, x6, x7;
  output y0, y1, y2, y3, y4, y5, y6, y7, y8, y9, y10, y11, y12, y13, y14, y15, y16, y17, y18, y19, y20, y21, y22, y23, y24, y25, y26, y27, y28, y29, y30, y31, y32, y33, y34, y35, y36, y37, y38, y39, y40, y41, y42, y43, y44, y45, y46, y47, y48, y49, y50, y51, y52, y53, y54, y55, y56, y57, y58, y59, y60, y61, y62, y63, y64, y65, y66, y67, y68, y69, y70, y71, y72, y73, y74, y75, y76, y77, y78, y79, y80, y81, y82, y83, y84, y85, y86, y87, y88, y89, y90, y91, y92, y93, y94, y95, y96, y97, y98, y99, y100, y101, y102, y103, y104, y105, y106, y107, y108, y109, y110, y111, y112, y113, y114, y115, y116, y117, y118, y119, y120, y121, y122, y123, y124, y125, y126, y127, y128, y129, y130, y131, y132, y133, y134, y135, y136, y137, y138, y139, y140, y141, y142, y143, y144, y145, y146, y147, y148, y149, y150, y151, y152, y153, y154, y155, y156, y157, y158, y159, y160, y161, y162, y163, y164, y165, y166, y167, y168, y169, y170, y171, y172, y173, y174, y175, y176, y177, y178, y179, y180, y181, y182, y183, y184, y185, y186, y187, y188, y189, y190, y191, y192, y193, y194, y195, y196, y197, y198, y199, y200, y201, y202, y203, y204, y205, y206, y207, y208, y209, y210, y211, y212, y213, y214, y215, y216, y217, y218, y219, y220, y221, y222, y223, y224, y225, y226, y227, y228, y229, y230, y231, y232, y233, y234, y235, y236, y237, y238, y239, y240, y241, y242, y243, y244, y245, y246, y247, y248, y249, y250, y251, y252, y253, y254, y255;
  wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349;
  assign n9 = ~x6 & x7;
  assign n10 = ~x2 & ~x3;
  assign n11 = n9 & n10;
  assign n12 = ~x4 & ~x5;
  assign n13 = ~x0 & ~x1;
  assign n14 = n12 & n13;
  assign n15 = n11 & n14;
  assign n16 = n9 & n12;
  assign n17 = x0 & ~x1;
  assign n18 = n10 & n17;
  assign n19 = n16 & n18;
  assign n20 = ~x0 & x1;
  assign n21 = n10 & n20;
  assign n22 = n16 & n21;
  assign n23 = x0 & x1;
  assign n24 = n10 & n23;
  assign n25 = n16 & n24;
  assign n26 = x2 & ~x3;
  assign n27 = n13 & n26;
  assign n28 = n16 & n27;
  assign n29 = n17 & n26;
  assign n30 = n16 & n29;
  assign n31 = n20 & n26;
  assign n32 = n16 & n31;
  assign n33 = n23 & n26;
  assign n34 = n16 & n33;
  assign n35 = ~x2 & x3;
  assign n36 = n13 & n35;
  assign n37 = n16 & n36;
  assign n38 = n17 & n35;
  assign n39 = n16 & n38;
  assign n40 = n20 & n35;
  assign n41 = n16 & n40;
  assign n42 = n23 & n35;
  assign n43 = n16 & n42;
  assign n44 = x2 & x3;
  assign n45 = n13 & n44;
  assign n46 = n16 & n45;
  assign n47 = n17 & n44;
  assign n48 = n16 & n47;
  assign n49 = n20 & n44;
  assign n50 = n16 & n49;
  assign n51 = n23 & n44;
  assign n52 = n16 & n51;
  assign n53 = ~x5 & ~x6;
  assign n54 = n10 & n53;
  assign n55 = x4 & x7;
  assign n56 = n13 & n55;
  assign n57 = n54 & n56;
  assign n58 = n17 & n55;
  assign n59 = n54 & n58;
  assign n60 = n20 & n55;
  assign n61 = n54 & n60;
  assign n62 = n23 & n55;
  assign n63 = n54 & n62;
  assign n64 = n26 & n53;
  assign n65 = n56 & n64;
  assign n66 = n58 & n64;
  assign n67 = n60 & n64;
  assign n68 = n62 & n64;
  assign n69 = n35 & n53;
  assign n70 = n56 & n69;
  assign n71 = n58 & n69;
  assign n72 = n60 & n69;
  assign n73 = n62 & n69;
  assign n74 = n44 & n53;
  assign n75 = n56 & n74;
  assign n76 = n58 & n74;
  assign n77 = n60 & n74;
  assign n78 = n62 & n74;
  assign n79 = ~x4 & x5;
  assign n80 = n13 & n79;
  assign n81 = n11 & n80;
  assign n82 = n9 & n17;
  assign n83 = n10 & n79;
  assign n84 = n82 & n83;
  assign n85 = n9 & n20;
  assign n86 = n83 & n85;
  assign n87 = n9 & n23;
  assign n88 = n83 & n87;
  assign n89 = n9 & n13;
  assign n90 = n26 & n79;
  assign n91 = n89 & n90;
  assign n92 = n82 & n90;
  assign n93 = n85 & n90;
  assign n94 = n87 & n90;
  assign n95 = n35 & n79;
  assign n96 = n89 & n95;
  assign n97 = n82 & n95;
  assign n98 = n85 & n95;
  assign n99 = n87 & n95;
  assign n100 = n44 & n79;
  assign n101 = n89 & n100;
  assign n102 = n82 & n100;
  assign n103 = n85 & n100;
  assign n104 = n87 & n100;
  assign n105 = x4 & x5;
  assign n106 = n10 & n105;
  assign n107 = n89 & n106;
  assign n108 = n82 & n106;
  assign n109 = n85 & n106;
  assign n110 = n87 & n106;
  assign n111 = n26 & n105;
  assign n112 = n89 & n111;
  assign n113 = n82 & n111;
  assign n114 = n85 & n111;
  assign n115 = n87 & n111;
  assign n116 = n35 & n105;
  assign n117 = n89 & n116;
  assign n118 = n82 & n116;
  assign n119 = n85 & n116;
  assign n120 = n87 & n116;
  assign n121 = n44 & n105;
  assign n122 = n89 & n121;
  assign n123 = n82 & n121;
  assign n124 = n85 & n121;
  assign n125 = n87 & n121;
  assign n126 = x6 & x7;
  assign n127 = n10 & n126;
  assign n128 = n14 & n127;
  assign n129 = n12 & n17;
  assign n130 = n127 & n129;
  assign n131 = n12 & n20;
  assign n132 = n127 & n131;
  assign n133 = n12 & n23;
  assign n134 = n127 & n133;
  assign n135 = n26 & n126;
  assign n136 = n14 & n135;
  assign n137 = n129 & n135;
  assign n138 = n131 & n135;
  assign n139 = n133 & n135;
  assign n140 = n35 & n126;
  assign n141 = n14 & n140;
  assign n142 = n129 & n140;
  assign n143 = n131 & n140;
  assign n144 = n133 & n140;
  assign n145 = n44 & n126;
  assign n146 = n14 & n145;
  assign n147 = n129 & n145;
  assign n148 = n131 & n145;
  assign n149 = n133 & n145;
  assign n150 = x4 & ~x5;
  assign n151 = n13 & n150;
  assign n152 = n127 & n151;
  assign n153 = n17 & n150;
  assign n154 = n127 & n153;
  assign n155 = n20 & n150;
  assign n156 = n127 & n155;
  assign n157 = n23 & n150;
  assign n158 = n127 & n157;
  assign n159 = n135 & n151;
  assign n160 = n135 & n153;
  assign n161 = n135 & n155;
  assign n162 = n135 & n157;
  assign n163 = n140 & n151;
  assign n164 = n140 & n153;
  assign n165 = n140 & n155;
  assign n166 = n140 & n157;
  assign n167 = n145 & n151;
  assign n168 = n145 & n153;
  assign n169 = n145 & n155;
  assign n170 = n145 & n157;
  assign n171 = n80 & n127;
  assign n172 = n17 & n126;
  assign n173 = n83 & n172;
  assign n174 = n20 & n126;
  assign n175 = n83 & n174;
  assign n176 = n23 & n126;
  assign n177 = n83 & n176;
  assign n178 = n80 & n135;
  assign n179 = n90 & n172;
  assign n180 = n90 & n174;
  assign n181 = n90 & n176;
  assign n182 = n80 & n140;
  assign n183 = n95 & n172;
  assign n184 = n95 & n174;
  assign n185 = n95 & n176;
  assign n186 = n80 & n145;
  assign n187 = n100 & n172;
  assign n188 = n100 & n174;
  assign n189 = n100 & n176;
  assign n190 = n10 & n13;
  assign n191 = n105 & n126;
  assign n192 = n190 & n191;
  assign n193 = n18 & n191;
  assign n194 = n21 & n191;
  assign n195 = n24 & n191;
  assign n196 = n27 & n191;
  assign n197 = n29 & n191;
  assign n198 = n31 & n191;
  assign n199 = n111 & n176;
  assign n200 = n36 & n191;
  assign n201 = n38 & n191;
  assign n202 = n116 & n174;
  assign n203 = n42 & n191;
  assign n204 = n45 & n191;
  assign n205 = n47 & n191;
  assign n206 = n49 & n191;
  assign n207 = n51 & n191;
  assign n208 = ~x6 & ~x7;
  assign n209 = n12 & n208;
  assign n210 = n190 & n209;
  assign n211 = n18 & n209;
  assign n212 = n21 & n209;
  assign n213 = n24 & n209;
  assign n214 = n27 & n209;
  assign n215 = n29 & n209;
  assign n216 = n31 & n209;
  assign n217 = n33 & n209;
  assign n218 = n36 & n209;
  assign n219 = n38 & n209;
  assign n220 = n40 & n209;
  assign n221 = n42 & n209;
  assign n222 = n45 & n209;
  assign n223 = n47 & n209;
  assign n224 = n49 & n209;
  assign n225 = n51 & n209;
  assign n226 = x4 & ~x7;
  assign n227 = n13 & n226;
  assign n228 = n54 & n227;
  assign n229 = n17 & n226;
  assign n230 = n54 & n229;
  assign n231 = n20 & n226;
  assign n232 = n54 & n231;
  assign n233 = n23 & n226;
  assign n234 = n54 & n233;
  assign n235 = n64 & n227;
  assign n236 = n64 & n229;
  assign n237 = n64 & n231;
  assign n238 = n64 & n233;
  assign n239 = n69 & n227;
  assign n240 = n69 & n229;
  assign n241 = n69 & n231;
  assign n242 = n69 & n233;
  assign n243 = n74 & n227;
  assign n244 = n74 & n229;
  assign n245 = n74 & n231;
  assign n246 = n74 & n233;
  assign n247 = n79 & n208;
  assign n248 = n190 & n247;
  assign n249 = n18 & n247;
  assign n250 = n21 & n247;
  assign n251 = n24 & n247;
  assign n252 = n27 & n247;
  assign n253 = n29 & n247;
  assign n254 = n31 & n247;
  assign n255 = n33 & n247;
  assign n256 = n36 & n247;
  assign n257 = n38 & n247;
  assign n258 = n40 & n247;
  assign n259 = n42 & n247;
  assign n260 = n45 & n247;
  assign n261 = n47 & n247;
  assign n262 = n49 & n247;
  assign n263 = n51 & n247;
  assign n264 = n105 & n208;
  assign n265 = n190 & n264;
  assign n266 = n18 & n264;
  assign n267 = n21 & n264;
  assign n268 = n24 & n264;
  assign n269 = n27 & n264;
  assign n270 = n29 & n264;
  assign n271 = n31 & n264;
  assign n272 = n33 & n264;
  assign n273 = n36 & n264;
  assign n274 = n38 & n264;
  assign n275 = n40 & n264;
  assign n276 = n42 & n264;
  assign n277 = n45 & n264;
  assign n278 = n47 & n264;
  assign n279 = n49 & n264;
  assign n280 = n51 & n264;
  assign n281 = x6 & ~x7;
  assign n282 = n12 & n281;
  assign n283 = n190 & n282;
  assign n284 = n18 & n282;
  assign n285 = n21 & n282;
  assign n286 = n24 & n282;
  assign n287 = n27 & n282;
  assign n288 = n29 & n282;
  assign n289 = n31 & n282;
  assign n290 = n33 & n282;
  assign n291 = n36 & n282;
  assign n292 = n38 & n282;
  assign n293 = n40 & n282;
  assign n294 = n42 & n282;
  assign n295 = n45 & n282;
  assign n296 = n47 & n282;
  assign n297 = n49 & n282;
  assign n298 = n51 & n282;
  assign n299 = n150 & n281;
  assign n300 = n190 & n299;
  assign n301 = n18 & n299;
  assign n302 = n21 & n299;
  assign n303 = n24 & n299;
  assign n304 = n27 & n299;
  assign n305 = n29 & n299;
  assign n306 = n31 & n299;
  assign n307 = n33 & n299;
  assign n308 = n36 & n299;
  assign n309 = n38 & n299;
  assign n310 = n40 & n299;
  assign n311 = n42 & n299;
  assign n312 = n45 & n299;
  assign n313 = n47 & n299;
  assign n314 = n49 & n299;
  assign n315 = n51 & n299;
  assign n316 = n79 & n281;
  assign n317 = n190 & n316;
  assign n318 = n18 & n316;
  assign n319 = n21 & n316;
  assign n320 = n24 & n316;
  assign n321 = n27 & n316;
  assign n322 = n29 & n316;
  assign n323 = n31 & n316;
  assign n324 = n33 & n316;
  assign n325 = n36 & n316;
  assign n326 = n38 & n316;
  assign n327 = n40 & n316;
  assign n328 = n42 & n316;
  assign n329 = n45 & n316;
  assign n330 = n47 & n316;
  assign n331 = n49 & n316;
  assign n332 = n51 & n316;
  assign n333 = n105 & n281;
  assign n334 = n190 & n333;
  assign n335 = n18 & n333;
  assign n336 = n21 & n333;
  assign n337 = n24 & n333;
  assign n338 = n27 & n333;
  assign n339 = n29 & n333;
  assign n340 = n31 & n333;
  assign n341 = n33 & n333;
  assign n342 = n36 & n333;
  assign n343 = n38 & n333;
  assign n344 = n40 & n333;
  assign n345 = n42 & n333;
  assign n346 = n45 & n333;
  assign n347 = n47 & n333;
  assign n348 = n49 & n333;
  assign n349 = n51 & n333;
  assign y0 = n15;
  assign y1 = n19;
  assign y2 = n22;
  assign y3 = n25;
  assign y4 = n28;
  assign y5 = n30;
  assign y6 = n32;
  assign y7 = n34;
  assign y8 = n37;
  assign y9 = n39;
  assign y10 = n41;
  assign y11 = n43;
  assign y12 = n46;
  assign y13 = n48;
  assign y14 = n50;
  assign y15 = n52;
  assign y16 = n57;
  assign y17 = n59;
  assign y18 = n61;
  assign y19 = n63;
  assign y20 = n65;
  assign y21 = n66;
  assign y22 = n67;
  assign y23 = n68;
  assign y24 = n70;
  assign y25 = n71;
  assign y26 = n72;
  assign y27 = n73;
  assign y28 = n75;
  assign y29 = n76;
  assign y30 = n77;
  assign y31 = n78;
  assign y32 = n81;
  assign y33 = n84;
  assign y34 = n86;
  assign y35 = n88;
  assign y36 = n91;
  assign y37 = n92;
  assign y38 = n93;
  assign y39 = n94;
  assign y40 = n96;
  assign y41 = n97;
  assign y42 = n98;
  assign y43 = n99;
  assign y44 = n101;
  assign y45 = n102;
  assign y46 = n103;
  assign y47 = n104;
  assign y48 = n107;
  assign y49 = n108;
  assign y50 = n109;
  assign y51 = n110;
  assign y52 = n112;
  assign y53 = n113;
  assign y54 = n114;
  assign y55 = n115;
  assign y56 = n117;
  assign y57 = n118;
  assign y58 = n119;
  assign y59 = n120;
  assign y60 = n122;
  assign y61 = n123;
  assign y62 = n124;
  assign y63 = n125;
  assign y64 = n128;
  assign y65 = n130;
  assign y66 = n132;
  assign y67 = n134;
  assign y68 = n136;
  assign y69 = n137;
  assign y70 = n138;
  assign y71 = n139;
  assign y72 = n141;
  assign y73 = n142;
  assign y74 = n143;
  assign y75 = n144;
  assign y76 = n146;
  assign y77 = n147;
  assign y78 = n148;
  assign y79 = n149;
  assign y80 = n152;
  assign y81 = n154;
  assign y82 = n156;
  assign y83 = n158;
  assign y84 = n159;
  assign y85 = n160;
  assign y86 = n161;
  assign y87 = n162;
  assign y88 = n163;
  assign y89 = n164;
  assign y90 = n165;
  assign y91 = n166;
  assign y92 = n167;
  assign y93 = n168;
  assign y94 = n169;
  assign y95 = n170;
  assign y96 = n171;
  assign y97 = n173;
  assign y98 = n175;
  assign y99 = n177;
  assign y100 = n178;
  assign y101 = n179;
  assign y102 = n180;
  assign y103 = n181;
  assign y104 = n182;
  assign y105 = n183;
  assign y106 = n184;
  assign y107 = n185;
  assign y108 = n186;
  assign y109 = n187;
  assign y110 = n188;
  assign y111 = n189;
  assign y112 = n192;
  assign y113 = n193;
  assign y114 = n194;
  assign y115 = n195;
  assign y116 = n196;
  assign y117 = n197;
  assign y118 = n198;
  assign y119 = n199;
  assign y120 = n200;
  assign y121 = n201;
  assign y122 = n202;
  assign y123 = n203;
  assign y124 = n204;
  assign y125 = n205;
  assign y126 = n206;
  assign y127 = n207;
  assign y128 = n210;
  assign y129 = n211;
  assign y130 = n212;
  assign y131 = n213;
  assign y132 = n214;
  assign y133 = n215;
  assign y134 = n216;
  assign y135 = n217;
  assign y136 = n218;
  assign y137 = n219;
  assign y138 = n220;
  assign y139 = n221;
  assign y140 = n222;
  assign y141 = n223;
  assign y142 = n224;
  assign y143 = n225;
  assign y144 = n228;
  assign y145 = n230;
  assign y146 = n232;
  assign y147 = n234;
  assign y148 = n235;
  assign y149 = n236;
  assign y150 = n237;
  assign y151 = n238;
  assign y152 = n239;
  assign y153 = n240;
  assign y154 = n241;
  assign y155 = n242;
  assign y156 = n243;
  assign y157 = n244;
  assign y158 = n245;
  assign y159 = n246;
  assign y160 = n248;
  assign y161 = n249;
  assign y162 = n250;
  assign y163 = n251;
  assign y164 = n252;
  assign y165 = n253;
  assign y166 = n254;
  assign y167 = n255;
  assign y168 = n256;
  assign y169 = n257;
  assign y170 = n258;
  assign y171 = n259;
  assign y172 = n260;
  assign y173 = n261;
  assign y174 = n262;
  assign y175 = n263;
  assign y176 = n265;
  assign y177 = n266;
  assign y178 = n267;
  assign y179 = n268;
  assign y180 = n269;
  assign y181 = n270;
  assign y182 = n271;
  assign y183 = n272;
  assign y184 = n273;
  assign y185 = n274;
  assign y186 = n275;
  assign y187 = n276;
  assign y188 = n277;
  assign y189 = n278;
  assign y190 = n279;
  assign y191 = n280;
  assign y192 = n283;
  assign y193 = n284;
  assign y194 = n285;
  assign y195 = n286;
  assign y196 = n287;
  assign y197 = n288;
  assign y198 = n289;
  assign y199 = n290;
  assign y200 = n291;
  assign y201 = n292;
  assign y202 = n293;
  assign y203 = n294;
  assign y204 = n295;
  assign y205 = n296;
  assign y206 = n297;
  assign y207 = n298;
  assign y208 = n300;
  assign y209 = n301;
  assign y210 = n302;
  assign y211 = n303;
  assign y212 = n304;
  assign y213 = n305;
  assign y214 = n306;
  assign y215 = n307;
  assign y216 = n308;
  assign y217 = n309;
  assign y218 = n310;
  assign y219 = n311;
  assign y220 = n312;
  assign y221 = n313;
  assign y222 = n314;
  assign y223 = n315;
  assign y224 = n317;
  assign y225 = n318;
  assign y226 = n319;
  assign y227 = n320;
  assign y228 = n321;
  assign y229 = n322;
  assign y230 = n323;
  assign y231 = n324;
  assign y232 = n325;
  assign y233 = n326;
  assign y234 = n327;
  assign y235 = n328;
  assign y236 = n329;
  assign y237 = n330;
  assign y238 = n331;
  assign y239 = n332;
  assign y240 = n334;
  assign y241 = n335;
  assign y242 = n336;
  assign y243 = n337;
  assign y244 = n338;
  assign y245 = n339;
  assign y246 = n340;
  assign y247 = n341;
  assign y248 = n342;
  assign y249 = n343;
  assign y250 = n344;
  assign y251 = n345;
  assign y252 = n346;
  assign y253 = n347;
  assign y254 = n348;
  assign y255 = n349;
endmodule
