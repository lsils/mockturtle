module top( N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 , N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 );
  input N1 , N101 , N105 , N109 , N113 , N117 , N121 , N125 , N129 , N13 , N130 , N131 , N132 , N133 , N134 , N135 , N136 , N137 , N17 , N21 , N25 , N29 , N33 , N37 , N41 , N45 , N49 , N5 , N53 , N57 , N61 , N65 , N69 , N73 , N77 , N81 , N85 , N89 , N9 , N93 , N97 ;
  output N724 , N725 , N726 , N727 , N728 , N729 , N730 , N731 , N732 , N733 , N734 , N735 , N736 , N737 , N738 , N739 , N740 , N741 , N742 , N743 , N744 , N745 , N746 , N747 , N748 , N749 , N750 , N751 , N752 , N753 , N754 , N755 ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 ;
  assign n42 = N33 & ~N49 ;
  assign n43 = ~N33 & N49 ;
  assign n44 = n42 | n43 ;
  assign n45 = N129 & N137 ;
  assign n46 = N1 & ~N17 ;
  assign n47 = ~N1 & N17 ;
  assign n48 = n46 | n47 ;
  assign n49 = n45 & ~n48 ;
  assign n50 = ~n45 & n48 ;
  assign n51 = n49 | n50 ;
  assign n52 = n44 | n51 ;
  assign n53 = n44 & n51 ;
  assign n54 = n52 & ~n53 ;
  assign n55 = N73 | N77 ;
  assign n56 = N73 & N77 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = N65 & ~N69 ;
  assign n59 = ~N65 & N69 ;
  assign n60 = n58 | n59 ;
  assign n61 = ~n57 & n60 ;
  assign n62 = n57 & ~n60 ;
  assign n63 = n61 | n62 ;
  assign n64 = N89 | N93 ;
  assign n65 = N89 & N93 ;
  assign n66 = n64 & ~n65 ;
  assign n67 = N81 & ~N85 ;
  assign n68 = ~N81 & N85 ;
  assign n69 = n67 | n68 ;
  assign n70 = ~n66 & n69 ;
  assign n71 = n66 & ~n69 ;
  assign n72 = n70 | n71 ;
  assign n73 = n63 & n72 ;
  assign n74 = n63 | n72 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = ~n54 & n75 ;
  assign n77 = n54 & ~n75 ;
  assign n78 = n76 | n77 ;
  assign n79 = N135 & N137 ;
  assign n80 = N105 & ~N121 ;
  assign n81 = ~N105 & N121 ;
  assign n82 = n80 | n81 ;
  assign n83 = N73 & ~N89 ;
  assign n84 = ~N73 & N89 ;
  assign n85 = n83 | n84 ;
  assign n86 = ~n82 & n85 ;
  assign n87 = n82 & ~n85 ;
  assign n88 = n86 | n87 ;
  assign n89 = n79 & n88 ;
  assign n90 = n79 | n88 ;
  assign n91 = ~n89 & n90 ;
  assign n92 = N13 | N9 ;
  assign n93 = N13 & N9 ;
  assign n94 = n92 & ~n93 ;
  assign n95 = N1 & ~N5 ;
  assign n96 = ~N1 & N5 ;
  assign n97 = n95 | n96 ;
  assign n98 = ~n94 & n97 ;
  assign n99 = n94 & ~n97 ;
  assign n100 = n98 | n99 ;
  assign n101 = N41 | N45 ;
  assign n102 = N41 & N45 ;
  assign n103 = n101 & ~n102 ;
  assign n104 = N33 & ~N37 ;
  assign n105 = ~N33 & N37 ;
  assign n106 = n104 | n105 ;
  assign n107 = ~n103 & n106 ;
  assign n108 = n103 & ~n106 ;
  assign n109 = n107 | n108 ;
  assign n110 = n100 & n109 ;
  assign n111 = n100 | n109 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = ~n91 & n112 ;
  assign n114 = n91 & ~n112 ;
  assign n115 = n113 | n114 ;
  assign n116 = N136 & N137 ;
  assign n117 = N109 & ~N125 ;
  assign n118 = ~N109 & N125 ;
  assign n119 = n117 | n118 ;
  assign n120 = N77 & ~N93 ;
  assign n121 = ~N77 & N93 ;
  assign n122 = n120 | n121 ;
  assign n123 = ~n119 & n122 ;
  assign n124 = n119 & ~n122 ;
  assign n125 = n123 | n124 ;
  assign n126 = n116 & n125 ;
  assign n127 = n116 | n125 ;
  assign n128 = ~n126 & n127 ;
  assign n129 = N25 | N29 ;
  assign n130 = N25 & N29 ;
  assign n131 = n129 & ~n130 ;
  assign n132 = N17 & ~N21 ;
  assign n133 = ~N17 & N21 ;
  assign n134 = n132 | n133 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = n131 & ~n134 ;
  assign n137 = n135 | n136 ;
  assign n138 = N57 | N61 ;
  assign n139 = N57 & N61 ;
  assign n140 = n138 & ~n139 ;
  assign n141 = N49 & ~N53 ;
  assign n142 = ~N49 & N53 ;
  assign n143 = n141 | n142 ;
  assign n144 = ~n140 & n143 ;
  assign n145 = n140 & ~n143 ;
  assign n146 = n144 | n145 ;
  assign n147 = n137 & n146 ;
  assign n148 = n137 | n146 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = ~n128 & n149 ;
  assign n151 = n128 & ~n149 ;
  assign n152 = n150 | n151 ;
  assign n153 = n115 & ~n152 ;
  assign n154 = N131 & N137 ;
  assign n155 = N41 & ~N57 ;
  assign n156 = ~N41 & N57 ;
  assign n157 = n155 | n156 ;
  assign n158 = ~N25 & N9 ;
  assign n159 = N25 & ~N9 ;
  assign n160 = n158 | n159 ;
  assign n161 = ~n157 & n160 ;
  assign n162 = n157 & ~n160 ;
  assign n163 = n161 | n162 ;
  assign n164 = n154 & n163 ;
  assign n165 = n154 | n163 ;
  assign n166 = ~n164 & n165 ;
  assign n167 = N105 | N109 ;
  assign n168 = N105 & N109 ;
  assign n169 = n167 & ~n168 ;
  assign n170 = ~N101 & N97 ;
  assign n171 = N101 & ~N97 ;
  assign n172 = n170 | n171 ;
  assign n173 = ~n169 & n172 ;
  assign n174 = n169 & ~n172 ;
  assign n175 = n173 | n174 ;
  assign n176 = n63 & n175 ;
  assign n177 = n63 | n175 ;
  assign n178 = ~n176 & n177 ;
  assign n179 = ~n166 & n178 ;
  assign n180 = n166 & ~n178 ;
  assign n181 = n179 | n180 ;
  assign n182 = N37 & ~N53 ;
  assign n183 = ~N37 & N53 ;
  assign n184 = n182 | n183 ;
  assign n185 = N130 & N137 ;
  assign n186 = ~N21 & N5 ;
  assign n187 = N21 & ~N5 ;
  assign n188 = n186 | n187 ;
  assign n189 = n185 & ~n188 ;
  assign n190 = ~n185 & n188 ;
  assign n191 = n189 | n190 ;
  assign n192 = n184 | n191 ;
  assign n193 = n184 & n191 ;
  assign n194 = n192 & ~n193 ;
  assign n195 = N121 | N125 ;
  assign n196 = N121 & N125 ;
  assign n197 = n195 & ~n196 ;
  assign n198 = N113 & ~N117 ;
  assign n199 = ~N113 & N117 ;
  assign n200 = n198 | n199 ;
  assign n201 = ~n197 & n200 ;
  assign n202 = n197 & ~n200 ;
  assign n203 = n201 | n202 ;
  assign n204 = n175 & n203 ;
  assign n205 = n175 | n203 ;
  assign n206 = ~n204 & n205 ;
  assign n207 = ~n194 & n206 ;
  assign n208 = n194 & ~n206 ;
  assign n209 = n207 | n208 ;
  assign n210 = ~n78 & n209 ;
  assign n211 = ~n181 & n210 ;
  assign n212 = n78 & ~n209 ;
  assign n213 = ~n181 & n212 ;
  assign n214 = n211 | n213 ;
  assign n215 = N132 & N137 ;
  assign n216 = N45 & ~N61 ;
  assign n217 = ~N45 & N61 ;
  assign n218 = n216 | n217 ;
  assign n219 = N13 & ~N29 ;
  assign n220 = ~N13 & N29 ;
  assign n221 = n219 | n220 ;
  assign n222 = ~n218 & n221 ;
  assign n223 = n218 & ~n221 ;
  assign n224 = n222 | n223 ;
  assign n225 = n215 & n224 ;
  assign n226 = n215 | n224 ;
  assign n227 = ~n225 & n226 ;
  assign n228 = n72 & n203 ;
  assign n229 = n72 | n203 ;
  assign n230 = ~n228 & n229 ;
  assign n231 = ~n227 & n230 ;
  assign n232 = n227 & ~n230 ;
  assign n233 = n231 | n232 ;
  assign n234 = n214 & ~n233 ;
  assign n235 = n181 & ~n233 ;
  assign n236 = ~n181 & n233 ;
  assign n237 = n235 | n236 ;
  assign n238 = n78 | n209 ;
  assign n239 = n237 & ~n238 ;
  assign n240 = n234 | n239 ;
  assign n241 = ~N113 & N97 ;
  assign n242 = N113 & ~N97 ;
  assign n243 = n241 | n242 ;
  assign n244 = N133 & N137 ;
  assign n245 = N65 & ~N81 ;
  assign n246 = ~N65 & N81 ;
  assign n247 = n245 | n246 ;
  assign n248 = n244 & ~n247 ;
  assign n249 = ~n244 & n247 ;
  assign n250 = n248 | n249 ;
  assign n251 = n243 | n250 ;
  assign n252 = n243 & n250 ;
  assign n253 = n251 & ~n252 ;
  assign n254 = n100 & n137 ;
  assign n255 = n100 | n137 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = ~n253 & n256 ;
  assign n258 = n253 & ~n256 ;
  assign n259 = n257 | n258 ;
  assign n260 = N101 & ~N117 ;
  assign n261 = ~N101 & N117 ;
  assign n262 = n260 | n261 ;
  assign n263 = N134 & N137 ;
  assign n264 = N69 & ~N85 ;
  assign n265 = ~N69 & N85 ;
  assign n266 = n264 | n265 ;
  assign n267 = n263 & ~n266 ;
  assign n268 = ~n263 & n266 ;
  assign n269 = n267 | n268 ;
  assign n270 = n262 | n269 ;
  assign n271 = n262 & n269 ;
  assign n272 = n270 & ~n271 ;
  assign n273 = n109 & n146 ;
  assign n274 = n109 | n146 ;
  assign n275 = ~n273 & n274 ;
  assign n276 = ~n272 & n275 ;
  assign n277 = n272 & ~n275 ;
  assign n278 = n276 | n277 ;
  assign n279 = n259 & ~n278 ;
  assign n280 = n240 & n279 ;
  assign n281 = n153 & n280 ;
  assign n282 = n78 & n281 ;
  assign n283 = N1 | n282 ;
  assign n284 = N1 & n282 ;
  assign n285 = n283 & ~n284 ;
  assign n286 = n209 & n281 ;
  assign n287 = N5 | n286 ;
  assign n288 = N5 & n286 ;
  assign n289 = n287 & ~n288 ;
  assign n290 = n181 & n281 ;
  assign n291 = N9 & n290 ;
  assign n292 = N9 | n290 ;
  assign n293 = ~n291 & n292 ;
  assign n294 = n233 & n281 ;
  assign n295 = ~N13 & n294 ;
  assign n296 = N13 & ~n294 ;
  assign n297 = n295 | n296 ;
  assign n298 = ~n115 & n152 ;
  assign n299 = n280 & n298 ;
  assign n300 = n78 & n299 ;
  assign n301 = N17 | n300 ;
  assign n302 = N17 & n300 ;
  assign n303 = n301 & ~n302 ;
  assign n304 = n209 & n299 ;
  assign n305 = N21 | n304 ;
  assign n306 = N21 & n304 ;
  assign n307 = n305 & ~n306 ;
  assign n308 = n181 & n299 ;
  assign n309 = N25 & n308 ;
  assign n310 = N25 | n308 ;
  assign n311 = ~n309 & n310 ;
  assign n312 = n233 & n299 ;
  assign n313 = ~N29 & n312 ;
  assign n314 = N29 & ~n312 ;
  assign n315 = n313 | n314 ;
  assign n316 = ~n259 & n278 ;
  assign n317 = n240 & n316 ;
  assign n318 = n153 & n317 ;
  assign n319 = n78 & n318 ;
  assign n320 = N33 | n319 ;
  assign n321 = N33 & n319 ;
  assign n322 = n320 & ~n321 ;
  assign n323 = n209 & n318 ;
  assign n324 = N37 | n323 ;
  assign n325 = N37 & n323 ;
  assign n326 = n324 & ~n325 ;
  assign n327 = n181 & n318 ;
  assign n328 = N41 & n327 ;
  assign n329 = N41 | n327 ;
  assign n330 = ~n328 & n329 ;
  assign n331 = n233 & n318 ;
  assign n332 = N45 | n331 ;
  assign n333 = N45 & n331 ;
  assign n334 = n332 & ~n333 ;
  assign n335 = n298 & n317 ;
  assign n336 = n78 & n335 ;
  assign n337 = N49 | n336 ;
  assign n338 = N49 & n336 ;
  assign n339 = n337 & ~n338 ;
  assign n340 = n209 & n335 ;
  assign n341 = N53 | n340 ;
  assign n342 = N53 & n340 ;
  assign n343 = n341 & ~n342 ;
  assign n344 = n181 & n335 ;
  assign n345 = N57 & n344 ;
  assign n346 = N57 | n344 ;
  assign n347 = ~n345 & n346 ;
  assign n348 = n233 & n335 ;
  assign n349 = N61 & n348 ;
  assign n350 = N61 | n348 ;
  assign n351 = ~n349 & n350 ;
  assign n352 = n279 | n316 ;
  assign n353 = n115 | n152 ;
  assign n354 = n352 & ~n353 ;
  assign n355 = n153 | n298 ;
  assign n356 = n259 | n278 ;
  assign n357 = n355 & ~n356 ;
  assign n358 = n354 | n357 ;
  assign n359 = n235 & n358 ;
  assign n360 = n212 & n359 ;
  assign n361 = n259 & n360 ;
  assign n362 = N65 | n361 ;
  assign n363 = N65 & n361 ;
  assign n364 = n362 & ~n363 ;
  assign n365 = n278 & n360 ;
  assign n366 = N69 | n365 ;
  assign n367 = N69 & n365 ;
  assign n368 = n366 & ~n367 ;
  assign n369 = n115 & n360 ;
  assign n370 = ~N73 & n369 ;
  assign n371 = N73 & ~n369 ;
  assign n372 = n370 | n371 ;
  assign n373 = n152 & n360 ;
  assign n374 = N77 & n373 ;
  assign n375 = N77 | n373 ;
  assign n376 = ~n374 & n375 ;
  assign n377 = n233 & n358 ;
  assign n378 = n213 & n377 ;
  assign n379 = n259 & n378 ;
  assign n380 = N81 | n379 ;
  assign n381 = N81 & n379 ;
  assign n382 = n380 & ~n381 ;
  assign n383 = n278 & n378 ;
  assign n384 = N85 | n383 ;
  assign n385 = N85 & n383 ;
  assign n386 = n384 & ~n385 ;
  assign n387 = n115 & n378 ;
  assign n388 = N89 & n387 ;
  assign n389 = N89 | n387 ;
  assign n390 = ~n388 & n389 ;
  assign n391 = n152 & n378 ;
  assign n392 = N93 | n391 ;
  assign n393 = N93 & n391 ;
  assign n394 = n392 & ~n393 ;
  assign n395 = n210 & n359 ;
  assign n396 = n259 & n395 ;
  assign n397 = N97 | n396 ;
  assign n398 = N97 & n396 ;
  assign n399 = n397 & ~n398 ;
  assign n400 = n278 & n395 ;
  assign n401 = N101 | n400 ;
  assign n402 = N101 & n400 ;
  assign n403 = n401 & ~n402 ;
  assign n404 = n115 & n395 ;
  assign n405 = ~N105 & n404 ;
  assign n406 = N105 & ~n404 ;
  assign n407 = n405 | n406 ;
  assign n408 = n152 & n395 ;
  assign n409 = N109 & n408 ;
  assign n410 = N109 | n408 ;
  assign n411 = ~n409 & n410 ;
  assign n412 = n211 & n377 ;
  assign n413 = n259 & n412 ;
  assign n414 = N113 | n413 ;
  assign n415 = N113 & n413 ;
  assign n416 = n414 & ~n415 ;
  assign n417 = n278 & n412 ;
  assign n418 = N117 | n417 ;
  assign n419 = N117 & n417 ;
  assign n420 = n418 & ~n419 ;
  assign n421 = n115 & n412 ;
  assign n422 = N121 & n421 ;
  assign n423 = N121 | n421 ;
  assign n424 = ~n422 & n423 ;
  assign n425 = n152 & n412 ;
  assign n426 = N125 | n425 ;
  assign n427 = N125 & n425 ;
  assign n428 = n426 & ~n427 ;
  assign N724 = n285 ;
  assign N725 = n289 ;
  assign N726 = n293 ;
  assign N727 = n297 ;
  assign N728 = n303 ;
  assign N729 = n307 ;
  assign N730 = n311 ;
  assign N731 = n315 ;
  assign N732 = n322 ;
  assign N733 = n326 ;
  assign N734 = n330 ;
  assign N735 = n334 ;
  assign N736 = n339 ;
  assign N737 = n343 ;
  assign N738 = n347 ;
  assign N739 = n351 ;
  assign N740 = n364 ;
  assign N741 = n368 ;
  assign N742 = n372 ;
  assign N743 = n376 ;
  assign N744 = n382 ;
  assign N745 = n386 ;
  assign N746 = n390 ;
  assign N747 = n394 ;
  assign N748 = n399 ;
  assign N749 = n403 ;
  assign N750 = n407 ;
  assign N751 = n411 ;
  assign N752 = n416 ;
  assign N753 = n420 ;
  assign N754 = n424 ;
  assign N755 = n428 ;
endmodule
