module top( G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G5 , G6 , G7 , G8 , G9 , G1324 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1343 , G1344 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 );
  input G1 , G10 , G11 , G12 , G13 , G14 , G15 , G16 , G17 , G18 , G19 , G2 , G20 , G21 , G22 , G23 , G24 , G25 , G26 , G27 , G28 , G29 , G3 , G30 , G31 , G32 , G33 , G34 , G35 , G36 , G37 , G38 , G39 , G4 , G40 , G41 , G5 , G6 , G7 , G8 , G9 ;
  output G1324 , G1325 , G1326 , G1327 , G1328 , G1329 , G1330 , G1331 , G1332 , G1333 , G1334 , G1335 , G1336 , G1337 , G1338 , G1339 , G1340 , G1341 , G1342 , G1343 , G1344 , G1345 , G1346 , G1347 , G1348 , G1349 , G1350 , G1351 , G1352 , G1353 , G1354 , G1355 ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 ;
  assign n42 = G33 & G41 ;
  assign n43 = G17 | G19 ;
  assign n44 = G17 & G19 ;
  assign n45 = n43 & ~n44 ;
  assign n46 = ~G18 & G20 ;
  assign n47 = G18 & ~G20 ;
  assign n48 = n46 | n47 ;
  assign n49 = ~n45 & n48 ;
  assign n50 = n45 & ~n48 ;
  assign n51 = n49 | n50 ;
  assign n52 = ~n42 & n51 ;
  assign n53 = n42 & ~n51 ;
  assign n54 = n52 | n53 ;
  assign n55 = G22 | G23 ;
  assign n56 = G22 & G23 ;
  assign n57 = n55 & ~n56 ;
  assign n58 = G21 & ~G24 ;
  assign n59 = ~G21 & G24 ;
  assign n60 = n58 | n59 ;
  assign n61 = ~n57 & n60 ;
  assign n62 = n57 & ~n60 ;
  assign n63 = n61 | n62 ;
  assign n64 = G13 | G5 ;
  assign n65 = G13 & G5 ;
  assign n66 = n64 & ~n65 ;
  assign n67 = G1 & ~G9 ;
  assign n68 = ~G1 & G9 ;
  assign n69 = n67 | n68 ;
  assign n70 = n66 | n69 ;
  assign n71 = n66 & n69 ;
  assign n72 = n70 & ~n71 ;
  assign n73 = n63 & n72 ;
  assign n74 = n63 | n72 ;
  assign n75 = ~n73 & n74 ;
  assign n76 = ~n54 & n75 ;
  assign n77 = n54 & ~n75 ;
  assign n78 = n76 | n77 ;
  assign n79 = G3 | G4 ;
  assign n80 = G3 & G4 ;
  assign n81 = n79 & ~n80 ;
  assign n82 = G1 & ~G2 ;
  assign n83 = ~G1 & G2 ;
  assign n84 = n82 | n83 ;
  assign n85 = ~n81 & n84 ;
  assign n86 = n81 & ~n84 ;
  assign n87 = n85 | n86 ;
  assign n88 = G39 & G41 ;
  assign n89 = n87 & ~n88 ;
  assign n90 = ~n87 & n88 ;
  assign n91 = n89 | n90 ;
  assign n92 = G10 | G12 ;
  assign n93 = G10 & G12 ;
  assign n94 = n92 & ~n93 ;
  assign n95 = ~G11 & G9 ;
  assign n96 = G11 & ~G9 ;
  assign n97 = n95 | n96 ;
  assign n98 = ~n94 & n97 ;
  assign n99 = n94 & ~n97 ;
  assign n100 = n98 | n99 ;
  assign n101 = G19 | G23 ;
  assign n102 = G19 & G23 ;
  assign n103 = n101 & ~n102 ;
  assign n104 = G27 & ~G31 ;
  assign n105 = ~G27 & G31 ;
  assign n106 = n104 | n105 ;
  assign n107 = n103 | n106 ;
  assign n108 = n103 & n106 ;
  assign n109 = n107 & ~n108 ;
  assign n110 = n100 & n109 ;
  assign n111 = n100 | n109 ;
  assign n112 = ~n110 & n111 ;
  assign n113 = ~n91 & n112 ;
  assign n114 = n91 & ~n112 ;
  assign n115 = n113 | n114 ;
  assign n116 = G7 | G8 ;
  assign n117 = G7 & G8 ;
  assign n118 = n116 & ~n117 ;
  assign n119 = ~G5 & G6 ;
  assign n120 = G5 & ~G6 ;
  assign n121 = n119 | n120 ;
  assign n122 = ~n118 & n121 ;
  assign n123 = n118 & ~n121 ;
  assign n124 = n122 | n123 ;
  assign n125 = G40 & G41 ;
  assign n126 = n124 & ~n125 ;
  assign n127 = ~n124 & n125 ;
  assign n128 = n126 | n127 ;
  assign n129 = G14 | G16 ;
  assign n130 = G14 & G16 ;
  assign n131 = n129 & ~n130 ;
  assign n132 = G13 & ~G15 ;
  assign n133 = ~G13 & G15 ;
  assign n134 = n132 | n133 ;
  assign n135 = ~n131 & n134 ;
  assign n136 = n131 & ~n134 ;
  assign n137 = n135 | n136 ;
  assign n138 = G20 | G24 ;
  assign n139 = G20 & G24 ;
  assign n140 = n138 & ~n139 ;
  assign n141 = ~G28 & G32 ;
  assign n142 = G28 & ~G32 ;
  assign n143 = n141 | n142 ;
  assign n144 = n140 | n143 ;
  assign n145 = n140 & n143 ;
  assign n146 = n144 & ~n145 ;
  assign n147 = n137 & n146 ;
  assign n148 = n137 | n146 ;
  assign n149 = ~n147 & n148 ;
  assign n150 = ~n128 & n149 ;
  assign n151 = n128 & ~n149 ;
  assign n152 = n150 | n151 ;
  assign n153 = n115 & ~n152 ;
  assign n154 = G37 & G41 ;
  assign n155 = n87 & ~n154 ;
  assign n156 = ~n87 & n154 ;
  assign n157 = n155 | n156 ;
  assign n158 = G21 & ~G25 ;
  assign n159 = ~G21 & G25 ;
  assign n160 = n158 | n159 ;
  assign n161 = G17 | G29 ;
  assign n162 = G17 & G29 ;
  assign n163 = n161 & ~n162 ;
  assign n164 = n160 | n163 ;
  assign n165 = n160 & n163 ;
  assign n166 = n164 & ~n165 ;
  assign n167 = n124 & n166 ;
  assign n168 = n124 | n166 ;
  assign n169 = ~n167 & n168 ;
  assign n170 = ~n157 & n169 ;
  assign n171 = n157 & ~n169 ;
  assign n172 = n170 | n171 ;
  assign n173 = G38 & G41 ;
  assign n174 = n100 & ~n173 ;
  assign n175 = ~n100 & n173 ;
  assign n176 = n174 | n175 ;
  assign n177 = ~G18 & G26 ;
  assign n178 = G18 & ~G26 ;
  assign n179 = n177 | n178 ;
  assign n180 = G22 | G30 ;
  assign n181 = G22 & G30 ;
  assign n182 = n180 & ~n181 ;
  assign n183 = n179 | n182 ;
  assign n184 = n179 & n182 ;
  assign n185 = n183 & ~n184 ;
  assign n186 = n137 & n185 ;
  assign n187 = n137 | n185 ;
  assign n188 = ~n186 & n187 ;
  assign n189 = ~n176 & n188 ;
  assign n190 = n176 & ~n188 ;
  assign n191 = n189 | n190 ;
  assign n192 = n172 & ~n191 ;
  assign n193 = G34 & G41 ;
  assign n194 = G29 | G30 ;
  assign n195 = G29 & G30 ;
  assign n196 = n194 & ~n195 ;
  assign n197 = ~G31 & G32 ;
  assign n198 = G31 & ~G32 ;
  assign n199 = n197 | n198 ;
  assign n200 = ~n196 & n199 ;
  assign n201 = n196 & ~n199 ;
  assign n202 = n200 | n201 ;
  assign n203 = ~n193 & n202 ;
  assign n204 = n193 & ~n202 ;
  assign n205 = n203 | n204 ;
  assign n206 = G25 | G28 ;
  assign n207 = G25 & G28 ;
  assign n208 = n206 & ~n207 ;
  assign n209 = G26 & ~G27 ;
  assign n210 = ~G26 & G27 ;
  assign n211 = n209 | n210 ;
  assign n212 = ~n208 & n211 ;
  assign n213 = n208 & ~n211 ;
  assign n214 = n212 | n213 ;
  assign n215 = G14 | G2 ;
  assign n216 = G14 & G2 ;
  assign n217 = n215 & ~n216 ;
  assign n218 = G10 & ~G6 ;
  assign n219 = ~G10 & G6 ;
  assign n220 = n218 | n219 ;
  assign n221 = n217 | n220 ;
  assign n222 = n217 & n220 ;
  assign n223 = n221 & ~n222 ;
  assign n224 = n214 & n223 ;
  assign n225 = n214 | n223 ;
  assign n226 = ~n224 & n225 ;
  assign n227 = ~n205 & n226 ;
  assign n228 = n205 & ~n226 ;
  assign n229 = n227 | n228 ;
  assign n230 = ~n78 & n229 ;
  assign n231 = G35 & G41 ;
  assign n232 = n51 & ~n231 ;
  assign n233 = ~n51 & n231 ;
  assign n234 = n232 | n233 ;
  assign n235 = G11 & ~G15 ;
  assign n236 = ~G11 & G15 ;
  assign n237 = n235 | n236 ;
  assign n238 = G3 | G7 ;
  assign n239 = G3 & G7 ;
  assign n240 = n238 & ~n239 ;
  assign n241 = n237 | n240 ;
  assign n242 = n237 & n240 ;
  assign n243 = n241 & ~n242 ;
  assign n244 = n214 & n243 ;
  assign n245 = n214 | n243 ;
  assign n246 = ~n244 & n245 ;
  assign n247 = ~n234 & n246 ;
  assign n248 = n234 & ~n246 ;
  assign n249 = n247 | n248 ;
  assign n250 = n230 & ~n249 ;
  assign n251 = n78 & ~n229 ;
  assign n252 = ~n249 & n251 ;
  assign n253 = n250 | n252 ;
  assign n254 = G36 & G41 ;
  assign n255 = n63 & ~n254 ;
  assign n256 = ~n63 & n254 ;
  assign n257 = n255 | n256 ;
  assign n258 = G12 & ~G4 ;
  assign n259 = ~G12 & G4 ;
  assign n260 = n258 | n259 ;
  assign n261 = G16 | G8 ;
  assign n262 = G16 & G8 ;
  assign n263 = n261 & ~n262 ;
  assign n264 = n260 | n263 ;
  assign n265 = n260 & n263 ;
  assign n266 = n264 & ~n265 ;
  assign n267 = n202 & n266 ;
  assign n268 = n202 | n266 ;
  assign n269 = ~n267 & n268 ;
  assign n270 = ~n257 & n269 ;
  assign n271 = n257 & ~n269 ;
  assign n272 = n270 | n271 ;
  assign n273 = n253 & ~n272 ;
  assign n274 = n249 & ~n272 ;
  assign n275 = ~n249 & n272 ;
  assign n276 = n274 | n275 ;
  assign n277 = n78 | n229 ;
  assign n278 = n276 & ~n277 ;
  assign n279 = n273 | n278 ;
  assign n280 = n192 & n279 ;
  assign n281 = n153 & n280 ;
  assign n282 = n78 & n281 ;
  assign n283 = G1 & ~n282 ;
  assign n284 = ~G1 & n282 ;
  assign n285 = n283 | n284 ;
  assign n286 = n229 & n281 ;
  assign n287 = G2 & ~n286 ;
  assign n288 = ~G2 & n286 ;
  assign n289 = n287 | n288 ;
  assign n290 = n249 & n281 ;
  assign n291 = G3 & ~n290 ;
  assign n292 = ~G3 & n290 ;
  assign n293 = n291 | n292 ;
  assign n294 = n272 & n281 ;
  assign n295 = G4 & ~n294 ;
  assign n296 = ~G4 & n294 ;
  assign n297 = n295 | n296 ;
  assign n298 = ~n115 & n152 ;
  assign n299 = n280 & n298 ;
  assign n300 = n78 & n299 ;
  assign n301 = G5 & ~n300 ;
  assign n302 = ~G5 & n300 ;
  assign n303 = n301 | n302 ;
  assign n304 = n229 & n299 ;
  assign n305 = G6 & ~n304 ;
  assign n306 = ~G6 & n304 ;
  assign n307 = n305 | n306 ;
  assign n308 = n249 & n299 ;
  assign n309 = G7 & ~n308 ;
  assign n310 = ~G7 & n308 ;
  assign n311 = n309 | n310 ;
  assign n312 = n272 & n299 ;
  assign n313 = G8 & ~n312 ;
  assign n314 = ~G8 & n312 ;
  assign n315 = n313 | n314 ;
  assign n316 = ~n172 & n191 ;
  assign n317 = n153 & n279 ;
  assign n318 = n316 & n317 ;
  assign n319 = n78 & n318 ;
  assign n320 = G9 & ~n319 ;
  assign n321 = ~G9 & n319 ;
  assign n322 = n320 | n321 ;
  assign n323 = n229 & n318 ;
  assign n324 = G10 & ~n323 ;
  assign n325 = ~G10 & n323 ;
  assign n326 = n324 | n325 ;
  assign n327 = n249 & n318 ;
  assign n328 = G11 & ~n327 ;
  assign n329 = ~G11 & n327 ;
  assign n330 = n328 | n329 ;
  assign n331 = n272 & n318 ;
  assign n332 = G12 & ~n331 ;
  assign n333 = ~G12 & n331 ;
  assign n334 = n332 | n333 ;
  assign n335 = n298 & n316 ;
  assign n336 = n279 & n335 ;
  assign n337 = n78 & n336 ;
  assign n338 = G13 | n337 ;
  assign n339 = G13 & n337 ;
  assign n340 = n338 & ~n339 ;
  assign n341 = n229 & n336 ;
  assign n342 = G14 | n341 ;
  assign n343 = G14 & n341 ;
  assign n344 = n342 & ~n343 ;
  assign n345 = n249 & n336 ;
  assign n346 = G15 & ~n345 ;
  assign n347 = ~G15 & n345 ;
  assign n348 = n346 | n347 ;
  assign n349 = n272 & n336 ;
  assign n350 = G16 | n349 ;
  assign n351 = G16 & n349 ;
  assign n352 = n350 & ~n351 ;
  assign n353 = n192 | n316 ;
  assign n354 = n115 | n152 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = n153 | n298 ;
  assign n357 = n172 | n191 ;
  assign n358 = n356 & ~n357 ;
  assign n359 = n355 | n358 ;
  assign n360 = n274 & n359 ;
  assign n361 = n251 & n360 ;
  assign n362 = n172 & n361 ;
  assign n363 = G17 & ~n362 ;
  assign n364 = ~G17 & n362 ;
  assign n365 = n363 | n364 ;
  assign n366 = n191 & n361 ;
  assign n367 = G18 & ~n366 ;
  assign n368 = ~G18 & n366 ;
  assign n369 = n367 | n368 ;
  assign n370 = n115 & n361 ;
  assign n371 = G19 & ~n370 ;
  assign n372 = ~G19 & n370 ;
  assign n373 = n371 | n372 ;
  assign n374 = n152 & n361 ;
  assign n375 = G20 & ~n374 ;
  assign n376 = ~G20 & n374 ;
  assign n377 = n375 | n376 ;
  assign n378 = n252 & n272 ;
  assign n379 = n359 & n378 ;
  assign n380 = n172 & n379 ;
  assign n381 = G21 & ~n380 ;
  assign n382 = ~G21 & n380 ;
  assign n383 = n381 | n382 ;
  assign n384 = n191 & n379 ;
  assign n385 = G22 & ~n384 ;
  assign n386 = ~G22 & n384 ;
  assign n387 = n385 | n386 ;
  assign n388 = n115 & n379 ;
  assign n389 = G23 & ~n388 ;
  assign n390 = ~G23 & n388 ;
  assign n391 = n389 | n390 ;
  assign n392 = n152 & n379 ;
  assign n393 = G24 & ~n392 ;
  assign n394 = ~G24 & n392 ;
  assign n395 = n393 | n394 ;
  assign n396 = n230 & n360 ;
  assign n397 = n172 & n396 ;
  assign n398 = G25 & ~n397 ;
  assign n399 = ~G25 & n397 ;
  assign n400 = n398 | n399 ;
  assign n401 = n191 & n396 ;
  assign n402 = G26 & ~n401 ;
  assign n403 = ~G26 & n401 ;
  assign n404 = n402 | n403 ;
  assign n405 = n115 & n396 ;
  assign n406 = G27 & ~n405 ;
  assign n407 = ~G27 & n405 ;
  assign n408 = n406 | n407 ;
  assign n409 = n152 & n396 ;
  assign n410 = G28 & ~n409 ;
  assign n411 = ~G28 & n409 ;
  assign n412 = n410 | n411 ;
  assign n413 = n250 & n272 ;
  assign n414 = n359 & n413 ;
  assign n415 = n172 & n414 ;
  assign n416 = G29 | n415 ;
  assign n417 = G29 & n415 ;
  assign n418 = n416 & ~n417 ;
  assign n419 = n191 & n414 ;
  assign n420 = G30 & ~n419 ;
  assign n421 = ~G30 & n419 ;
  assign n422 = n420 | n421 ;
  assign n423 = n115 & n414 ;
  assign n424 = G31 & ~n423 ;
  assign n425 = ~G31 & n423 ;
  assign n426 = n424 | n425 ;
  assign n427 = n152 & n414 ;
  assign n428 = G32 | n427 ;
  assign n429 = G32 & n427 ;
  assign n430 = n428 & ~n429 ;
  assign G1324 = ~n285 ;
  assign G1325 = ~n289 ;
  assign G1326 = ~n293 ;
  assign G1327 = ~n297 ;
  assign G1328 = ~n303 ;
  assign G1329 = ~n307 ;
  assign G1330 = ~n311 ;
  assign G1331 = ~n315 ;
  assign G1332 = ~n322 ;
  assign G1333 = ~n326 ;
  assign G1334 = ~n330 ;
  assign G1335 = ~n334 ;
  assign G1336 = ~n340 ;
  assign G1337 = ~n344 ;
  assign G1338 = ~n348 ;
  assign G1339 = ~n352 ;
  assign G1340 = ~n365 ;
  assign G1341 = ~n369 ;
  assign G1342 = ~n373 ;
  assign G1343 = ~n377 ;
  assign G1344 = ~n383 ;
  assign G1345 = ~n387 ;
  assign G1346 = ~n391 ;
  assign G1347 = ~n395 ;
  assign G1348 = ~n400 ;
  assign G1349 = ~n404 ;
  assign G1350 = ~n408 ;
  assign G1351 = ~n412 ;
  assign G1352 = ~n418 ;
  assign G1353 = ~n422 ;
  assign G1354 = ~n426 ;
  assign G1355 = ~n430 ;
endmodule
