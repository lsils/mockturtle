module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 ;
  wire n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 ;
  assign n179 = x152 & x155 ;
  assign n180 = x65 & x66 ;
  assign n181 = x0 & x133 ;
  assign n182 = x62 & ~x164 ;
  assign n183 = x10 & ~x163 ;
  assign n184 = x135 & x153 ;
  assign n185 = x10 & x11 ;
  assign n186 = x64 & n185 ;
  assign n187 = ( x32 & x162 ) | ( x32 & n185 ) | ( x162 & n185 ) ;
  assign n188 = ( x33 & ~x162 ) | ( x33 & n185 ) | ( ~x162 & n185 ) ;
  assign n189 = n187 & n188 ;
  assign n190 = ( x34 & x162 ) | ( x34 & n185 ) | ( x162 & n185 ) ;
  assign n191 = ( x12 & ~x162 ) | ( x12 & n185 ) | ( ~x162 & n185 ) ;
  assign n192 = n190 & n191 ;
  assign n193 = x31 & n185 ;
  assign n194 = ( ~x7 & x162 ) | ( ~x7 & n185 ) | ( x162 & n185 ) ;
  assign n195 = ( x8 & x162 ) | ( x8 & ~n185 ) | ( x162 & ~n185 ) ;
  assign n196 = n194 & ~n195 ;
  assign n197 = x65 & ~n196 ;
  assign n198 = ( ~x9 & x162 ) | ( ~x9 & n185 ) | ( x162 & n185 ) ;
  assign n199 = ( x29 & x162 ) | ( x29 & ~n185 ) | ( x162 & ~n185 ) ;
  assign n200 = n198 & ~n199 ;
  assign n201 = x65 & ~n200 ;
  assign n202 = ( ~x27 & x162 ) | ( ~x27 & n185 ) | ( x162 & n185 ) ;
  assign n203 = ( x6 & x162 ) | ( x6 & ~n185 ) | ( x162 & ~n185 ) ;
  assign n204 = n202 & ~n203 ;
  assign n205 = x65 & ~n204 ;
  assign n206 = ( ~x30 & x162 ) | ( ~x30 & n185 ) | ( x162 & n185 ) ;
  assign n207 = ( x28 & x162 ) | ( x28 & ~n185 ) | ( x162 & ~n185 ) ;
  assign n208 = n206 & ~n207 ;
  assign n209 = x65 & ~n208 ;
  assign n213 = ( x120 & ~x146 ) | ( x120 & x166 ) | ( ~x146 & x166 ) ;
  assign n214 = ( x120 & x146 ) | ( x120 & ~x165 ) | ( x146 & ~x165 ) ;
  assign n215 = n213 & ~n214 ;
  assign n216 = ( x120 & ~x146 ) | ( x120 & x168 ) | ( ~x146 & x168 ) ;
  assign n217 = ( x120 & x146 ) | ( x120 & ~x167 ) | ( x146 & ~x167 ) ;
  assign n218 = ~n216 & n217 ;
  assign n219 = n215 | n218 ;
  assign n227 = ( x125 & ~x148 ) | ( x125 & x166 ) | ( ~x148 & x166 ) ;
  assign n228 = ( x125 & x148 ) | ( x125 & ~x165 ) | ( x148 & ~x165 ) ;
  assign n229 = n227 & ~n228 ;
  assign n230 = ( x125 & ~x148 ) | ( x125 & x168 ) | ( ~x148 & x168 ) ;
  assign n231 = ( x125 & x148 ) | ( x125 & ~x167 ) | ( x148 & ~x167 ) ;
  assign n232 = ~n230 & n231 ;
  assign n233 = n229 | n232 ;
  assign n220 = ( x127 & ~x149 ) | ( x127 & x166 ) | ( ~x149 & x166 ) ;
  assign n221 = ( x127 & x149 ) | ( x127 & ~x165 ) | ( x149 & ~x165 ) ;
  assign n222 = n220 & ~n221 ;
  assign n223 = ( x127 & ~x149 ) | ( x127 & x168 ) | ( ~x149 & x168 ) ;
  assign n224 = ( x127 & x149 ) | ( x127 & ~x167 ) | ( x149 & ~x167 ) ;
  assign n225 = ~n223 & n224 ;
  assign n226 = n222 | n225 ;
  assign n234 = x147 & ~x168 ;
  assign n235 = x147 | x165 ;
  assign n236 = ( ~x147 & n234 ) | ( ~x147 & n235 ) | ( n234 & n235 ) ;
  assign n237 = n226 & n236 ;
  assign n238 = ( ~n219 & n233 ) | ( ~n219 & n237 ) | ( n233 & n237 ) ;
  assign n239 = n219 & n238 ;
  assign n210 = ~x99 & x129 ;
  assign n211 = x100 & ~x129 ;
  assign n212 = ( x129 & ~n210 ) | ( x129 & n211 ) | ( ~n210 & n211 ) ;
  assign n240 = ( x101 & ~x118 ) | ( x101 & x145 ) | ( ~x118 & x145 ) ;
  assign n241 = ( x97 & x118 ) | ( x97 & x145 ) | ( x118 & x145 ) ;
  assign n242 = n240 | n241 ;
  assign n243 = ( x99 & ~x118 ) | ( x99 & x145 ) | ( ~x118 & x145 ) ;
  assign n244 = ( x100 & x118 ) | ( x100 & x145 ) | ( x118 & x145 ) ;
  assign n245 = n243 & n244 ;
  assign n246 = n242 & ~n245 ;
  assign n254 = ~x99 & x114 ;
  assign n255 = x100 & ~x114 ;
  assign n256 = ( x114 & ~n254 ) | ( x114 & n255 ) | ( ~n254 & n255 ) ;
  assign n247 = ( x101 & ~x116 ) | ( x101 & x144 ) | ( ~x116 & x144 ) ;
  assign n248 = ( x97 & x116 ) | ( x97 & x144 ) | ( x116 & x144 ) ;
  assign n249 = n247 | n248 ;
  assign n250 = ( x99 & ~x116 ) | ( x99 & x144 ) | ( ~x116 & x144 ) ;
  assign n251 = ( x100 & x116 ) | ( x100 & x144 ) | ( x116 & x144 ) ;
  assign n252 = n250 & n251 ;
  assign n253 = n249 & ~n252 ;
  assign n257 = ~x97 & x112 ;
  assign n258 = x101 & ~x112 ;
  assign n259 = ( x112 & ~n257 ) | ( x112 & n258 ) | ( ~n257 & n258 ) ;
  assign n260 = n253 | n259 ;
  assign n261 = ( n246 & n256 ) | ( n246 & ~n260 ) | ( n256 & ~n260 ) ;
  assign n262 = ~n246 & n261 ;
  assign n263 = n212 & n262 ;
  assign n264 = n239 & n263 ;
  assign n272 = ( x102 & ~x136 ) | ( x102 & x166 ) | ( ~x136 & x166 ) ;
  assign n273 = ( x102 & x136 ) | ( x102 & ~x165 ) | ( x136 & ~x165 ) ;
  assign n274 = n272 & ~n273 ;
  assign n275 = ( x102 & ~x136 ) | ( x102 & x168 ) | ( ~x136 & x168 ) ;
  assign n276 = ( x102 & x136 ) | ( x102 & ~x167 ) | ( x136 & ~x167 ) ;
  assign n277 = ~n275 & n276 ;
  assign n278 = n274 | n277 ;
  assign n286 = ( x108 & ~x134 ) | ( x108 & x166 ) | ( ~x134 & x166 ) ;
  assign n287 = ( x108 & x134 ) | ( x108 & ~x165 ) | ( x134 & ~x165 ) ;
  assign n288 = n286 & ~n287 ;
  assign n289 = ( x108 & ~x134 ) | ( x108 & x168 ) | ( ~x134 & x168 ) ;
  assign n290 = ( x108 & x134 ) | ( x108 & ~x167 ) | ( x134 & ~x167 ) ;
  assign n291 = ~n289 & n290 ;
  assign n292 = n288 | n291 ;
  assign n279 = ( x104 & ~x137 ) | ( x104 & x166 ) | ( ~x137 & x166 ) ;
  assign n280 = ( x104 & x137 ) | ( x104 & ~x165 ) | ( x137 & ~x165 ) ;
  assign n281 = n279 & ~n280 ;
  assign n282 = ( x104 & ~x137 ) | ( x104 & x168 ) | ( ~x137 & x168 ) ;
  assign n283 = ( x104 & x137 ) | ( x104 & ~x167 ) | ( x137 & ~x167 ) ;
  assign n284 = ~n282 & n283 ;
  assign n285 = n281 | n284 ;
  assign n293 = ( x106 & ~x138 ) | ( x106 & x166 ) | ( ~x138 & x166 ) ;
  assign n294 = ( x106 & x138 ) | ( x106 & ~x165 ) | ( x138 & ~x165 ) ;
  assign n295 = n293 & ~n294 ;
  assign n296 = ( x106 & ~x138 ) | ( x106 & x168 ) | ( ~x138 & x168 ) ;
  assign n297 = ( x106 & x138 ) | ( x106 & ~x167 ) | ( x138 & ~x167 ) ;
  assign n298 = ~n296 & n297 ;
  assign n299 = n295 | n298 ;
  assign n300 = n285 & n299 ;
  assign n301 = ( ~n278 & n292 ) | ( ~n278 & n300 ) | ( n292 & n300 ) ;
  assign n302 = n278 & n301 ;
  assign n265 = ( ~x87 & x101 ) | ( ~x87 & x141 ) | ( x101 & x141 ) ;
  assign n266 = ( x87 & x97 ) | ( x87 & x141 ) | ( x97 & x141 ) ;
  assign n267 = n265 | n266 ;
  assign n268 = ( ~x87 & x99 ) | ( ~x87 & x141 ) | ( x99 & x141 ) ;
  assign n269 = ( x87 & x100 ) | ( x87 & x141 ) | ( x100 & x141 ) ;
  assign n270 = n268 & n269 ;
  assign n271 = n267 & ~n270 ;
  assign n303 = ( x89 & ~x142 ) | ( x89 & x166 ) | ( ~x142 & x166 ) ;
  assign n304 = ( x89 & x142 ) | ( x89 & ~x165 ) | ( x142 & ~x165 ) ;
  assign n305 = n303 & ~n304 ;
  assign n306 = ( x89 & ~x142 ) | ( x89 & x168 ) | ( ~x142 & x168 ) ;
  assign n307 = ( x89 & x142 ) | ( x89 & ~x167 ) | ( x142 & ~x167 ) ;
  assign n308 = ~n306 & n307 ;
  assign n309 = n305 | n308 ;
  assign n317 = ( x95 & ~x140 ) | ( x95 & x166 ) | ( ~x140 & x166 ) ;
  assign n318 = ( x95 & x140 ) | ( x95 & ~x165 ) | ( x140 & ~x165 ) ;
  assign n319 = n317 & ~n318 ;
  assign n320 = ( x95 & ~x140 ) | ( x95 & x168 ) | ( ~x140 & x168 ) ;
  assign n321 = ( x95 & x140 ) | ( x95 & ~x167 ) | ( x140 & ~x167 ) ;
  assign n322 = ~n320 & n321 ;
  assign n323 = n319 | n322 ;
  assign n310 = ( x91 & ~x143 ) | ( x91 & x166 ) | ( ~x143 & x166 ) ;
  assign n311 = ( x91 & x143 ) | ( x91 & ~x165 ) | ( x143 & ~x165 ) ;
  assign n312 = n310 & ~n311 ;
  assign n313 = ( x91 & ~x143 ) | ( x91 & x168 ) | ( ~x143 & x168 ) ;
  assign n314 = ( x91 & x143 ) | ( x91 & ~x167 ) | ( x143 & ~x167 ) ;
  assign n315 = ~n313 & n314 ;
  assign n316 = n312 | n315 ;
  assign n324 = ( x93 & ~x139 ) | ( x93 & x166 ) | ( ~x139 & x166 ) ;
  assign n325 = ( x93 & x139 ) | ( x93 & ~x165 ) | ( x139 & ~x165 ) ;
  assign n326 = n324 & ~n325 ;
  assign n327 = ( x93 & ~x139 ) | ( x93 & x168 ) | ( ~x139 & x168 ) ;
  assign n328 = ( x93 & x139 ) | ( x93 & ~x167 ) | ( x139 & ~x167 ) ;
  assign n329 = ~n327 & n328 ;
  assign n330 = n326 | n329 ;
  assign n331 = n316 & n330 ;
  assign n332 = ( ~n309 & n323 ) | ( ~n309 & n331 ) | ( n323 & n331 ) ;
  assign n333 = n309 & n332 ;
  assign n334 = ~n271 & n333 ;
  assign n335 = n302 & n334 ;
  assign n336 = ~x96 & x123 ;
  assign n337 = x95 & ~x123 ;
  assign n338 = ( x123 & ~n336 ) | ( x123 & n337 ) | ( ~n336 & n337 ) ;
  assign n339 = x140 | n338 ;
  assign n340 = ~x140 & n338 ;
  assign n341 = ( ~n338 & n339 ) | ( ~n338 & n340 ) | ( n339 & n340 ) ;
  assign n342 = ~x103 & x123 ;
  assign n343 = x102 & ~x123 ;
  assign n344 = ( x123 & ~n342 ) | ( x123 & n343 ) | ( ~n342 & n343 ) ;
  assign n345 = x136 | n344 ;
  assign n346 = ~x136 & n344 ;
  assign n347 = ( ~n344 & n345 ) | ( ~n344 & n346 ) | ( n345 & n346 ) ;
  assign n354 = ~x109 & x123 ;
  assign n355 = x108 & ~x123 ;
  assign n356 = ( x123 & ~n354 ) | ( x123 & n355 ) | ( ~n354 & n355 ) ;
  assign n357 = x134 | n356 ;
  assign n358 = ~x134 & n356 ;
  assign n359 = ( ~n356 & n357 ) | ( ~n356 & n358 ) | ( n357 & n358 ) ;
  assign n348 = ~x105 & x123 ;
  assign n349 = x104 & ~x123 ;
  assign n350 = ( x123 & ~n348 ) | ( x123 & n349 ) | ( ~n348 & n349 ) ;
  assign n351 = x137 | n350 ;
  assign n352 = ~x137 & n350 ;
  assign n353 = ( ~n350 & n351 ) | ( ~n350 & n352 ) | ( n351 & n352 ) ;
  assign n360 = ~x107 & x123 ;
  assign n361 = x106 & ~x123 ;
  assign n362 = ( x123 & ~n360 ) | ( x123 & n361 ) | ( ~n360 & n361 ) ;
  assign n363 = x138 | n362 ;
  assign n364 = ~x138 & n362 ;
  assign n365 = ( ~n362 & n363 ) | ( ~n362 & n364 ) | ( n363 & n364 ) ;
  assign n366 = n353 & n365 ;
  assign n367 = ( ~n347 & n359 ) | ( ~n347 & n366 ) | ( n359 & n366 ) ;
  assign n368 = n347 & n367 ;
  assign n369 = n341 & n368 ;
  assign n370 = ~x88 & x123 ;
  assign n371 = x87 & ~x123 ;
  assign n372 = ( x123 & ~n370 ) | ( x123 & n371 ) | ( ~n370 & n371 ) ;
  assign n373 = x141 | n372 ;
  assign n374 = ~x141 & n372 ;
  assign n375 = ( ~n372 & n373 ) | ( ~n372 & n374 ) | ( n373 & n374 ) ;
  assign n382 = ~x94 & x123 ;
  assign n383 = x93 & ~x123 ;
  assign n384 = ( x123 & ~n382 ) | ( x123 & n383 ) | ( ~n382 & n383 ) ;
  assign n385 = x139 | n384 ;
  assign n386 = ~x139 & n384 ;
  assign n387 = ( ~n384 & n385 ) | ( ~n384 & n386 ) | ( n385 & n386 ) ;
  assign n376 = ~x90 & x123 ;
  assign n377 = x89 & ~x123 ;
  assign n378 = ( x123 & ~n376 ) | ( x123 & n377 ) | ( ~n376 & n377 ) ;
  assign n379 = x142 | n378 ;
  assign n380 = ~x142 & n378 ;
  assign n381 = ( ~n378 & n379 ) | ( ~n378 & n380 ) | ( n379 & n380 ) ;
  assign n388 = ~x92 & x123 ;
  assign n389 = x91 & ~x123 ;
  assign n390 = ( x123 & ~n388 ) | ( x123 & n389 ) | ( ~n388 & n389 ) ;
  assign n391 = x143 | n390 ;
  assign n392 = ~x143 & n390 ;
  assign n393 = ( ~n390 & n391 ) | ( ~n390 & n392 ) | ( n391 & n392 ) ;
  assign n394 = n381 & n393 ;
  assign n395 = ( ~n375 & n387 ) | ( ~n375 & n394 ) | ( n387 & n394 ) ;
  assign n396 = n375 & n395 ;
  assign n397 = n369 & n396 ;
  assign n398 = x122 & ~x128 ;
  assign n399 = ~x122 & x127 ;
  assign n400 = ( x122 & ~n398 ) | ( x122 & n399 ) | ( ~n398 & n399 ) ;
  assign n401 = x149 | n400 ;
  assign n402 = ~x149 & n400 ;
  assign n403 = ( ~n400 & n401 ) | ( ~n400 & n402 ) | ( n401 & n402 ) ;
  assign n410 = x122 & ~x126 ;
  assign n411 = ~x122 & x125 ;
  assign n412 = ( x122 & ~n410 ) | ( x122 & n411 ) | ( ~n410 & n411 ) ;
  assign n413 = x148 | n412 ;
  assign n414 = ~x148 & n412 ;
  assign n415 = ( ~n412 & n413 ) | ( ~n412 & n414 ) | ( n413 & n414 ) ;
  assign n404 = ~x121 & x122 ;
  assign n405 = x120 & ~x122 ;
  assign n406 = ( x122 & ~n404 ) | ( x122 & n405 ) | ( ~n404 & n405 ) ;
  assign n407 = x146 | n406 ;
  assign n408 = ~x146 & n406 ;
  assign n409 = ( ~n406 & n407 ) | ( ~n406 & n408 ) | ( n407 & n408 ) ;
  assign n416 = x122 & ~x124 ;
  assign n417 = ~x147 & n416 ;
  assign n418 = x147 | n416 ;
  assign n419 = ( ~n416 & n417 ) | ( ~n416 & n418 ) | ( n417 & n418 ) ;
  assign n420 = x122 & ~x130 ;
  assign n421 = ~x122 & x129 ;
  assign n422 = ( x122 & ~n420 ) | ( x122 & n421 ) | ( ~n420 & n421 ) ;
  assign n423 = n419 | n422 ;
  assign n424 = n409 & ~n423 ;
  assign n425 = ( ~n403 & n415 ) | ( ~n403 & n424 ) | ( n415 & n424 ) ;
  assign n426 = n403 & n425 ;
  assign n427 = ~x117 & x122 ;
  assign n428 = x116 & ~x122 ;
  assign n429 = ( x122 & ~n427 ) | ( x122 & n428 ) | ( ~n427 & n428 ) ;
  assign n430 = x144 | n429 ;
  assign n431 = ~x144 & n429 ;
  assign n432 = ( ~n429 & n430 ) | ( ~n429 & n431 ) | ( n430 & n431 ) ;
  assign n439 = ~x113 & x122 ;
  assign n440 = x112 & ~x122 ;
  assign n441 = ( x122 & ~n439 ) | ( x122 & n440 ) | ( ~n439 & n440 ) ;
  assign n433 = ~x119 & x122 ;
  assign n434 = x118 & ~x122 ;
  assign n435 = ( x122 & ~n433 ) | ( x122 & n434 ) | ( ~n433 & n434 ) ;
  assign n436 = x145 | n435 ;
  assign n437 = ~x145 & n435 ;
  assign n438 = ( ~n435 & n436 ) | ( ~n435 & n437 ) | ( n436 & n437 ) ;
  assign n442 = ~x115 & x122 ;
  assign n443 = x114 & ~x122 ;
  assign n444 = ( x122 & ~n442 ) | ( x122 & n443 ) | ( ~n442 & n443 ) ;
  assign n445 = n438 & ~n444 ;
  assign n446 = ( n432 & n441 ) | ( n432 & ~n445 ) | ( n441 & ~n445 ) ;
  assign n447 = n432 & ~n446 ;
  assign n448 = n426 & n447 ;
  assign n449 = n403 & ~n422 ;
  assign n450 = n415 & n449 ;
  assign n451 = ( n409 & n419 ) | ( n409 & ~n450 ) | ( n419 & ~n450 ) ;
  assign n452 = n409 & ~n451 ;
  assign n453 = n447 & n452 ;
  assign n454 = n347 & n359 ;
  assign n455 = ( ~n341 & n353 ) | ( ~n341 & n454 ) | ( n353 & n454 ) ;
  assign n456 = n341 & n455 ;
  assign n457 = n365 & n456 ;
  assign n458 = n396 & n457 ;
  assign n459 = x125 & ~x127 ;
  assign n460 = x125 | x127 ;
  assign n461 = ( ~x125 & n459 ) | ( ~x125 & n460 ) | ( n459 & n460 ) ;
  assign n462 = ( x120 & x129 ) | ( x120 & ~n461 ) | ( x129 & ~n461 ) ;
  assign n463 = ( ~x120 & n461 ) | ( ~x120 & n462 ) | ( n461 & n462 ) ;
  assign n464 = ( ~x129 & n462 ) | ( ~x129 & n463 ) | ( n462 & n463 ) ;
  assign n465 = x131 | n464 ;
  assign n466 = x131 & n464 ;
  assign n467 = n465 & ~n466 ;
  assign n468 = ( x112 & x114 ) | ( x112 & x116 ) | ( x114 & x116 ) ;
  assign n469 = ( x112 & x114 ) | ( x112 & ~n468 ) | ( x114 & ~n468 ) ;
  assign n470 = ( x116 & ~n468 ) | ( x116 & n469 ) | ( ~n468 & n469 ) ;
  assign n471 = ~x118 & n470 ;
  assign n472 = x118 & ~n470 ;
  assign n473 = n471 | n472 ;
  assign n474 = n467 & n473 ;
  assign n475 = ~n467 & n473 ;
  assign n476 = ( n467 & ~n474 ) | ( n467 & n475 ) | ( ~n474 & n475 ) ;
  assign n477 = x108 & ~x110 ;
  assign n478 = x108 | x110 ;
  assign n479 = ( ~x108 & n477 ) | ( ~x108 & n478 ) | ( n477 & n478 ) ;
  assign n480 = x104 & ~x106 ;
  assign n481 = x104 | x106 ;
  assign n482 = ( ~x104 & n480 ) | ( ~x104 & n481 ) | ( n480 & n481 ) ;
  assign n483 = ( ~x95 & n479 ) | ( ~x95 & n482 ) | ( n479 & n482 ) ;
  assign n484 = ( n479 & n482 ) | ( n479 & ~n483 ) | ( n482 & ~n483 ) ;
  assign n485 = ( x95 & n483 ) | ( x95 & ~n484 ) | ( n483 & ~n484 ) ;
  assign n486 = ~x102 & n485 ;
  assign n487 = x102 & ~n485 ;
  assign n488 = n486 | n487 ;
  assign n489 = ( x87 & x89 ) | ( x87 & x91 ) | ( x89 & x91 ) ;
  assign n490 = ( x87 & x89 ) | ( x87 & ~n489 ) | ( x89 & ~n489 ) ;
  assign n491 = ( x91 & ~n489 ) | ( x91 & n490 ) | ( ~n489 & n490 ) ;
  assign n492 = ~x93 & n491 ;
  assign n493 = x93 & ~n491 ;
  assign n494 = n492 | n493 ;
  assign n495 = ~n488 & n494 ;
  assign n496 = n488 & n494 ;
  assign n497 = ( n488 & n495 ) | ( n488 & ~n496 ) | ( n495 & ~n496 ) ;
  assign n515 = x143 & n390 ;
  assign n519 = ( ~n375 & n381 ) | ( ~n375 & n515 ) | ( n381 & n515 ) ;
  assign n516 = x139 & n384 ;
  assign n517 = n375 & n516 ;
  assign n518 = n393 & n517 ;
  assign n520 = n381 & n518 ;
  assign n521 = ( n375 & n519 ) | ( n375 & n520 ) | ( n519 & n520 ) ;
  assign n514 = x142 & n378 ;
  assign n522 = ( x141 & n372 ) | ( x141 & n514 ) | ( n372 & n514 ) ;
  assign n523 = n521 | n522 ;
  assign n498 = x138 & n353 ;
  assign n499 = ( ~n341 & n362 ) | ( ~n341 & n498 ) | ( n362 & n498 ) ;
  assign n500 = n341 & n499 ;
  assign n501 = x134 & n356 ;
  assign n502 = n353 & n501 ;
  assign n503 = ( ~n341 & n365 ) | ( ~n341 & n502 ) | ( n365 & n502 ) ;
  assign n504 = n341 & n503 ;
  assign n505 = x137 & n350 ;
  assign n506 = x136 & n344 ;
  assign n507 = ( x140 & n338 ) | ( x140 & n506 ) | ( n338 & n506 ) ;
  assign n508 = ( n341 & n347 ) | ( n341 & n507 ) | ( n347 & n507 ) ;
  assign n509 = n505 & ~n508 ;
  assign n510 = ( n505 & n507 ) | ( n505 & ~n509 ) | ( n507 & ~n509 ) ;
  assign n511 = ( ~n500 & n504 ) | ( ~n500 & n510 ) | ( n504 & n510 ) ;
  assign n512 = n347 | n510 ;
  assign n513 = ( n500 & n511 ) | ( n500 & n512 ) | ( n511 & n512 ) ;
  assign n524 = n513 | n523 ;
  assign n525 = ( n396 & n523 ) | ( n396 & n524 ) | ( n523 & n524 ) ;
  assign n541 = x145 & n435 ;
  assign n542 = n432 & ~n441 ;
  assign n543 = n541 & n542 ;
  assign n544 = x144 & n429 ;
  assign n545 = n444 | n544 ;
  assign n546 = ( n441 & ~n543 ) | ( n441 & n545 ) | ( ~n543 & n545 ) ;
  assign n547 = n543 | n546 ;
  assign n526 = x149 & n415 ;
  assign n527 = ( n400 & ~n409 ) | ( n400 & n526 ) | ( ~n409 & n526 ) ;
  assign n528 = n409 & n527 ;
  assign n529 = n409 & n422 ;
  assign n530 = ( ~n403 & n415 ) | ( ~n403 & n529 ) | ( n415 & n529 ) ;
  assign n531 = n403 & n530 ;
  assign n532 = x148 & n412 ;
  assign n533 = x147 & ~n416 ;
  assign n534 = ( x146 & n406 ) | ( x146 & n533 ) | ( n406 & n533 ) ;
  assign n535 = ( n409 & ~n419 ) | ( n409 & n534 ) | ( ~n419 & n534 ) ;
  assign n536 = n532 & ~n535 ;
  assign n537 = ( n532 & n534 ) | ( n532 & ~n536 ) | ( n534 & ~n536 ) ;
  assign n538 = ( ~n528 & n531 ) | ( ~n528 & n537 ) | ( n531 & n537 ) ;
  assign n539 = n419 & ~n537 ;
  assign n540 = ( n528 & n538 ) | ( n528 & ~n539 ) | ( n538 & ~n539 ) ;
  assign n548 = n540 | n547 ;
  assign n549 = ( n447 & n547 ) | ( n447 & n548 ) | ( n547 & n548 ) ;
  assign n553 = ( ~x175 & x176 ) | ( ~x175 & n212 ) | ( x176 & n212 ) ;
  assign n550 = x20 | n422 ;
  assign n551 = ~x20 & n422 ;
  assign n552 = ( ~n422 & n550 ) | ( ~n422 & n551 ) | ( n550 & n551 ) ;
  assign n554 = ( x175 & x176 ) | ( x175 & n552 ) | ( x176 & n552 ) ;
  assign n555 = n553 | n554 ;
  assign n556 = ( ~x59 & x175 ) | ( ~x59 & n555 ) | ( x175 & n555 ) ;
  assign n557 = x176 & n556 ;
  assign n558 = ( ~x176 & n555 ) | ( ~x176 & n557 ) | ( n555 & n557 ) ;
  assign n562 = ( ~x175 & x176 ) | ( ~x175 & n226 ) | ( x176 & n226 ) ;
  assign n559 = ( x20 & n403 ) | ( x20 & ~n551 ) | ( n403 & ~n551 ) ;
  assign n560 = ( x20 & ~n403 ) | ( x20 & n551 ) | ( ~n403 & n551 ) ;
  assign n561 = ( ~x20 & n559 ) | ( ~x20 & n560 ) | ( n559 & n560 ) ;
  assign n563 = ( x175 & x176 ) | ( x175 & ~n561 ) | ( x176 & ~n561 ) ;
  assign n564 = n562 | n563 ;
  assign n565 = ( ~x57 & x175 ) | ( ~x57 & n564 ) | ( x175 & n564 ) ;
  assign n566 = x176 & n565 ;
  assign n567 = ( ~x176 & n564 ) | ( ~x176 & n566 ) | ( n564 & n566 ) ;
  assign n571 = ( ~x175 & x176 ) | ( ~x175 & n292 ) | ( x176 & n292 ) ;
  assign n568 = x1 | n359 ;
  assign n569 = ~x1 & n359 ;
  assign n570 = ( ~n359 & n568 ) | ( ~n359 & n569 ) | ( n568 & n569 ) ;
  assign n572 = ( x175 & x176 ) | ( x175 & ~n570 ) | ( x176 & ~n570 ) ;
  assign n573 = n571 | n572 ;
  assign n574 = ( ~x47 & x175 ) | ( ~x47 & n573 ) | ( x175 & n573 ) ;
  assign n575 = x176 & n574 ;
  assign n576 = ( ~x176 & n573 ) | ( ~x176 & n575 ) | ( n573 & n575 ) ;
  assign n577 = ( x144 & n429 ) | ( x144 & n541 ) | ( n429 & n541 ) ;
  assign n578 = n444 | n577 ;
  assign n583 = x20 | n540 ;
  assign n584 = ( n426 & n540 ) | ( n426 & n583 ) | ( n540 & n583 ) ;
  assign n585 = n578 & ~n584 ;
  assign n579 = x145 & ~n435 ;
  assign n580 = n432 & ~n444 ;
  assign n581 = ( n435 & n579 ) | ( n435 & n580 ) | ( n579 & n580 ) ;
  assign n582 = n545 | n581 ;
  assign n586 = n582 & n584 ;
  assign n587 = ( ~n441 & n585 ) | ( ~n441 & n586 ) | ( n585 & n586 ) ;
  assign n588 = ( n441 & ~n586 ) | ( n441 & n587 ) | ( ~n586 & n587 ) ;
  assign n589 = ( ~n585 & n587 ) | ( ~n585 & n588 ) | ( n587 & n588 ) ;
  assign n590 = ( x171 & ~x172 ) | ( x171 & n558 ) | ( ~x172 & n558 ) ;
  assign n591 = ( x171 & x172 ) | ( x171 & n576 ) | ( x172 & n576 ) ;
  assign n592 = n590 | n591 ;
  assign n593 = ( x21 & x171 ) | ( x21 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n594 = ( x2 & x171 ) | ( x2 & x172 ) | ( x171 & x172 ) ;
  assign n595 = n593 & n594 ;
  assign n596 = n592 & ~n595 ;
  assign n611 = ( ~x175 & x176 ) | ( ~x175 & n219 ) | ( x176 & n219 ) ;
  assign n597 = n403 & n422 ;
  assign n598 = n415 & n597 ;
  assign n599 = x20 & n415 ;
  assign n600 = ( n403 & n422 ) | ( n403 & ~n599 ) | ( n422 & ~n599 ) ;
  assign n601 = n403 & ~n600 ;
  assign n602 = n400 & n526 ;
  assign n603 = n532 | n602 ;
  assign n604 = ( x147 & ~n416 ) | ( x147 & n603 ) | ( ~n416 & n603 ) ;
  assign n605 = ( ~n598 & n601 ) | ( ~n598 & n604 ) | ( n601 & n604 ) ;
  assign n606 = n419 & ~n604 ;
  assign n607 = ( n598 & n605 ) | ( n598 & ~n606 ) | ( n605 & ~n606 ) ;
  assign n608 = n409 & ~n607 ;
  assign n609 = n409 & n607 ;
  assign n610 = ( n607 & n608 ) | ( n607 & ~n609 ) | ( n608 & ~n609 ) ;
  assign n612 = ( x175 & x176 ) | ( x175 & ~n610 ) | ( x176 & ~n610 ) ;
  assign n613 = n611 | n612 ;
  assign n614 = ( ~x18 & x175 ) | ( ~x18 & n613 ) | ( x175 & n613 ) ;
  assign n615 = x176 & n614 ;
  assign n616 = ( ~x176 & n613 ) | ( ~x176 & n615 ) | ( n613 & n615 ) ;
  assign n622 = ( ~x175 & x176 ) | ( ~x175 & n236 ) | ( x176 & n236 ) ;
  assign n617 = n598 | n601 ;
  assign n618 = n603 | n617 ;
  assign n619 = n419 & n618 ;
  assign n620 = n419 | n618 ;
  assign n621 = ~n619 & n620 ;
  assign n623 = ( x175 & x176 ) | ( x175 & n621 ) | ( x176 & n621 ) ;
  assign n624 = n622 | n623 ;
  assign n625 = ( ~x58 & x175 ) | ( ~x58 & n624 ) | ( x175 & n624 ) ;
  assign n626 = x176 & n625 ;
  assign n627 = ( ~x176 & n624 ) | ( ~x176 & n626 ) | ( n624 & n626 ) ;
  assign n632 = ( ~x175 & x176 ) | ( ~x175 & n233 ) | ( x176 & n233 ) ;
  assign n628 = ( x149 & n400 ) | ( x149 & n550 ) | ( n400 & n550 ) ;
  assign n629 = ~n415 & n628 ;
  assign n630 = n415 & n628 ;
  assign n631 = ( n415 & n629 ) | ( n415 & ~n630 ) | ( n629 & ~n630 ) ;
  assign n633 = ( x175 & x176 ) | ( x175 & ~n631 ) | ( x176 & ~n631 ) ;
  assign n634 = n632 | n633 ;
  assign n635 = ( ~x49 & x175 ) | ( ~x49 & n634 ) | ( x175 & n634 ) ;
  assign n636 = x176 & n635 ;
  assign n637 = ( ~x176 & n634 ) | ( ~x176 & n636 ) | ( n634 & n636 ) ;
  assign n638 = ( ~x173 & x174 ) | ( ~x173 & n558 ) | ( x174 & n558 ) ;
  assign n639 = ( x173 & x174 ) | ( x173 & n576 ) | ( x174 & n576 ) ;
  assign n640 = n638 | n639 ;
  assign n641 = ( x21 & ~x173 ) | ( x21 & x174 ) | ( ~x173 & x174 ) ;
  assign n642 = ( x2 & x173 ) | ( x2 & x174 ) | ( x173 & x174 ) ;
  assign n643 = n641 & n642 ;
  assign n644 = n640 & ~n643 ;
  assign n658 = ( ~x175 & x176 ) | ( ~x175 & n323 ) | ( x176 & n323 ) ;
  assign n645 = n365 & n502 ;
  assign n646 = x1 & n359 ;
  assign n647 = ( ~n353 & n365 ) | ( ~n353 & n646 ) | ( n365 & n646 ) ;
  assign n648 = n353 & n647 ;
  assign n649 = n362 & n498 ;
  assign n650 = n505 | n649 ;
  assign n651 = ( x136 & n344 ) | ( x136 & n650 ) | ( n344 & n650 ) ;
  assign n652 = ( ~n645 & n648 ) | ( ~n645 & n651 ) | ( n648 & n651 ) ;
  assign n653 = n347 | n651 ;
  assign n654 = ( n645 & n652 ) | ( n645 & n653 ) | ( n652 & n653 ) ;
  assign n655 = n341 & ~n654 ;
  assign n656 = n341 & n654 ;
  assign n657 = ( n654 & n655 ) | ( n654 & ~n656 ) | ( n655 & ~n656 ) ;
  assign n659 = ( x175 & x176 ) | ( x175 & ~n657 ) | ( x176 & ~n657 ) ;
  assign n660 = n658 | n659 ;
  assign n661 = ( ~x52 & x175 ) | ( ~x52 & n660 ) | ( x175 & n660 ) ;
  assign n662 = x176 & n661 ;
  assign n663 = ( ~x176 & n660 ) | ( ~x176 & n662 ) | ( n660 & n662 ) ;
  assign n669 = ( ~x175 & x176 ) | ( ~x175 & n278 ) | ( x176 & n278 ) ;
  assign n664 = n645 | n648 ;
  assign n665 = n650 | n664 ;
  assign n666 = ~n347 & n665 ;
  assign n667 = n347 & ~n665 ;
  assign n668 = n666 | n667 ;
  assign n670 = ( x175 & x176 ) | ( x175 & ~n668 ) | ( x176 & ~n668 ) ;
  assign n671 = n669 | n670 ;
  assign n672 = ( ~x56 & x175 ) | ( ~x56 & n671 ) | ( x175 & n671 ) ;
  assign n673 = x176 & n672 ;
  assign n674 = ( ~x176 & n671 ) | ( ~x176 & n673 ) | ( n671 & n673 ) ;
  assign n682 = ( ~x175 & x176 ) | ( ~x175 & n285 ) | ( x176 & n285 ) ;
  assign n675 = ( x138 & n362 ) | ( x138 & n501 ) | ( n362 & n501 ) ;
  assign n676 = ( n359 & n365 ) | ( n359 & n675 ) | ( n365 & n675 ) ;
  assign n677 = x1 & ~n676 ;
  assign n678 = ( x1 & n675 ) | ( x1 & ~n677 ) | ( n675 & ~n677 ) ;
  assign n679 = n353 & ~n678 ;
  assign n680 = n353 & n678 ;
  assign n681 = ( n678 & n679 ) | ( n678 & ~n680 ) | ( n679 & ~n680 ) ;
  assign n683 = ( x175 & x176 ) | ( x175 & ~n681 ) | ( x176 & ~n681 ) ;
  assign n684 = n682 | n683 ;
  assign n685 = ( ~x55 & x175 ) | ( ~x55 & n684 ) | ( x175 & n684 ) ;
  assign n686 = x176 & n685 ;
  assign n687 = ( ~x176 & n684 ) | ( ~x176 & n686 ) | ( n684 & n686 ) ;
  assign n692 = ( ~x175 & x176 ) | ( ~x175 & n299 ) | ( x176 & n299 ) ;
  assign n688 = ( x1 & x134 ) | ( x1 & n356 ) | ( x134 & n356 ) ;
  assign n689 = n365 | n688 ;
  assign n690 = n365 & n688 ;
  assign n691 = n689 & ~n690 ;
  assign n693 = ( x175 & x176 ) | ( x175 & ~n691 ) | ( x176 & ~n691 ) ;
  assign n694 = n692 | n693 ;
  assign n695 = ( ~x54 & x175 ) | ( ~x54 & n694 ) | ( x175 & n694 ) ;
  assign n696 = x176 & n695 ;
  assign n697 = ( ~x176 & n694 ) | ( ~x176 & n696 ) | ( n694 & n696 ) ;
  assign n698 = ~n400 & n412 ;
  assign n699 = n400 & n412 ;
  assign n700 = ( n400 & n698 ) | ( n400 & ~n699 ) | ( n698 & ~n699 ) ;
  assign n701 = x122 & ~x132 ;
  assign n702 = x122 | x131 ;
  assign n703 = ( n422 & ~n701 ) | ( n422 & n702 ) | ( ~n701 & n702 ) ;
  assign n704 = ( n422 & n702 ) | ( n422 & ~n703 ) | ( n702 & ~n703 ) ;
  assign n705 = ( n701 & n703 ) | ( n701 & ~n704 ) | ( n703 & ~n704 ) ;
  assign n706 = ( n406 & n700 ) | ( n406 & n705 ) | ( n700 & n705 ) ;
  assign n707 = ( n700 & n705 ) | ( n700 & ~n706 ) | ( n705 & ~n706 ) ;
  assign n708 = ( n406 & ~n706 ) | ( n406 & n707 ) | ( ~n706 & n707 ) ;
  assign n709 = n416 | n708 ;
  assign n710 = n416 & n708 ;
  assign n711 = n709 & ~n710 ;
  assign n712 = ~n429 & n435 ;
  assign n713 = n429 & n435 ;
  assign n714 = ( n429 & n712 ) | ( n429 & ~n713 ) | ( n712 & ~n713 ) ;
  assign n715 = ( n441 & ~n711 ) | ( n441 & n714 ) | ( ~n711 & n714 ) ;
  assign n716 = ( n711 & ~n714 ) | ( n711 & n715 ) | ( ~n714 & n715 ) ;
  assign n717 = ( ~n441 & n715 ) | ( ~n441 & n716 ) | ( n715 & n716 ) ;
  assign n718 = n444 & n717 ;
  assign n719 = n444 | n717 ;
  assign n720 = ~n718 & n719 ;
  assign n721 = ~x111 & x123 ;
  assign n722 = x110 | x123 ;
  assign n723 = ( n372 & ~n721 ) | ( n372 & n722 ) | ( ~n721 & n722 ) ;
  assign n724 = ( n372 & n722 ) | ( n372 & ~n723 ) | ( n722 & ~n723 ) ;
  assign n725 = ( n721 & n723 ) | ( n721 & ~n724 ) | ( n723 & ~n724 ) ;
  assign n726 = ~n378 & n390 ;
  assign n727 = n378 & n390 ;
  assign n728 = ( n378 & n726 ) | ( n378 & ~n727 ) | ( n726 & ~n727 ) ;
  assign n729 = ( n384 & n725 ) | ( n384 & n728 ) | ( n725 & n728 ) ;
  assign n730 = ( n725 & n728 ) | ( n725 & ~n729 ) | ( n728 & ~n729 ) ;
  assign n731 = ( n384 & ~n729 ) | ( n384 & n730 ) | ( ~n729 & n730 ) ;
  assign n732 = n338 & ~n731 ;
  assign n733 = ~n338 & n731 ;
  assign n734 = n732 | n733 ;
  assign n735 = ~n344 & n350 ;
  assign n736 = n344 & n350 ;
  assign n737 = ( n344 & n735 ) | ( n344 & ~n736 ) | ( n735 & ~n736 ) ;
  assign n738 = ( n356 & n734 ) | ( n356 & n737 ) | ( n734 & n737 ) ;
  assign n739 = ( n734 & n737 ) | ( n734 & ~n738 ) | ( n737 & ~n738 ) ;
  assign n740 = ( n356 & ~n738 ) | ( n356 & n739 ) | ( ~n738 & n739 ) ;
  assign n741 = n362 & ~n740 ;
  assign n742 = ~n362 & n740 ;
  assign n743 = n741 | n742 ;
  assign n749 = n681 | n691 ;
  assign n750 = n570 | n749 ;
  assign n744 = x1 | n513 ;
  assign n745 = ( n457 & n513 ) | ( n457 & n744 ) | ( n513 & n744 ) ;
  assign n746 = n387 & ~n745 ;
  assign n747 = n387 & n745 ;
  assign n748 = ( n745 & n746 ) | ( n745 & ~n747 ) | ( n746 & ~n747 ) ;
  assign n751 = n668 | n748 ;
  assign n752 = ( ~n657 & n750 ) | ( ~n657 & n751 ) | ( n750 & n751 ) ;
  assign n753 = n657 | n752 ;
  assign n754 = n393 & n516 ;
  assign n767 = n515 | n754 ;
  assign n770 = ~n745 & n767 ;
  assign n768 = n393 | n767 ;
  assign n769 = ( n387 & n767 ) | ( n387 & n768 ) | ( n767 & n768 ) ;
  assign n771 = n745 & n769 ;
  assign n772 = ( ~n381 & n770 ) | ( ~n381 & n771 ) | ( n770 & n771 ) ;
  assign n773 = ( n381 & ~n771 ) | ( n381 & n772 ) | ( ~n771 & n772 ) ;
  assign n774 = ( ~n770 & n772 ) | ( ~n770 & n773 ) | ( n772 & n773 ) ;
  assign n755 = ( n514 & n515 ) | ( n514 & ~n754 ) | ( n515 & ~n754 ) ;
  assign n756 = n381 | n514 ;
  assign n757 = ( n754 & n755 ) | ( n754 & n756 ) | ( n755 & n756 ) ;
  assign n762 = ~n745 & n757 ;
  assign n758 = x139 & ~n384 ;
  assign n759 = ( n384 & n394 ) | ( n384 & n758 ) | ( n394 & n758 ) ;
  assign n760 = ( x142 & n378 ) | ( x142 & n515 ) | ( n378 & n515 ) ;
  assign n761 = n759 | n760 ;
  assign n763 = n745 & n761 ;
  assign n764 = ( ~n375 & n762 ) | ( ~n375 & n763 ) | ( n762 & n763 ) ;
  assign n765 = ( n375 & ~n763 ) | ( n375 & n764 ) | ( ~n763 & n764 ) ;
  assign n766 = ( ~n762 & n764 ) | ( ~n762 & n765 ) | ( n764 & n765 ) ;
  assign n775 = ( x139 & n384 ) | ( x139 & n745 ) | ( n384 & n745 ) ;
  assign n776 = n393 | n775 ;
  assign n777 = n393 & n775 ;
  assign n778 = n776 & ~n777 ;
  assign n779 = n766 | n778 ;
  assign n780 = ( ~n753 & n774 ) | ( ~n753 & n779 ) | ( n774 & n779 ) ;
  assign n781 = n753 | n780 ;
  assign n782 = n438 & ~n584 ;
  assign n783 = n438 & n584 ;
  assign n784 = ( n584 & n782 ) | ( n584 & ~n783 ) | ( n782 & ~n783 ) ;
  assign n785 = n552 & ~n561 ;
  assign n786 = ~n631 & n785 ;
  assign n787 = ~n784 & n786 ;
  assign n788 = ( n610 & n621 ) | ( n610 & n787 ) | ( n621 & n787 ) ;
  assign n789 = ~n610 & n788 ;
  assign n792 = n577 & ~n584 ;
  assign n790 = n438 | n577 ;
  assign n791 = ( n432 & n577 ) | ( n432 & n790 ) | ( n577 & n790 ) ;
  assign n793 = n584 & n791 ;
  assign n794 = ( ~n444 & n792 ) | ( ~n444 & n793 ) | ( n792 & n793 ) ;
  assign n795 = ( n444 & ~n793 ) | ( n444 & n794 ) | ( ~n793 & n794 ) ;
  assign n796 = ( ~n792 & n794 ) | ( ~n792 & n795 ) | ( n794 & n795 ) ;
  assign n797 = ( x145 & n435 ) | ( x145 & n584 ) | ( n435 & n584 ) ;
  assign n798 = n432 | n797 ;
  assign n799 = n432 & n797 ;
  assign n800 = n798 & ~n799 ;
  assign n801 = n589 & ~n800 ;
  assign n802 = ( ~n789 & n796 ) | ( ~n789 & n801 ) | ( n796 & n801 ) ;
  assign n803 = n789 & n802 ;
  assign n807 = ( ~x157 & x158 ) | ( ~x157 & n558 ) | ( x158 & n558 ) ;
  assign n808 = ( x157 & x158 ) | ( x157 & n576 ) | ( x158 & n576 ) ;
  assign n809 = n807 | n808 ;
  assign n804 = ( x80 & ~x157 ) | ( x80 & x158 ) | ( ~x157 & x158 ) ;
  assign n805 = ( x79 & x157 ) | ( x79 & x158 ) | ( x157 & x158 ) ;
  assign n806 = n804 & n805 ;
  assign n810 = x63 & n806 ;
  assign n811 = ( x63 & ~n809 ) | ( x63 & n810 ) | ( ~n809 & n810 ) ;
  assign n815 = ( ~x159 & x160 ) | ( ~x159 & n558 ) | ( x160 & n558 ) ;
  assign n816 = ( x159 & x160 ) | ( x159 & n576 ) | ( x160 & n576 ) ;
  assign n817 = n815 | n816 ;
  assign n812 = ( x80 & ~x159 ) | ( x80 & x160 ) | ( ~x159 & x160 ) ;
  assign n813 = ( x79 & x159 ) | ( x79 & x160 ) | ( x159 & x160 ) ;
  assign n814 = n812 & n813 ;
  assign n818 = x63 & n814 ;
  assign n819 = ( x63 & ~n817 ) | ( x63 & n818 ) | ( ~n817 & n818 ) ;
  assign n820 = ( x171 & ~x172 ) | ( x171 & n616 ) | ( ~x172 & n616 ) ;
  assign n821 = ( x171 & x172 ) | ( x171 & n663 ) | ( x172 & n663 ) ;
  assign n822 = n820 | n821 ;
  assign n823 = ( x13 & x171 ) | ( x13 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n824 = ( x15 & x171 ) | ( x15 & x172 ) | ( x171 & x172 ) ;
  assign n825 = n823 & n824 ;
  assign n826 = n822 & ~n825 ;
  assign n827 = ( x171 & ~x172 ) | ( x171 & n627 ) | ( ~x172 & n627 ) ;
  assign n828 = ( x171 & x172 ) | ( x171 & n674 ) | ( x172 & n674 ) ;
  assign n829 = n827 | n828 ;
  assign n830 = ( x5 & x171 ) | ( x5 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n831 = ( x26 & x171 ) | ( x26 & x172 ) | ( x171 & x172 ) ;
  assign n832 = n830 & n831 ;
  assign n833 = n829 & ~n832 ;
  assign n834 = ( x171 & ~x172 ) | ( x171 & n637 ) | ( ~x172 & n637 ) ;
  assign n835 = ( x171 & x172 ) | ( x171 & n687 ) | ( x172 & n687 ) ;
  assign n836 = n834 | n835 ;
  assign n837 = ( x4 & x171 ) | ( x4 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n838 = ( x25 & x171 ) | ( x25 & x172 ) | ( x171 & x172 ) ;
  assign n839 = n837 & n838 ;
  assign n840 = n836 & ~n839 ;
  assign n841 = ( x171 & ~x172 ) | ( x171 & n567 ) | ( ~x172 & n567 ) ;
  assign n842 = ( x171 & x172 ) | ( x171 & n697 ) | ( x172 & n697 ) ;
  assign n843 = n841 | n842 ;
  assign n844 = ( x24 & x171 ) | ( x24 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n845 = ( x23 & x171 ) | ( x23 & x172 ) | ( x171 & x172 ) ;
  assign n846 = n844 & n845 ;
  assign n847 = n843 & ~n846 ;
  assign n848 = ( ~x173 & x174 ) | ( ~x173 & n616 ) | ( x174 & n616 ) ;
  assign n849 = ( x173 & x174 ) | ( x173 & n663 ) | ( x174 & n663 ) ;
  assign n850 = n848 | n849 ;
  assign n851 = ( x13 & ~x173 ) | ( x13 & x174 ) | ( ~x173 & x174 ) ;
  assign n852 = ( x15 & x173 ) | ( x15 & x174 ) | ( x173 & x174 ) ;
  assign n853 = n851 & n852 ;
  assign n854 = n850 & ~n853 ;
  assign n855 = ( ~x173 & x174 ) | ( ~x173 & n627 ) | ( x174 & n627 ) ;
  assign n856 = ( x173 & x174 ) | ( x173 & n674 ) | ( x174 & n674 ) ;
  assign n857 = n855 | n856 ;
  assign n858 = ( x5 & ~x173 ) | ( x5 & x174 ) | ( ~x173 & x174 ) ;
  assign n859 = ( x26 & x173 ) | ( x26 & x174 ) | ( x173 & x174 ) ;
  assign n860 = n858 & n859 ;
  assign n861 = n857 & ~n860 ;
  assign n862 = ( ~x173 & x174 ) | ( ~x173 & n637 ) | ( x174 & n637 ) ;
  assign n863 = ( x173 & x174 ) | ( x173 & n687 ) | ( x174 & n687 ) ;
  assign n864 = n862 | n863 ;
  assign n865 = ( x4 & ~x173 ) | ( x4 & x174 ) | ( ~x173 & x174 ) ;
  assign n866 = ( x25 & x173 ) | ( x25 & x174 ) | ( x173 & x174 ) ;
  assign n867 = n865 & n866 ;
  assign n868 = n864 & ~n867 ;
  assign n869 = ( ~x173 & x174 ) | ( ~x173 & n567 ) | ( x174 & n567 ) ;
  assign n870 = ( x173 & x174 ) | ( x173 & n697 ) | ( x174 & n697 ) ;
  assign n871 = n869 | n870 ;
  assign n872 = ( x24 & ~x173 ) | ( x24 & x174 ) | ( ~x173 & x174 ) ;
  assign n873 = ( x23 & x173 ) | ( x23 & x174 ) | ( x173 & x174 ) ;
  assign n874 = n872 & n873 ;
  assign n875 = n871 & ~n874 ;
  assign n879 = ( ~x157 & x158 ) | ( ~x157 & n616 ) | ( x158 & n616 ) ;
  assign n880 = ( x157 & x158 ) | ( x157 & n663 ) | ( x158 & n663 ) ;
  assign n881 = n879 | n880 ;
  assign n876 = ( x75 & ~x157 ) | ( x75 & x158 ) | ( ~x157 & x158 ) ;
  assign n877 = ( x85 & x157 ) | ( x85 & x158 ) | ( x157 & x158 ) ;
  assign n878 = n876 & n877 ;
  assign n882 = x63 & n878 ;
  assign n883 = ( x63 & ~n881 ) | ( x63 & n882 ) | ( ~n881 & n882 ) ;
  assign n887 = ( ~x157 & x158 ) | ( ~x157 & n567 ) | ( x158 & n567 ) ;
  assign n888 = ( x157 & x158 ) | ( x157 & n697 ) | ( x158 & n697 ) ;
  assign n889 = n887 | n888 ;
  assign n884 = ( x71 & ~x157 ) | ( x71 & x158 ) | ( ~x157 & x158 ) ;
  assign n885 = ( x81 & x157 ) | ( x81 & x158 ) | ( x157 & x158 ) ;
  assign n886 = n884 & n885 ;
  assign n890 = x63 & n886 ;
  assign n891 = ( x63 & ~n889 ) | ( x63 & n890 ) | ( ~n889 & n890 ) ;
  assign n895 = ( ~x157 & x158 ) | ( ~x157 & n637 ) | ( x158 & n637 ) ;
  assign n896 = ( x157 & x158 ) | ( x157 & n687 ) | ( x158 & n687 ) ;
  assign n897 = n895 | n896 ;
  assign n892 = ( x69 & ~x157 ) | ( x69 & x158 ) | ( ~x157 & x158 ) ;
  assign n893 = ( x70 & x157 ) | ( x70 & x158 ) | ( x157 & x158 ) ;
  assign n894 = n892 & n893 ;
  assign n898 = x63 & n894 ;
  assign n899 = ( x63 & ~n897 ) | ( x63 & n898 ) | ( ~n897 & n898 ) ;
  assign n903 = ( ~x157 & x158 ) | ( ~x157 & n627 ) | ( x158 & n627 ) ;
  assign n904 = ( x157 & x158 ) | ( x157 & n674 ) | ( x158 & n674 ) ;
  assign n905 = n903 | n904 ;
  assign n900 = ( x67 & ~x157 ) | ( x67 & x158 ) | ( ~x157 & x158 ) ;
  assign n901 = ( x68 & x157 ) | ( x68 & x158 ) | ( x157 & x158 ) ;
  assign n902 = n900 & n901 ;
  assign n906 = x63 & n902 ;
  assign n907 = ( x63 & ~n905 ) | ( x63 & n906 ) | ( ~n905 & n906 ) ;
  assign n911 = ( ~x159 & x160 ) | ( ~x159 & n616 ) | ( x160 & n616 ) ;
  assign n912 = ( x159 & x160 ) | ( x159 & n663 ) | ( x160 & n663 ) ;
  assign n913 = n911 | n912 ;
  assign n908 = ( x75 & ~x159 ) | ( x75 & x160 ) | ( ~x159 & x160 ) ;
  assign n909 = ( x85 & x159 ) | ( x85 & x160 ) | ( x159 & x160 ) ;
  assign n910 = n908 & n909 ;
  assign n914 = x63 & n910 ;
  assign n915 = ( x63 & ~n913 ) | ( x63 & n914 ) | ( ~n913 & n914 ) ;
  assign n919 = ( ~x159 & x160 ) | ( ~x159 & n567 ) | ( x160 & n567 ) ;
  assign n920 = ( x159 & x160 ) | ( x159 & n697 ) | ( x160 & n697 ) ;
  assign n921 = n919 | n920 ;
  assign n916 = ( x71 & ~x159 ) | ( x71 & x160 ) | ( ~x159 & x160 ) ;
  assign n917 = ( x81 & x159 ) | ( x81 & x160 ) | ( x159 & x160 ) ;
  assign n918 = n916 & n917 ;
  assign n922 = x63 & n918 ;
  assign n923 = ( x63 & ~n921 ) | ( x63 & n922 ) | ( ~n921 & n922 ) ;
  assign n927 = ( ~x159 & x160 ) | ( ~x159 & n637 ) | ( x160 & n637 ) ;
  assign n928 = ( x159 & x160 ) | ( x159 & n687 ) | ( x160 & n687 ) ;
  assign n929 = n927 | n928 ;
  assign n924 = ( x69 & ~x159 ) | ( x69 & x160 ) | ( ~x159 & x160 ) ;
  assign n925 = ( x70 & x159 ) | ( x70 & x160 ) | ( x159 & x160 ) ;
  assign n926 = n924 & n925 ;
  assign n930 = x63 & n926 ;
  assign n931 = ( x63 & ~n929 ) | ( x63 & n930 ) | ( ~n929 & n930 ) ;
  assign n935 = ( ~x159 & x160 ) | ( ~x159 & n627 ) | ( x160 & n627 ) ;
  assign n936 = ( x159 & x160 ) | ( x159 & n674 ) | ( x160 & n674 ) ;
  assign n937 = n935 | n936 ;
  assign n932 = ( x67 & ~x159 ) | ( x67 & x160 ) | ( ~x159 & x160 ) ;
  assign n933 = ( x68 & x159 ) | ( x68 & x160 ) | ( x159 & x160 ) ;
  assign n934 = n932 & n933 ;
  assign n938 = x63 & n934 ;
  assign n939 = ( x63 & ~n937 ) | ( x63 & n938 ) | ( ~n937 & n938 ) ;
  assign n940 = ( ~x169 & x170 ) | ( ~x169 & n589 ) | ( x170 & n589 ) ;
  assign n941 = ( x53 & x169 ) | ( x53 & x170 ) | ( x169 & x170 ) ;
  assign n942 = ~n940 & n941 ;
  assign n946 = ( ~x169 & x170 ) | ( ~x169 & n259 ) | ( x170 & n259 ) ;
  assign n943 = x60 | n441 ;
  assign n944 = ~x60 & n441 ;
  assign n945 = ( ~n441 & n943 ) | ( ~n441 & n944 ) | ( n943 & n944 ) ;
  assign n947 = ( x169 & x170 ) | ( x169 & n945 ) | ( x170 & n945 ) ;
  assign n948 = n946 & ~n947 ;
  assign n949 = n942 | n948 ;
  assign n950 = ~x177 & n949 ;
  assign n951 = ( ~x61 & n949 ) | ( ~x61 & n950 ) | ( n949 & n950 ) ;
  assign n952 = n589 & ~n945 ;
  assign n953 = n589 | n945 ;
  assign n954 = ( ~n589 & n952 ) | ( ~n589 & n953 ) | ( n952 & n953 ) ;
  assign n955 = ( x175 & ~x176 ) | ( x175 & n259 ) | ( ~x176 & n259 ) ;
  assign n956 = ( x175 & x176 ) | ( x175 & n589 ) | ( x176 & n589 ) ;
  assign n957 = n955 & ~n956 ;
  assign n958 = ( x53 & ~x175 ) | ( x53 & n957 ) | ( ~x175 & n957 ) ;
  assign n959 = x176 & ~n958 ;
  assign n960 = ( x176 & n957 ) | ( x176 & ~n959 ) | ( n957 & ~n959 ) ;
  assign n961 = ( ~x175 & x176 ) | ( ~x175 & n256 ) | ( x176 & n256 ) ;
  assign n962 = ( x175 & x176 ) | ( x175 & n796 ) | ( x176 & n796 ) ;
  assign n963 = n961 | n962 ;
  assign n964 = ( ~x51 & x175 ) | ( ~x51 & n963 ) | ( x175 & n963 ) ;
  assign n965 = x176 & n964 ;
  assign n966 = ( ~x176 & n963 ) | ( ~x176 & n965 ) | ( n963 & n965 ) ;
  assign n967 = ( x175 & ~x176 ) | ( x175 & n253 ) | ( ~x176 & n253 ) ;
  assign n968 = ( x175 & x176 ) | ( x175 & ~n800 ) | ( x176 & ~n800 ) ;
  assign n969 = n967 & ~n968 ;
  assign n970 = ( x46 & ~x175 ) | ( x46 & n969 ) | ( ~x175 & n969 ) ;
  assign n971 = x176 & ~n970 ;
  assign n972 = ( x176 & n969 ) | ( x176 & ~n971 ) | ( n969 & ~n971 ) ;
  assign n973 = ( x175 & ~x176 ) | ( x175 & n246 ) | ( ~x176 & n246 ) ;
  assign n974 = ( x175 & x176 ) | ( x175 & ~n784 ) | ( x176 & ~n784 ) ;
  assign n975 = n973 & ~n974 ;
  assign n976 = ( x42 & ~x175 ) | ( x42 & n975 ) | ( ~x175 & n975 ) ;
  assign n977 = x176 & ~n976 ;
  assign n978 = ( x176 & n975 ) | ( x176 & ~n977 ) | ( n975 & ~n977 ) ;
  assign n982 = x152 & x154 ;
  assign n983 = ( ~x135 & x153 ) | ( ~x135 & n982 ) | ( x153 & n982 ) ;
  assign n984 = x135 & n983 ;
  assign n979 = x155 & ~n743 ;
  assign n980 = ( n476 & ~n720 ) | ( n476 & n979 ) | ( ~n720 & n979 ) ;
  assign n981 = n720 & n980 ;
  assign n985 = x98 & n981 ;
  assign n986 = ( n497 & n984 ) | ( n497 & n985 ) | ( n984 & n985 ) ;
  assign n987 = ~n497 & n986 ;
  assign n988 = ( x175 & ~x176 ) | ( x175 & n271 ) | ( ~x176 & n271 ) ;
  assign n989 = ( x175 & x176 ) | ( x175 & ~n766 ) | ( x176 & ~n766 ) ;
  assign n990 = n988 & ~n989 ;
  assign n991 = ( x45 & ~x175 ) | ( x45 & n990 ) | ( ~x175 & n990 ) ;
  assign n992 = x176 & ~n991 ;
  assign n993 = ( x176 & n990 ) | ( x176 & ~n992 ) | ( n990 & ~n992 ) ;
  assign n994 = ( ~x175 & x176 ) | ( ~x175 & n309 ) | ( x176 & n309 ) ;
  assign n995 = ( x175 & x176 ) | ( x175 & ~n774 ) | ( x176 & ~n774 ) ;
  assign n996 = n994 | n995 ;
  assign n997 = ( ~x44 & x175 ) | ( ~x44 & n996 ) | ( x175 & n996 ) ;
  assign n998 = x176 & n997 ;
  assign n999 = ( ~x176 & n996 ) | ( ~x176 & n998 ) | ( n996 & n998 ) ;
  assign n1000 = ( ~x175 & x176 ) | ( ~x175 & n316 ) | ( x176 & n316 ) ;
  assign n1001 = ( x175 & x176 ) | ( x175 & ~n778 ) | ( x176 & ~n778 ) ;
  assign n1002 = n1000 | n1001 ;
  assign n1003 = ( ~x19 & x175 ) | ( ~x19 & n1002 ) | ( x175 & n1002 ) ;
  assign n1004 = x176 & n1003 ;
  assign n1005 = ( ~x176 & n1002 ) | ( ~x176 & n1004 ) | ( n1002 & n1004 ) ;
  assign n1006 = ( ~x175 & x176 ) | ( ~x175 & n330 ) | ( x176 & n330 ) ;
  assign n1007 = ( x175 & x176 ) | ( x175 & ~n748 ) | ( x176 & ~n748 ) ;
  assign n1008 = n1006 | n1007 ;
  assign n1009 = ( ~x43 & x175 ) | ( ~x43 & n1008 ) | ( x175 & n1008 ) ;
  assign n1010 = x176 & n1009 ;
  assign n1011 = ( ~x176 & n1008 ) | ( ~x176 & n1010 ) | ( n1008 & n1010 ) ;
  assign n1012 = ( x173 & ~x174 ) | ( x173 & n960 ) | ( ~x174 & n960 ) ;
  assign n1013 = ( x173 & x174 ) | ( x173 & ~n993 ) | ( x174 & ~n993 ) ;
  assign n1014 = n1012 & ~n1013 ;
  assign n1015 = ( x40 & ~x173 ) | ( x40 & x174 ) | ( ~x173 & x174 ) ;
  assign n1016 = ( x41 & x173 ) | ( x41 & x174 ) | ( x173 & x174 ) ;
  assign n1017 = n1015 & n1016 ;
  assign n1018 = n1014 | n1017 ;
  assign n1019 = ( ~x171 & x172 ) | ( ~x171 & n960 ) | ( x172 & n960 ) ;
  assign n1020 = ( x171 & x172 ) | ( x171 & ~n993 ) | ( x172 & ~n993 ) ;
  assign n1021 = n1019 & ~n1020 ;
  assign n1022 = ( x40 & x171 ) | ( x40 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n1023 = ( x41 & x171 ) | ( x41 & x172 ) | ( x171 & x172 ) ;
  assign n1024 = n1022 & n1023 ;
  assign n1025 = n1021 | n1024 ;
  assign n1026 = ( x171 & ~x172 ) | ( x171 & n966 ) | ( ~x172 & n966 ) ;
  assign n1027 = ( x171 & x172 ) | ( x171 & n999 ) | ( x172 & n999 ) ;
  assign n1028 = n1026 | n1027 ;
  assign n1029 = ( x17 & x171 ) | ( x17 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n1030 = ( x16 & x171 ) | ( x16 & x172 ) | ( x171 & x172 ) ;
  assign n1031 = n1029 & n1030 ;
  assign n1032 = n1028 & ~n1031 ;
  assign n1033 = ( ~x171 & x172 ) | ( ~x171 & n972 ) | ( x172 & n972 ) ;
  assign n1034 = ( x171 & x172 ) | ( x171 & n1005 ) | ( x172 & n1005 ) ;
  assign n1035 = n1033 & ~n1034 ;
  assign n1036 = ( x39 & x171 ) | ( x39 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n1037 = ( x38 & x171 ) | ( x38 & x172 ) | ( x171 & x172 ) ;
  assign n1038 = n1036 & n1037 ;
  assign n1039 = n1035 | n1038 ;
  assign n1040 = ( ~x171 & x172 ) | ( ~x171 & n978 ) | ( x172 & n978 ) ;
  assign n1041 = ( x171 & x172 ) | ( x171 & n1011 ) | ( x172 & n1011 ) ;
  assign n1042 = n1040 & ~n1041 ;
  assign n1043 = ( x14 & x171 ) | ( x14 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n1044 = ( x35 & x171 ) | ( x35 & x172 ) | ( x171 & x172 ) ;
  assign n1045 = n1043 & n1044 ;
  assign n1046 = n1042 | n1045 ;
  assign n1047 = ( ~x173 & x174 ) | ( ~x173 & n966 ) | ( x174 & n966 ) ;
  assign n1048 = ( x173 & x174 ) | ( x173 & n999 ) | ( x174 & n999 ) ;
  assign n1049 = n1047 | n1048 ;
  assign n1050 = ( x17 & ~x173 ) | ( x17 & x174 ) | ( ~x173 & x174 ) ;
  assign n1051 = ( x16 & x173 ) | ( x16 & x174 ) | ( x173 & x174 ) ;
  assign n1052 = n1050 & n1051 ;
  assign n1053 = n1049 & ~n1052 ;
  assign n1054 = ( x173 & ~x174 ) | ( x173 & n972 ) | ( ~x174 & n972 ) ;
  assign n1055 = ( x173 & x174 ) | ( x173 & n1005 ) | ( x174 & n1005 ) ;
  assign n1056 = n1054 & ~n1055 ;
  assign n1057 = ( x39 & ~x173 ) | ( x39 & x174 ) | ( ~x173 & x174 ) ;
  assign n1058 = ( x38 & x173 ) | ( x38 & x174 ) | ( x173 & x174 ) ;
  assign n1059 = n1057 & n1058 ;
  assign n1060 = n1056 | n1059 ;
  assign n1061 = ( x173 & ~x174 ) | ( x173 & n978 ) | ( ~x174 & n978 ) ;
  assign n1062 = ( x173 & x174 ) | ( x173 & n1011 ) | ( x174 & n1011 ) ;
  assign n1063 = n1061 & ~n1062 ;
  assign n1064 = ( x14 & ~x173 ) | ( x14 & x174 ) | ( ~x173 & x174 ) ;
  assign n1065 = ( x35 & x173 ) | ( x35 & x174 ) | ( x173 & x174 ) ;
  assign n1066 = n1064 & n1065 ;
  assign n1067 = n1063 | n1066 ;
  assign n1071 = ( x157 & ~x158 ) | ( x157 & n978 ) | ( ~x158 & n978 ) ;
  assign n1072 = ( x157 & x158 ) | ( x157 & n1011 ) | ( x158 & n1011 ) ;
  assign n1073 = n1071 & ~n1072 ;
  assign n1068 = ( x76 & ~x157 ) | ( x76 & x158 ) | ( ~x157 & x158 ) ;
  assign n1069 = ( x86 & x157 ) | ( x86 & x158 ) | ( x157 & x158 ) ;
  assign n1070 = n1068 & n1069 ;
  assign n1074 = x63 & n1070 ;
  assign n1075 = ( x63 & n1073 ) | ( x63 & n1074 ) | ( n1073 & n1074 ) ;
  assign n1079 = ( x157 & ~x158 ) | ( x157 & n972 ) | ( ~x158 & n972 ) ;
  assign n1080 = ( x157 & x158 ) | ( x157 & n1005 ) | ( x158 & n1005 ) ;
  assign n1081 = n1079 & ~n1080 ;
  assign n1076 = ( x74 & ~x157 ) | ( x74 & x158 ) | ( ~x157 & x158 ) ;
  assign n1077 = ( x84 & x157 ) | ( x84 & x158 ) | ( x157 & x158 ) ;
  assign n1078 = n1076 & n1077 ;
  assign n1082 = x63 & n1078 ;
  assign n1083 = ( x63 & n1081 ) | ( x63 & n1082 ) | ( n1081 & n1082 ) ;
  assign n1087 = ( ~x157 & x158 ) | ( ~x157 & n966 ) | ( x158 & n966 ) ;
  assign n1088 = ( x157 & x158 ) | ( x157 & n999 ) | ( x158 & n999 ) ;
  assign n1089 = n1087 | n1088 ;
  assign n1084 = ( x73 & ~x157 ) | ( x73 & x158 ) | ( ~x157 & x158 ) ;
  assign n1085 = ( x83 & x157 ) | ( x83 & x158 ) | ( x157 & x158 ) ;
  assign n1086 = n1084 & n1085 ;
  assign n1090 = x63 & n1086 ;
  assign n1091 = ( x63 & ~n1089 ) | ( x63 & n1090 ) | ( ~n1089 & n1090 ) ;
  assign n1095 = ( x157 & ~x158 ) | ( x157 & n960 ) | ( ~x158 & n960 ) ;
  assign n1096 = ( x157 & x158 ) | ( x157 & ~n993 ) | ( x158 & ~n993 ) ;
  assign n1097 = n1095 & ~n1096 ;
  assign n1092 = ( x72 & ~x157 ) | ( x72 & x158 ) | ( ~x157 & x158 ) ;
  assign n1093 = ( x82 & x157 ) | ( x82 & x158 ) | ( x157 & x158 ) ;
  assign n1094 = n1092 & n1093 ;
  assign n1098 = x63 & n1094 ;
  assign n1099 = ( x63 & n1097 ) | ( x63 & n1098 ) | ( n1097 & n1098 ) ;
  assign n1103 = ( x159 & ~x160 ) | ( x159 & n978 ) | ( ~x160 & n978 ) ;
  assign n1104 = ( x159 & x160 ) | ( x159 & n1011 ) | ( x160 & n1011 ) ;
  assign n1105 = n1103 & ~n1104 ;
  assign n1100 = ( x76 & ~x159 ) | ( x76 & x160 ) | ( ~x159 & x160 ) ;
  assign n1101 = ( x86 & x159 ) | ( x86 & x160 ) | ( x159 & x160 ) ;
  assign n1102 = n1100 & n1101 ;
  assign n1106 = x63 & n1102 ;
  assign n1107 = ( x63 & n1105 ) | ( x63 & n1106 ) | ( n1105 & n1106 ) ;
  assign n1111 = ( x159 & ~x160 ) | ( x159 & n972 ) | ( ~x160 & n972 ) ;
  assign n1112 = ( x159 & x160 ) | ( x159 & n1005 ) | ( x160 & n1005 ) ;
  assign n1113 = n1111 & ~n1112 ;
  assign n1108 = ( x74 & ~x159 ) | ( x74 & x160 ) | ( ~x159 & x160 ) ;
  assign n1109 = ( x84 & x159 ) | ( x84 & x160 ) | ( x159 & x160 ) ;
  assign n1110 = n1108 & n1109 ;
  assign n1114 = x63 & n1110 ;
  assign n1115 = ( x63 & n1113 ) | ( x63 & n1114 ) | ( n1113 & n1114 ) ;
  assign n1119 = ( ~x159 & x160 ) | ( ~x159 & n966 ) | ( x160 & n966 ) ;
  assign n1120 = ( x159 & x160 ) | ( x159 & n999 ) | ( x160 & n999 ) ;
  assign n1121 = n1119 | n1120 ;
  assign n1116 = ( x73 & ~x159 ) | ( x73 & x160 ) | ( ~x159 & x160 ) ;
  assign n1117 = ( x83 & x159 ) | ( x83 & x160 ) | ( x159 & x160 ) ;
  assign n1118 = n1116 & n1117 ;
  assign n1122 = x63 & n1118 ;
  assign n1123 = ( x63 & ~n1121 ) | ( x63 & n1122 ) | ( ~n1121 & n1122 ) ;
  assign n1127 = ( x159 & ~x160 ) | ( x159 & n960 ) | ( ~x160 & n960 ) ;
  assign n1128 = ( x159 & x160 ) | ( x159 & ~n993 ) | ( x160 & ~n993 ) ;
  assign n1129 = n1127 & ~n1128 ;
  assign n1124 = ( x72 & ~x159 ) | ( x72 & x160 ) | ( ~x159 & x160 ) ;
  assign n1125 = ( x82 & x159 ) | ( x82 & x160 ) | ( x159 & x160 ) ;
  assign n1126 = n1124 & n1125 ;
  assign n1130 = x63 & n1126 ;
  assign n1131 = ( x63 & n1129 ) | ( x63 & n1130 ) | ( n1129 & n1130 ) ;
  assign n1160 = ( x99 & ~x125 ) | ( x99 & x148 ) | ( ~x125 & x148 ) ;
  assign n1161 = ( x100 & x125 ) | ( x100 & x148 ) | ( x125 & x148 ) ;
  assign n1162 = n1160 & n1161 ;
  assign n1151 = ( x99 & ~x127 ) | ( x99 & x149 ) | ( ~x127 & x149 ) ;
  assign n1152 = ( x100 & x127 ) | ( x100 & x149 ) | ( x127 & x149 ) ;
  assign n1153 = n1151 & n1152 ;
  assign n1157 = ( x101 & ~x127 ) | ( x101 & x149 ) | ( ~x127 & x149 ) ;
  assign n1158 = ( x97 & x127 ) | ( x97 & x149 ) | ( x127 & x149 ) ;
  assign n1159 = n1157 | n1158 ;
  assign n1163 = ~n1153 & n1159 ;
  assign n1164 = n1162 & ~n1163 ;
  assign n1154 = ( x101 & ~x125 ) | ( x101 & x148 ) | ( ~x125 & x148 ) ;
  assign n1155 = ( x97 & x125 ) | ( x97 & x148 ) | ( x125 & x148 ) ;
  assign n1156 = n1154 | n1155 ;
  assign n1165 = n1156 & ~n1163 ;
  assign n1166 = ( ~n1156 & n1162 ) | ( ~n1156 & n1163 ) | ( n1162 & n1163 ) ;
  assign n1167 = ( ~n1164 & n1165 ) | ( ~n1164 & n1166 ) | ( n1165 & n1166 ) ;
  assign n1132 = ( n246 & n253 ) | ( n246 & ~n259 ) | ( n253 & ~n259 ) ;
  assign n1133 = ( n246 & n253 ) | ( n246 & ~n1132 ) | ( n253 & ~n1132 ) ;
  assign n1134 = ( n259 & n1132 ) | ( n259 & ~n1133 ) | ( n1132 & ~n1133 ) ;
  assign n1135 = n256 & ~n1134 ;
  assign n1136 = ~n256 & n1134 ;
  assign n1137 = n1135 | n1136 ;
  assign n1138 = ( x101 & ~x120 ) | ( x101 & x146 ) | ( ~x120 & x146 ) ;
  assign n1139 = ( x97 & x120 ) | ( x97 & x146 ) | ( x120 & x146 ) ;
  assign n1140 = n1138 | n1139 ;
  assign n1144 = x99 & x147 ;
  assign n1145 = x97 & ~x147 ;
  assign n1146 = ( x147 & ~n1144 ) | ( x147 & n1145 ) | ( ~n1144 & n1145 ) ;
  assign n1141 = ( x99 & ~x120 ) | ( x99 & x146 ) | ( ~x120 & x146 ) ;
  assign n1142 = ( x100 & x120 ) | ( x100 & x146 ) | ( x120 & x146 ) ;
  assign n1143 = n1141 & n1142 ;
  assign n1147 = n1140 & n1143 ;
  assign n1148 = ( n1140 & n1146 ) | ( n1140 & n1147 ) | ( n1146 & n1147 ) ;
  assign n1149 = ( ~n1140 & n1146 ) | ( ~n1140 & n1147 ) | ( n1146 & n1147 ) ;
  assign n1150 = ( n1140 & ~n1148 ) | ( n1140 & n1149 ) | ( ~n1148 & n1149 ) ;
  assign n1168 = ( ~n1137 & n1150 ) | ( ~n1137 & n1167 ) | ( n1150 & n1167 ) ;
  assign n1169 = ( n1137 & ~n1150 ) | ( n1137 & n1168 ) | ( ~n1150 & n1168 ) ;
  assign n1170 = ( ~n1167 & n1168 ) | ( ~n1167 & n1169 ) | ( n1168 & n1169 ) ;
  assign n1171 = n212 & n1170 ;
  assign n1172 = n212 | n1170 ;
  assign n1173 = ~n1171 & n1172 ;
  assign n1243 = ( x175 & ~x176 ) | ( x175 & n1173 ) | ( ~x176 & n1173 ) ;
  assign n1193 = ( ~n436 & n577 ) | ( ~n436 & n578 ) | ( n577 & n578 ) ;
  assign n1194 = ( n436 & ~n578 ) | ( n436 & n1193 ) | ( ~n578 & n1193 ) ;
  assign n1195 = ( ~n577 & n1193 ) | ( ~n577 & n1194 ) | ( n1193 & n1194 ) ;
  assign n1196 = ( n432 & n441 ) | ( n432 & n1195 ) | ( n441 & n1195 ) ;
  assign n1197 = ( n432 & n1195 ) | ( n432 & ~n1196 ) | ( n1195 & ~n1196 ) ;
  assign n1198 = ( n441 & ~n1196 ) | ( n441 & n1197 ) | ( ~n1196 & n1197 ) ;
  assign n1199 = n444 & ~n1198 ;
  assign n1200 = ~n444 & n1198 ;
  assign n1201 = n1199 | n1200 ;
  assign n1214 = n452 | n540 ;
  assign n1215 = ( x161 & n1201 ) | ( x161 & n1214 ) | ( n1201 & n1214 ) ;
  assign n1202 = ( n541 & n582 ) | ( n541 & n791 ) | ( n582 & n791 ) ;
  assign n1203 = ( n541 & n582 ) | ( n541 & ~n1202 ) | ( n582 & ~n1202 ) ;
  assign n1204 = ( n791 & ~n1202 ) | ( n791 & n1203 ) | ( ~n1202 & n1203 ) ;
  assign n1205 = ( n432 & n441 ) | ( n432 & ~n1204 ) | ( n441 & ~n1204 ) ;
  assign n1206 = ( ~n432 & n1204 ) | ( ~n432 & n1205 ) | ( n1204 & n1205 ) ;
  assign n1207 = ( ~n441 & n1205 ) | ( ~n441 & n1206 ) | ( n1205 & n1206 ) ;
  assign n1208 = n444 & n1207 ;
  assign n1209 = n444 | n1207 ;
  assign n1210 = ~n1208 & n1209 ;
  assign n1216 = ( ~x161 & n1210 ) | ( ~x161 & n1214 ) | ( n1210 & n1214 ) ;
  assign n1217 = n1215 & ~n1216 ;
  assign n1175 = n598 | n603 ;
  assign n1176 = ( x149 & ~n400 ) | ( x149 & n1175 ) | ( ~n400 & n1175 ) ;
  assign n1177 = ( x149 & n422 ) | ( x149 & ~n1176 ) | ( n422 & ~n1176 ) ;
  assign n1178 = ( n400 & n422 ) | ( n400 & n1176 ) | ( n422 & n1176 ) ;
  assign n1179 = ( n1175 & n1177 ) | ( n1175 & ~n1178 ) | ( n1177 & ~n1178 ) ;
  assign n1174 = ~n419 & n598 ;
  assign n1180 = n604 | n1174 ;
  assign n1181 = ( n422 & n1179 ) | ( n422 & ~n1180 ) | ( n1179 & ~n1180 ) ;
  assign n1182 = ( ~n1179 & n1180 ) | ( ~n1179 & n1181 ) | ( n1180 & n1181 ) ;
  assign n1183 = ( ~n422 & n1181 ) | ( ~n422 & n1182 ) | ( n1181 & n1182 ) ;
  assign n1184 = ( n403 & n409 ) | ( n403 & n1183 ) | ( n409 & n1183 ) ;
  assign n1185 = ( n403 & n1183 ) | ( n403 & ~n1184 ) | ( n1183 & ~n1184 ) ;
  assign n1186 = ( n409 & ~n1184 ) | ( n409 & n1185 ) | ( ~n1184 & n1185 ) ;
  assign n1187 = n415 & ~n1186 ;
  assign n1188 = ~n415 & n1186 ;
  assign n1189 = n1187 | n1188 ;
  assign n1190 = ( ~x161 & n419 ) | ( ~x161 & n1189 ) | ( n419 & n1189 ) ;
  assign n1191 = ~n419 & n1190 ;
  assign n1192 = ( ~n1189 & n1190 ) | ( ~n1189 & n1191 ) | ( n1190 & n1191 ) ;
  assign n1220 = n415 | n603 ;
  assign n1221 = ( n403 & n603 ) | ( n403 & n1220 ) | ( n603 & n1220 ) ;
  assign n1222 = ( x149 & ~n402 ) | ( x149 & n1221 ) | ( ~n402 & n1221 ) ;
  assign n1223 = ( x149 & n402 ) | ( x149 & ~n1221 ) | ( n402 & ~n1221 ) ;
  assign n1224 = ( ~x149 & n1222 ) | ( ~x149 & n1223 ) | ( n1222 & n1223 ) ;
  assign n1218 = n403 & n415 ;
  assign n1219 = ~n419 & n1218 ;
  assign n1225 = n604 | n1219 ;
  assign n1226 = ( n422 & n1224 ) | ( n422 & ~n1225 ) | ( n1224 & ~n1225 ) ;
  assign n1227 = ( ~n1224 & n1225 ) | ( ~n1224 & n1226 ) | ( n1225 & n1226 ) ;
  assign n1228 = ( ~n422 & n1226 ) | ( ~n422 & n1227 ) | ( n1226 & n1227 ) ;
  assign n1229 = ( n403 & n409 ) | ( n403 & ~n1228 ) | ( n409 & ~n1228 ) ;
  assign n1230 = ( ~n403 & n1228 ) | ( ~n403 & n1229 ) | ( n1228 & n1229 ) ;
  assign n1231 = ( ~n409 & n1229 ) | ( ~n409 & n1230 ) | ( n1229 & n1230 ) ;
  assign n1232 = n415 & n1231 ;
  assign n1233 = n415 | n1231 ;
  assign n1234 = ~n1232 & n1233 ;
  assign n1235 = ( x161 & n419 ) | ( x161 & n1234 ) | ( n419 & n1234 ) ;
  assign n1236 = ~n419 & n1235 ;
  assign n1237 = ( ~n1234 & n1235 ) | ( ~n1234 & n1236 ) | ( n1235 & n1236 ) ;
  assign n1238 = n1192 | n1237 ;
  assign n1239 = n1217 & n1238 ;
  assign n1211 = ( x161 & n540 ) | ( x161 & n1210 ) | ( n540 & n1210 ) ;
  assign n1212 = ( ~x161 & n540 ) | ( ~x161 & n1201 ) | ( n540 & n1201 ) ;
  assign n1213 = ~n1211 & n1212 ;
  assign n1240 = ~n1213 & n1238 ;
  assign n1241 = ( n1213 & n1217 ) | ( n1213 & ~n1238 ) | ( n1217 & ~n1238 ) ;
  assign n1242 = ( ~n1239 & n1240 ) | ( ~n1239 & n1241 ) | ( n1240 & n1241 ) ;
  assign n1244 = ( x175 & x176 ) | ( x175 & ~n1242 ) | ( x176 & ~n1242 ) ;
  assign n1245 = n1243 & ~n1244 ;
  assign n1246 = ( ~x50 & x175 ) | ( ~x50 & n1245 ) | ( x175 & n1245 ) ;
  assign n1247 = x176 | n1245 ;
  assign n1248 = ( x50 & n1246 ) | ( x50 & n1247 ) | ( n1246 & n1247 ) ;
  assign n1309 = ( x99 & ~x104 ) | ( x99 & x137 ) | ( ~x104 & x137 ) ;
  assign n1310 = ( x100 & x104 ) | ( x100 & x137 ) | ( x104 & x137 ) ;
  assign n1311 = n1309 & n1310 ;
  assign n1300 = ( x99 & ~x106 ) | ( x99 & x138 ) | ( ~x106 & x138 ) ;
  assign n1301 = ( x100 & x106 ) | ( x100 & x138 ) | ( x106 & x138 ) ;
  assign n1302 = n1300 & n1301 ;
  assign n1306 = ( x101 & ~x106 ) | ( x101 & x138 ) | ( ~x106 & x138 ) ;
  assign n1307 = ( x97 & x106 ) | ( x97 & x138 ) | ( x106 & x138 ) ;
  assign n1308 = n1306 | n1307 ;
  assign n1312 = ~n1302 & n1308 ;
  assign n1313 = n1311 & ~n1312 ;
  assign n1303 = ( x101 & ~x104 ) | ( x101 & x137 ) | ( ~x104 & x137 ) ;
  assign n1304 = ( x97 & x104 ) | ( x97 & x137 ) | ( x104 & x137 ) ;
  assign n1305 = n1303 | n1304 ;
  assign n1314 = n1305 & ~n1312 ;
  assign n1315 = ( ~n1305 & n1311 ) | ( ~n1305 & n1312 ) | ( n1311 & n1312 ) ;
  assign n1316 = ( ~n1313 & n1314 ) | ( ~n1313 & n1315 ) | ( n1314 & n1315 ) ;
  assign n1293 = ( x101 & ~x108 ) | ( x101 & x134 ) | ( ~x108 & x134 ) ;
  assign n1294 = ( x97 & x108 ) | ( x97 & x134 ) | ( x108 & x134 ) ;
  assign n1295 = n1293 | n1294 ;
  assign n1296 = ( x99 & ~x108 ) | ( x99 & x134 ) | ( ~x108 & x134 ) ;
  assign n1297 = ( x100 & x108 ) | ( x100 & x134 ) | ( x108 & x134 ) ;
  assign n1298 = n1296 & n1297 ;
  assign n1299 = n1295 & ~n1298 ;
  assign n1264 = ( ~x91 & x99 ) | ( ~x91 & x143 ) | ( x99 & x143 ) ;
  assign n1265 = ( x91 & x100 ) | ( x91 & x143 ) | ( x100 & x143 ) ;
  assign n1266 = n1264 & n1265 ;
  assign n1255 = ( ~x93 & x99 ) | ( ~x93 & x139 ) | ( x99 & x139 ) ;
  assign n1256 = ( x93 & x100 ) | ( x93 & x139 ) | ( x100 & x139 ) ;
  assign n1257 = n1255 & n1256 ;
  assign n1261 = ( ~x93 & x101 ) | ( ~x93 & x139 ) | ( x101 & x139 ) ;
  assign n1262 = ( x93 & x97 ) | ( x93 & x139 ) | ( x97 & x139 ) ;
  assign n1263 = n1261 | n1262 ;
  assign n1267 = ~n1257 & n1263 ;
  assign n1268 = n1266 & ~n1267 ;
  assign n1258 = ( ~x91 & x101 ) | ( ~x91 & x143 ) | ( x101 & x143 ) ;
  assign n1259 = ( x91 & x97 ) | ( x91 & x143 ) | ( x97 & x143 ) ;
  assign n1260 = n1258 | n1259 ;
  assign n1269 = n1260 & ~n1267 ;
  assign n1270 = ( ~n1260 & n1266 ) | ( ~n1260 & n1267 ) | ( n1266 & n1267 ) ;
  assign n1271 = ( ~n1268 & n1269 ) | ( ~n1268 & n1270 ) | ( n1269 & n1270 ) ;
  assign n1249 = ( ~x89 & x101 ) | ( ~x89 & x142 ) | ( x101 & x142 ) ;
  assign n1250 = ( x89 & x97 ) | ( x89 & x142 ) | ( x97 & x142 ) ;
  assign n1251 = n1249 | n1250 ;
  assign n1252 = ( ~x89 & x99 ) | ( ~x89 & x142 ) | ( x99 & x142 ) ;
  assign n1253 = ( x89 & x100 ) | ( x89 & x142 ) | ( x100 & x142 ) ;
  assign n1254 = n1252 & n1253 ;
  assign n1272 = n1251 & ~n1254 ;
  assign n1273 = ( ~n271 & n1271 ) | ( ~n271 & n1272 ) | ( n1271 & n1272 ) ;
  assign n1274 = ( n271 & ~n1272 ) | ( n271 & n1273 ) | ( ~n1272 & n1273 ) ;
  assign n1275 = ( ~n1271 & n1273 ) | ( ~n1271 & n1274 ) | ( n1273 & n1274 ) ;
  assign n1285 = ( ~x95 & x99 ) | ( ~x95 & x140 ) | ( x99 & x140 ) ;
  assign n1286 = ( x95 & x100 ) | ( x95 & x140 ) | ( x100 & x140 ) ;
  assign n1287 = n1285 & n1286 ;
  assign n1276 = ( x99 & ~x102 ) | ( x99 & x136 ) | ( ~x102 & x136 ) ;
  assign n1277 = ( x100 & x102 ) | ( x100 & x136 ) | ( x102 & x136 ) ;
  assign n1278 = n1276 & n1277 ;
  assign n1282 = ( x101 & ~x102 ) | ( x101 & x136 ) | ( ~x102 & x136 ) ;
  assign n1283 = ( x97 & x102 ) | ( x97 & x136 ) | ( x102 & x136 ) ;
  assign n1284 = n1282 | n1283 ;
  assign n1288 = ~n1278 & n1284 ;
  assign n1289 = n1287 & ~n1288 ;
  assign n1279 = ( ~x95 & x101 ) | ( ~x95 & x140 ) | ( x101 & x140 ) ;
  assign n1280 = ( x95 & x97 ) | ( x95 & x140 ) | ( x97 & x140 ) ;
  assign n1281 = n1279 | n1280 ;
  assign n1290 = n1281 & ~n1288 ;
  assign n1291 = ( ~n1281 & n1287 ) | ( ~n1281 & n1288 ) | ( n1287 & n1288 ) ;
  assign n1292 = ( ~n1289 & n1290 ) | ( ~n1289 & n1291 ) | ( n1290 & n1291 ) ;
  assign n1317 = ( n1275 & n1292 ) | ( n1275 & ~n1299 ) | ( n1292 & ~n1299 ) ;
  assign n1318 = ( n1275 & n1292 ) | ( n1275 & ~n1317 ) | ( n1292 & ~n1317 ) ;
  assign n1319 = ( n1299 & n1317 ) | ( n1299 & ~n1318 ) | ( n1317 & ~n1318 ) ;
  assign n1320 = n1316 & n1319 ;
  assign n1321 = n1316 | n1319 ;
  assign n1322 = ~n1320 & n1321 ;
  assign n1401 = ( x175 & ~x176 ) | ( x175 & n1322 ) | ( ~x176 & n1322 ) ;
  assign n1351 = ( ~n385 & n757 ) | ( ~n385 & n767 ) | ( n757 & n767 ) ;
  assign n1352 = ( n385 & ~n757 ) | ( n385 & n1351 ) | ( ~n757 & n1351 ) ;
  assign n1353 = ( ~n767 & n1351 ) | ( ~n767 & n1352 ) | ( n1351 & n1352 ) ;
  assign n1354 = ( n375 & n381 ) | ( n375 & n1353 ) | ( n381 & n1353 ) ;
  assign n1355 = ( n375 & n1353 ) | ( n375 & ~n1354 ) | ( n1353 & ~n1354 ) ;
  assign n1356 = ( n381 & ~n1354 ) | ( n381 & n1355 ) | ( ~n1354 & n1355 ) ;
  assign n1357 = n393 & ~n1356 ;
  assign n1358 = ~n393 & n1356 ;
  assign n1359 = n1357 | n1358 ;
  assign n1372 = n369 | n513 ;
  assign n1373 = ( x156 & n1359 ) | ( x156 & n1372 ) | ( n1359 & n1372 ) ;
  assign n1360 = ( n516 & n761 ) | ( n516 & n769 ) | ( n761 & n769 ) ;
  assign n1361 = ( n516 & n769 ) | ( n516 & ~n1360 ) | ( n769 & ~n1360 ) ;
  assign n1362 = ( n761 & ~n1360 ) | ( n761 & n1361 ) | ( ~n1360 & n1361 ) ;
  assign n1363 = ( n375 & n381 ) | ( n375 & ~n1362 ) | ( n381 & ~n1362 ) ;
  assign n1364 = ( ~n375 & n1362 ) | ( ~n375 & n1363 ) | ( n1362 & n1363 ) ;
  assign n1365 = ( ~n381 & n1363 ) | ( ~n381 & n1364 ) | ( n1363 & n1364 ) ;
  assign n1366 = n393 & n1365 ;
  assign n1367 = n393 | n1365 ;
  assign n1368 = ~n1366 & n1367 ;
  assign n1374 = ( ~x156 & n1368 ) | ( ~x156 & n1372 ) | ( n1368 & n1372 ) ;
  assign n1375 = n1373 & ~n1374 ;
  assign n1333 = n359 | n675 ;
  assign n1334 = ( n365 & n675 ) | ( n365 & n1333 ) | ( n675 & n1333 ) ;
  assign n1323 = n353 & n359 ;
  assign n1327 = n365 | n645 ;
  assign n1328 = ( n645 & n1323 ) | ( n645 & n1327 ) | ( n1323 & n1327 ) ;
  assign n1329 = n357 & n1328 ;
  assign n1330 = n357 & ~n650 ;
  assign n1331 = ( ~n357 & n650 ) | ( ~n357 & n1328 ) | ( n650 & n1328 ) ;
  assign n1332 = ( ~n1329 & n1330 ) | ( ~n1329 & n1331 ) | ( n1330 & n1331 ) ;
  assign n1335 = ~n1332 & n1334 ;
  assign n1336 = n1332 | n1334 ;
  assign n1337 = ( ~n1334 & n1335 ) | ( ~n1334 & n1336 ) | ( n1335 & n1336 ) ;
  assign n1324 = ( n347 & ~n365 ) | ( n347 & n1323 ) | ( ~n365 & n1323 ) ;
  assign n1325 = n347 & n645 ;
  assign n1326 = ( n365 & n1324 ) | ( n365 & n1325 ) | ( n1324 & n1325 ) ;
  assign n1338 = n651 | n1326 ;
  assign n1339 = ( ~n359 & n1337 ) | ( ~n359 & n1338 ) | ( n1337 & n1338 ) ;
  assign n1340 = ( n1337 & n1338 ) | ( n1337 & ~n1339 ) | ( n1338 & ~n1339 ) ;
  assign n1341 = ( n359 & n1339 ) | ( n359 & ~n1340 ) | ( n1339 & ~n1340 ) ;
  assign n1342 = ( n341 & n353 ) | ( n341 & ~n1341 ) | ( n353 & ~n1341 ) ;
  assign n1343 = ( ~n341 & n1341 ) | ( ~n341 & n1342 ) | ( n1341 & n1342 ) ;
  assign n1344 = ( ~n353 & n1342 ) | ( ~n353 & n1343 ) | ( n1342 & n1343 ) ;
  assign n1345 = n365 & n1344 ;
  assign n1346 = n365 | n1344 ;
  assign n1347 = ~n1345 & n1346 ;
  assign n1348 = ( x156 & ~n347 ) | ( x156 & n1347 ) | ( ~n347 & n1347 ) ;
  assign n1349 = n347 & n1348 ;
  assign n1350 = ( ~n1347 & n1348 ) | ( ~n1347 & n1349 ) | ( n1348 & n1349 ) ;
  assign n1376 = ( n645 & n651 ) | ( n645 & n653 ) | ( n651 & n653 ) ;
  assign n1377 = ~n645 & n650 ;
  assign n1378 = ( n501 & ~n645 ) | ( n501 & n1377 ) | ( ~n645 & n1377 ) ;
  assign n1379 = ( n501 & n645 ) | ( n501 & n1377 ) | ( n645 & n1377 ) ;
  assign n1380 = ( n645 & n1378 ) | ( n645 & ~n1379 ) | ( n1378 & ~n1379 ) ;
  assign n1381 = ( n675 & n1376 ) | ( n675 & ~n1380 ) | ( n1376 & ~n1380 ) ;
  assign n1382 = ( ~n1376 & n1380 ) | ( ~n1376 & n1381 ) | ( n1380 & n1381 ) ;
  assign n1383 = ( ~n675 & n1381 ) | ( ~n675 & n1382 ) | ( n1381 & n1382 ) ;
  assign n1384 = n359 & n1383 ;
  assign n1385 = n359 | n1383 ;
  assign n1386 = ~n1384 & n1385 ;
  assign n1387 = ( n341 & n353 ) | ( n341 & ~n1386 ) | ( n353 & ~n1386 ) ;
  assign n1388 = ( ~n341 & n1386 ) | ( ~n341 & n1387 ) | ( n1386 & n1387 ) ;
  assign n1389 = ( ~n353 & n1387 ) | ( ~n353 & n1388 ) | ( n1387 & n1388 ) ;
  assign n1390 = n365 & n1389 ;
  assign n1391 = n365 | n1389 ;
  assign n1392 = ~n1390 & n1391 ;
  assign n1393 = ( x156 & n347 ) | ( x156 & n1392 ) | ( n347 & n1392 ) ;
  assign n1394 = n347 & ~n1393 ;
  assign n1395 = ( n1392 & ~n1393 ) | ( n1392 & n1394 ) | ( ~n1393 & n1394 ) ;
  assign n1396 = n1350 | n1395 ;
  assign n1397 = n1375 & n1396 ;
  assign n1369 = ( x156 & n513 ) | ( x156 & n1368 ) | ( n513 & n1368 ) ;
  assign n1370 = ( ~x156 & n513 ) | ( ~x156 & n1359 ) | ( n513 & n1359 ) ;
  assign n1371 = ~n1369 & n1370 ;
  assign n1398 = ~n1371 & n1396 ;
  assign n1399 = ( n1371 & n1375 ) | ( n1371 & ~n1396 ) | ( n1375 & ~n1396 ) ;
  assign n1400 = ( ~n1397 & n1398 ) | ( ~n1397 & n1399 ) | ( n1398 & n1399 ) ;
  assign n1402 = ( x175 & x176 ) | ( x175 & ~n1400 ) | ( x176 & ~n1400 ) ;
  assign n1403 = n1401 & ~n1402 ;
  assign n1404 = ( ~x48 & x175 ) | ( ~x48 & n1403 ) | ( x175 & n1403 ) ;
  assign n1405 = x176 | n1403 ;
  assign n1406 = ( x48 & n1404 ) | ( x48 & n1405 ) | ( n1404 & n1405 ) ;
  assign n1416 = x36 & x176 ;
  assign n1413 = x175 & n1242 ;
  assign n1414 = x175 | n1173 ;
  assign n1415 = ( ~x175 & n1413 ) | ( ~x175 & n1414 ) | ( n1413 & n1414 ) ;
  assign n1417 = ~x176 & n1415 ;
  assign n1418 = ( x176 & ~n1416 ) | ( x176 & n1417 ) | ( ~n1416 & n1417 ) ;
  assign n1419 = ( x171 & ~x172 ) | ( x171 & n1418 ) | ( ~x172 & n1418 ) ;
  assign n1410 = x37 & x176 ;
  assign n1407 = x175 & n1400 ;
  assign n1408 = x175 | n1322 ;
  assign n1409 = ( ~x175 & n1407 ) | ( ~x175 & n1408 ) | ( n1407 & n1408 ) ;
  assign n1411 = ~x176 & n1409 ;
  assign n1412 = ( x176 & ~n1410 ) | ( x176 & n1411 ) | ( ~n1410 & n1411 ) ;
  assign n1420 = ( x171 & x172 ) | ( x171 & n1412 ) | ( x172 & n1412 ) ;
  assign n1421 = n1419 | n1420 ;
  assign n1422 = ( x22 & x171 ) | ( x22 & ~x172 ) | ( x171 & ~x172 ) ;
  assign n1423 = ( x3 & x171 ) | ( x3 & x172 ) | ( x171 & x172 ) ;
  assign n1424 = n1422 & n1423 ;
  assign n1425 = n1421 & ~n1424 ;
  assign n1426 = ( ~x173 & x174 ) | ( ~x173 & n1418 ) | ( x174 & n1418 ) ;
  assign n1427 = ( x173 & x174 ) | ( x173 & n1412 ) | ( x174 & n1412 ) ;
  assign n1428 = n1426 | n1427 ;
  assign n1429 = ( x22 & ~x173 ) | ( x22 & x174 ) | ( ~x173 & x174 ) ;
  assign n1430 = ( x3 & x173 ) | ( x3 & x174 ) | ( x173 & x174 ) ;
  assign n1431 = n1429 & n1430 ;
  assign n1432 = n1428 & ~n1431 ;
  assign n1436 = ( ~x157 & x158 ) | ( ~x157 & n1418 ) | ( x158 & n1418 ) ;
  assign n1437 = ( x157 & x158 ) | ( x157 & n1412 ) | ( x158 & n1412 ) ;
  assign n1438 = n1436 | n1437 ;
  assign n1433 = ( x78 & ~x157 ) | ( x78 & x158 ) | ( ~x157 & x158 ) ;
  assign n1434 = ( x77 & x157 ) | ( x77 & x158 ) | ( x157 & x158 ) ;
  assign n1435 = n1433 & n1434 ;
  assign n1439 = x63 & n1435 ;
  assign n1440 = ( x63 & ~n1438 ) | ( x63 & n1439 ) | ( ~n1438 & n1439 ) ;
  assign n1444 = ( ~x159 & x160 ) | ( ~x159 & n1418 ) | ( x160 & n1418 ) ;
  assign n1445 = ( x159 & x160 ) | ( x159 & n1412 ) | ( x160 & n1412 ) ;
  assign n1446 = n1444 | n1445 ;
  assign n1441 = ( x78 & ~x159 ) | ( x78 & x160 ) | ( ~x159 & x160 ) ;
  assign n1442 = ( x77 & x159 ) | ( x77 & x160 ) | ( x159 & x160 ) ;
  assign n1443 = n1441 & n1442 ;
  assign n1447 = x63 & n1443 ;
  assign n1448 = ( x63 & ~n1446 ) | ( x63 & n1447 ) | ( ~n1446 & n1447 ) ;
  assign y0 = x65 ;
  assign y1 = x112 ;
  assign y2 = x164 ;
  assign y3 = ~x150 ;
  assign y4 = ~x126 ;
  assign y5 = ~x130 ;
  assign y6 = n179 ;
  assign y7 = ~x151 ;
  assign y8 = ~x150 ;
  assign y9 = ~x150 ;
  assign y10 = ~x124 ;
  assign y11 = ~x128 ;
  assign y12 = n180 ;
  assign y13 = ~x98 ;
  assign y14 = ~x152 ;
  assign y15 = ~x155 ;
  assign y16 = ~x154 ;
  assign y17 = n181 ;
  assign y18 = n182 ;
  assign y19 = ~n183 ;
  assign y20 = ~n184 ;
  assign y21 = x63 ;
  assign y22 = x65 ;
  assign y23 = x0 ;
  assign y24 = x151 ;
  assign y25 = x113 ;
  assign y26 = ~x151 ;
  assign y27 = ~n186 ;
  assign y28 = ~n185 ;
  assign y29 = x0 ;
  assign y30 = x0 ;
  assign y31 = x0 ;
  assign y32 = x0 ;
  assign y33 = x113 ;
  assign y34 = ~x113 ;
  assign y35 = ~n189 ;
  assign y36 = ~n192 ;
  assign y37 = ~n192 ;
  assign y38 = ~n193 ;
  assign y39 = n197 ;
  assign y40 = n201 ;
  assign y41 = n205 ;
  assign y42 = n209 ;
  assign y43 = n264 ;
  assign y44 = n335 ;
  assign y45 = n397 ;
  assign y46 = n448 ;
  assign y47 = n453 ;
  assign y48 = n458 ;
  assign y49 = ~n476 ;
  assign y50 = n497 ;
  assign y51 = n525 ;
  assign y52 = n549 ;
  assign y53 = n525 ;
  assign y54 = n549 ;
  assign y55 = n558 ;
  assign y56 = n567 ;
  assign y57 = n576 ;
  assign y58 = n589 ;
  assign y59 = ~n596 ;
  assign y60 = n616 ;
  assign y61 = n627 ;
  assign y62 = n637 ;
  assign y63 = ~n644 ;
  assign y64 = n663 ;
  assign y65 = n674 ;
  assign y66 = n687 ;
  assign y67 = n697 ;
  assign y68 = ~n720 ;
  assign y69 = n743 ;
  assign y70 = ~n781 ;
  assign y71 = n803 ;
  assign y72 = n811 ;
  assign y73 = n819 ;
  assign y74 = ~n826 ;
  assign y75 = ~n833 ;
  assign y76 = ~n840 ;
  assign y77 = ~n847 ;
  assign y78 = ~n854 ;
  assign y79 = ~n861 ;
  assign y80 = ~n868 ;
  assign y81 = ~n875 ;
  assign y82 = n883 ;
  assign y83 = n891 ;
  assign y84 = n899 ;
  assign y85 = n907 ;
  assign y86 = n915 ;
  assign y87 = n923 ;
  assign y88 = n931 ;
  assign y89 = n939 ;
  assign y90 = n951 ;
  assign y91 = n954 ;
  assign y92 = ~n960 ;
  assign y93 = n966 ;
  assign y94 = ~n972 ;
  assign y95 = ~n978 ;
  assign y96 = n987 ;
  assign y97 = ~n993 ;
  assign y98 = n999 ;
  assign y99 = n1005 ;
  assign y100 = n1011 ;
  assign y101 = n1018 ;
  assign y102 = n1025 ;
  assign y103 = ~n1032 ;
  assign y104 = n1039 ;
  assign y105 = n1046 ;
  assign y106 = ~n1053 ;
  assign y107 = n1060 ;
  assign y108 = n1067 ;
  assign y109 = n1075 ;
  assign y110 = n1083 ;
  assign y111 = n1091 ;
  assign y112 = n1099 ;
  assign y113 = n1107 ;
  assign y114 = n1115 ;
  assign y115 = n1123 ;
  assign y116 = n1131 ;
  assign y117 = n1248 ;
  assign y118 = n1406 ;
  assign y119 = ~n1425 ;
  assign y120 = ~n1432 ;
  assign y121 = ~n1440 ;
  assign y122 = ~n1448 ;
endmodule
