module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , x128 , x129 , x130 , x131 , x132 , x133 , x134 , x135 , x136 , x137 , x138 , x139 , x140 , x141 , x142 , x143 , x144 , x145 , x146 , x147 , x148 , x149 , x150 , x151 , x152 , x153 , x154 , x155 , x156 , x157 , x158 , x159 , x160 , x161 , x162 , x163 , x164 , x165 , x166 , x167 , x168 , x169 , x170 , x171 , x172 , x173 , x174 , x175 , x176 , x177 , x178 , x179 , x180 , x181 , x182 , x183 , x184 , x185 , x186 , x187 , x188 , x189 , x190 , x191 , x192 , x193 , x194 , x195 , x196 , x197 , x198 , x199 , x200 , x201 , x202 , x203 , x204 , x205 , x206 , x207 , x208 , x209 , x210 , x211 , x212 , x213 , x214 , x215 , x216 , x217 , x218 , x219 , x220 , x221 , x222 , x223 , x224 , x225 , x226 , x227 , x228 , x229 , x230 , x231 , x232 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 ;
  wire n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 ;
  assign n234 = x215 & x217 ;
  assign n235 = ( ~x214 & x216 ) | ( ~x214 & n234 ) | ( x216 & n234 ) ;
  assign n236 = x214 & n235 ;
  assign n237 = x1 & x196 ;
  assign n238 = x10 & n237 ;
  assign n239 = x73 & x190 ;
  assign n240 = x6 & x196 ;
  assign n241 = x194 & n240 ;
  assign n242 = x222 & n240 ;
  assign n243 = x52 & x95 ;
  assign n244 = ( ~x42 & x85 ) | ( ~x42 & n243 ) | ( x85 & n243 ) ;
  assign n245 = x42 & n244 ;
  assign n246 = x63 & x105 ;
  assign n247 = ( ~x31 & x75 ) | ( ~x31 & n246 ) | ( x75 & n246 ) ;
  assign n248 = x31 & n247 ;
  assign n249 = n245 & n248 ;
  assign n250 = x194 & ~n245 ;
  assign n251 = x222 | n250 ;
  assign n252 = ( ~n248 & n250 ) | ( ~n248 & n251 ) | ( n250 & n251 ) ;
  assign n253 = ( x108 & x220 ) | ( x108 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n254 = ( ~x78 & x220 ) | ( ~x78 & x221 ) | ( x220 & x221 ) ;
  assign n255 = n253 & ~n254 ;
  assign n256 = ( x88 & ~x220 ) | ( x88 & x221 ) | ( ~x220 & x221 ) ;
  assign n257 = ( x98 & x220 ) | ( x98 & x221 ) | ( x220 & x221 ) ;
  assign n258 = n256 & n257 ;
  assign n259 = n255 | n258 ;
  assign n260 = ( x107 & x220 ) | ( x107 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n261 = ( ~x77 & x220 ) | ( ~x77 & x221 ) | ( x220 & x221 ) ;
  assign n262 = n260 & ~n261 ;
  assign n263 = ( x87 & ~x220 ) | ( x87 & x221 ) | ( ~x220 & x221 ) ;
  assign n264 = ( x97 & x220 ) | ( x97 & x221 ) | ( x220 & x221 ) ;
  assign n265 = n263 & n264 ;
  assign n266 = n262 | n265 ;
  assign n267 = ( x109 & x220 ) | ( x109 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n268 = ( ~x79 & x220 ) | ( ~x79 & x221 ) | ( x220 & x221 ) ;
  assign n269 = n267 & ~n268 ;
  assign n270 = ( x89 & ~x220 ) | ( x89 & x221 ) | ( ~x220 & x221 ) ;
  assign n271 = ( x99 & x220 ) | ( x99 & x221 ) | ( x220 & x221 ) ;
  assign n272 = n270 & n271 ;
  assign n273 = n269 | n272 ;
  assign n274 = ( x67 & x192 ) | ( x67 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n275 = ( ~x35 & x192 ) | ( ~x35 & x195 ) | ( x192 & x195 ) ;
  assign n276 = n274 & ~n275 ;
  assign n277 = ( x56 & ~x192 ) | ( x56 & x195 ) | ( ~x192 & x195 ) ;
  assign n278 = ( x45 & x192 ) | ( x45 & x195 ) | ( x192 & x195 ) ;
  assign n279 = n277 & n278 ;
  assign n280 = n276 | n279 ;
  assign n281 = ( x68 & x192 ) | ( x68 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n282 = ( ~x36 & x192 ) | ( ~x36 & x195 ) | ( x192 & x195 ) ;
  assign n283 = n281 & ~n282 ;
  assign n284 = ( x57 & ~x192 ) | ( x57 & x195 ) | ( ~x192 & x195 ) ;
  assign n285 = ( x46 & x192 ) | ( x46 & x195 ) | ( x192 & x195 ) ;
  assign n286 = n284 & n285 ;
  assign n287 = n283 | n286 ;
  assign n288 = ( x69 & x192 ) | ( x69 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n289 = ( ~x37 & x192 ) | ( ~x37 & x195 ) | ( x192 & x195 ) ;
  assign n290 = n288 & ~n289 ;
  assign n291 = ( x58 & ~x192 ) | ( x58 & x195 ) | ( ~x192 & x195 ) ;
  assign n292 = ( x47 & x192 ) | ( x47 & x195 ) | ( x192 & x195 ) ;
  assign n293 = n291 & n292 ;
  assign n294 = n290 | n293 ;
  assign n295 = ( x62 & x192 ) | ( x62 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n296 = ( ~x30 & x192 ) | ( ~x30 & x195 ) | ( x192 & x195 ) ;
  assign n297 = n295 & ~n296 ;
  assign n298 = ( x51 & ~x192 ) | ( x51 & x195 ) | ( ~x192 & x195 ) ;
  assign n299 = ( x41 & x192 ) | ( x41 & x195 ) | ( x192 & x195 ) ;
  assign n300 = n298 & n299 ;
  assign n301 = n297 | n300 ;
  assign n302 = x197 & ~n301 ;
  assign n303 = x27 & x196 ;
  assign n304 = ( x191 & n252 ) | ( x191 & n303 ) | ( n252 & n303 ) ;
  assign n305 = ~n252 & n304 ;
  assign n306 = x196 & ~n252 ;
  assign n307 = x191 & n306 ;
  assign n308 = ~x0 & n307 ;
  assign n309 = ( ~x2 & n307 ) | ( ~x2 & n308 ) | ( n307 & n308 ) ;
  assign n310 = ( x70 & x192 ) | ( x70 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n311 = ( ~x38 & x192 ) | ( ~x38 & x195 ) | ( x192 & x195 ) ;
  assign n312 = n310 & ~n311 ;
  assign n313 = ( x59 & ~x192 ) | ( x59 & x195 ) | ( ~x192 & x195 ) ;
  assign n314 = ( x48 & x192 ) | ( x48 & x195 ) | ( x192 & x195 ) ;
  assign n315 = n313 & n314 ;
  assign n316 = n312 | n315 ;
  assign n317 = ( x66 & x192 ) | ( x66 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n318 = ( ~x34 & x192 ) | ( ~x34 & x195 ) | ( x192 & x195 ) ;
  assign n319 = n317 & ~n318 ;
  assign n320 = ( x55 & x192 ) | ( x55 & ~n319 ) | ( x192 & ~n319 ) ;
  assign n321 = x195 | n319 ;
  assign n322 = ( x55 & ~n320 ) | ( x55 & n321 ) | ( ~n320 & n321 ) ;
  assign n323 = ( x65 & x192 ) | ( x65 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n324 = ( ~x33 & x192 ) | ( ~x33 & x195 ) | ( x192 & x195 ) ;
  assign n325 = n323 & ~n324 ;
  assign n326 = ( x54 & ~x192 ) | ( x54 & x195 ) | ( ~x192 & x195 ) ;
  assign n327 = ( x44 & x192 ) | ( x44 & x195 ) | ( x192 & x195 ) ;
  assign n328 = n326 & n327 ;
  assign n329 = n325 | n328 ;
  assign n330 = ( x64 & x192 ) | ( x64 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n331 = ( ~x32 & x192 ) | ( ~x32 & x195 ) | ( x192 & x195 ) ;
  assign n332 = n330 & ~n331 ;
  assign n333 = ( x53 & ~x192 ) | ( x53 & x195 ) | ( ~x192 & x195 ) ;
  assign n334 = ( x43 & x192 ) | ( x43 & x195 ) | ( x192 & x195 ) ;
  assign n335 = n333 & n334 ;
  assign n336 = n332 | n335 ;
  assign n337 = x198 & n294 ;
  assign n338 = ( x71 & x192 ) | ( x71 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n339 = ( ~x39 & x192 ) | ( ~x39 & x195 ) | ( x192 & x195 ) ;
  assign n340 = n338 & ~n339 ;
  assign n341 = ( x60 & ~x192 ) | ( x60 & x195 ) | ( ~x192 & x195 ) ;
  assign n342 = ( x49 & x192 ) | ( x49 & x195 ) | ( x192 & x195 ) ;
  assign n343 = n341 & n342 ;
  assign n344 = n340 | n343 ;
  assign n345 = x198 | n344 ;
  assign n346 = ( ~x198 & n337 ) | ( ~x198 & n345 ) | ( n337 & n345 ) ;
  assign n347 = x198 & n287 ;
  assign n348 = x198 | n316 ;
  assign n349 = ( ~x198 & n347 ) | ( ~x198 & n348 ) | ( n347 & n348 ) ;
  assign n350 = x197 & ~n344 ;
  assign n351 = ( x193 & n344 ) | ( x193 & ~n350 ) | ( n344 & ~n350 ) ;
  assign n352 = x193 | n344 ;
  assign n353 = x198 & n352 ;
  assign n354 = x198 | n301 ;
  assign n355 = ( ~x198 & n353 ) | ( ~x198 & n354 ) | ( n353 & n354 ) ;
  assign n356 = ( x106 & x220 ) | ( x106 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n357 = ( ~x76 & x220 ) | ( ~x76 & x221 ) | ( x220 & x221 ) ;
  assign n358 = n356 & ~n357 ;
  assign n359 = ( x86 & ~x220 ) | ( x86 & x221 ) | ( ~x220 & x221 ) ;
  assign n360 = ( x96 & x220 ) | ( x96 & x221 ) | ( x220 & x221 ) ;
  assign n361 = n359 & n360 ;
  assign n362 = n358 | n361 ;
  assign n363 = ( x218 & ~x219 ) | ( x218 & n362 ) | ( ~x219 & n362 ) ;
  assign n364 = ~x218 & n363 ;
  assign n365 = ( ~n362 & n363 ) | ( ~n362 & n364 ) | ( n363 & n364 ) ;
  assign n366 = x225 & ~x226 ;
  assign n367 = x225 | x226 ;
  assign n368 = ( ~x225 & n366 ) | ( ~x225 & n367 ) | ( n366 & n367 ) ;
  assign n369 = x223 & ~x224 ;
  assign n370 = x223 | x224 ;
  assign n371 = ( ~x223 & n369 ) | ( ~x223 & n370 ) | ( n369 & n370 ) ;
  assign n372 = ( x200 & x201 ) | ( x200 & x229 ) | ( x201 & x229 ) ;
  assign n373 = ( x200 & x201 ) | ( x200 & ~n372 ) | ( x201 & ~n372 ) ;
  assign n374 = ( x229 & ~n372 ) | ( x229 & n373 ) | ( ~n372 & n373 ) ;
  assign n375 = ~x230 & n374 ;
  assign n376 = x230 & ~n374 ;
  assign n377 = n375 | n376 ;
  assign n378 = x227 & ~x228 ;
  assign n379 = x227 | x228 ;
  assign n380 = ( ~x227 & n378 ) | ( ~x227 & n379 ) | ( n378 & n379 ) ;
  assign n381 = ( n371 & n377 ) | ( n371 & n380 ) | ( n377 & n380 ) ;
  assign n382 = ( n377 & n380 ) | ( n377 & ~n381 ) | ( n380 & ~n381 ) ;
  assign n383 = ( n371 & ~n381 ) | ( n371 & n382 ) | ( ~n381 & n382 ) ;
  assign n384 = n368 & ~n383 ;
  assign n385 = ~n368 & n383 ;
  assign n386 = n384 | n385 ;
  assign n387 = x9 & ~n386 ;
  assign n388 = x213 & ~x232 ;
  assign n389 = x213 | x232 ;
  assign n390 = ( ~x213 & n388 ) | ( ~x213 & n389 ) | ( n388 & n389 ) ;
  assign n391 = x214 & ~x215 ;
  assign n392 = x214 | x215 ;
  assign n393 = ( ~x214 & n391 ) | ( ~x214 & n392 ) | ( n391 & n392 ) ;
  assign n394 = ( ~x216 & n390 ) | ( ~x216 & n393 ) | ( n390 & n393 ) ;
  assign n395 = ( n390 & n393 ) | ( n390 & ~n394 ) | ( n393 & ~n394 ) ;
  assign n396 = ( x216 & n394 ) | ( x216 & ~n395 ) | ( n394 & ~n395 ) ;
  assign n397 = ~x217 & n396 ;
  assign n398 = x217 & ~n396 ;
  assign n399 = n397 | n398 ;
  assign n400 = ( x218 & ~x219 ) | ( x218 & n399 ) | ( ~x219 & n399 ) ;
  assign n401 = ( x218 & n399 ) | ( x218 & ~n400 ) | ( n399 & ~n400 ) ;
  assign n402 = ( x219 & n400 ) | ( x219 & ~n401 ) | ( n400 & ~n401 ) ;
  assign n403 = x203 & ~x231 ;
  assign n404 = x203 | x231 ;
  assign n405 = ( ~x203 & n403 ) | ( ~x203 & n404 ) | ( n403 & n404 ) ;
  assign n406 = x204 & ~x205 ;
  assign n407 = x204 | x205 ;
  assign n408 = ( ~x204 & n406 ) | ( ~x204 & n407 ) | ( n406 & n407 ) ;
  assign n409 = ( ~x206 & n405 ) | ( ~x206 & n408 ) | ( n405 & n408 ) ;
  assign n410 = ( n405 & n408 ) | ( n405 & ~n409 ) | ( n408 & ~n409 ) ;
  assign n411 = ( x206 & n409 ) | ( x206 & ~n410 ) | ( n409 & ~n410 ) ;
  assign n412 = ~x207 & n411 ;
  assign n413 = x207 & ~n411 ;
  assign n414 = n412 | n413 ;
  assign n415 = ( x208 & x209 ) | ( x208 & x210 ) | ( x209 & x210 ) ;
  assign n416 = ( x208 & x209 ) | ( x208 & ~n415 ) | ( x209 & ~n415 ) ;
  assign n417 = ( x210 & ~n415 ) | ( x210 & n416 ) | ( ~n415 & n416 ) ;
  assign n418 = ~x211 & n417 ;
  assign n419 = x211 & ~n417 ;
  assign n420 = n418 | n419 ;
  assign n421 = ~n414 & n420 ;
  assign n422 = n414 & n420 ;
  assign n423 = ( n414 & n421 ) | ( n414 & ~n422 ) | ( n421 & ~n422 ) ;
  assign n424 = ( x111 & x220 ) | ( x111 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n425 = ( ~x81 & x220 ) | ( ~x81 & x221 ) | ( x220 & x221 ) ;
  assign n426 = n424 & ~n425 ;
  assign n427 = ( x91 & ~x220 ) | ( x91 & x221 ) | ( ~x220 & x221 ) ;
  assign n428 = ( x101 & x220 ) | ( x101 & x221 ) | ( x220 & x221 ) ;
  assign n429 = n427 & n428 ;
  assign n430 = n426 | n429 ;
  assign n431 = x22 & ~n430 ;
  assign n432 = x19 | x22 ;
  assign n433 = ( x213 & n431 ) | ( x213 & ~n432 ) | ( n431 & ~n432 ) ;
  assign n434 = ( ~x213 & n432 ) | ( ~x213 & n433 ) | ( n432 & n433 ) ;
  assign n435 = ( ~n431 & n433 ) | ( ~n431 & n434 ) | ( n433 & n434 ) ;
  assign n436 = x22 & ~n259 ;
  assign n437 = x22 | x25 ;
  assign n438 = ( x216 & n436 ) | ( x216 & ~n437 ) | ( n436 & ~n437 ) ;
  assign n439 = ( ~x216 & n437 ) | ( ~x216 & n438 ) | ( n437 & n438 ) ;
  assign n440 = ( ~n436 & n438 ) | ( ~n436 & n439 ) | ( n438 & n439 ) ;
  assign n441 = ( x110 & x220 ) | ( x110 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n442 = ( ~x80 & x220 ) | ( ~x80 & x221 ) | ( x220 & x221 ) ;
  assign n443 = n441 & ~n442 ;
  assign n444 = ( x90 & ~x220 ) | ( x90 & x221 ) | ( ~x220 & x221 ) ;
  assign n445 = ( x100 & x220 ) | ( x100 & x221 ) | ( x220 & x221 ) ;
  assign n446 = n444 & n445 ;
  assign n447 = n443 | n446 ;
  assign n448 = x22 & ~n447 ;
  assign n449 = x22 | x24 ;
  assign n450 = ( x214 & n448 ) | ( x214 & ~n449 ) | ( n448 & ~n449 ) ;
  assign n451 = ( ~x214 & n449 ) | ( ~x214 & n450 ) | ( n449 & n450 ) ;
  assign n452 = ( ~n448 & n450 ) | ( ~n448 & n451 ) | ( n450 & n451 ) ;
  assign n453 = x22 & ~n273 ;
  assign n454 = x20 | x22 ;
  assign n455 = ( x215 & n453 ) | ( x215 & ~n454 ) | ( n453 & ~n454 ) ;
  assign n456 = ( ~x215 & n454 ) | ( ~x215 & n455 ) | ( n454 & n455 ) ;
  assign n457 = ( ~n453 & n455 ) | ( ~n453 & n456 ) | ( n455 & n456 ) ;
  assign n458 = n452 & n457 ;
  assign n459 = ( ~n435 & n440 ) | ( ~n435 & n458 ) | ( n440 & n458 ) ;
  assign n460 = n435 & n459 ;
  assign n461 = x22 & ~n266 ;
  assign n462 = x22 | x26 ;
  assign n463 = ( x217 & n461 ) | ( x217 & ~n462 ) | ( n461 & ~n462 ) ;
  assign n464 = ( ~x217 & n462 ) | ( ~x217 & n463 ) | ( n462 & n463 ) ;
  assign n465 = ( ~n461 & n463 ) | ( ~n461 & n464 ) | ( n463 & n464 ) ;
  assign n466 = ( ~x22 & n362 ) | ( ~x22 & n465 ) | ( n362 & n465 ) ;
  assign n467 = ( x21 & x22 ) | ( x21 & n465 ) | ( x22 & n465 ) ;
  assign n468 = n466 & n467 ;
  assign n469 = ( x112 & x220 ) | ( x112 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n470 = ( ~x82 & x220 ) | ( ~x82 & x221 ) | ( x220 & x221 ) ;
  assign n471 = n469 & ~n470 ;
  assign n472 = ( x92 & ~x220 ) | ( x92 & x221 ) | ( ~x220 & x221 ) ;
  assign n473 = ( x102 & x220 ) | ( x102 & x221 ) | ( x220 & x221 ) ;
  assign n474 = n472 & n473 ;
  assign n475 = n471 | n474 ;
  assign n476 = x22 & ~n475 ;
  assign n477 = x22 | x23 ;
  assign n478 = ( x211 & n476 ) | ( x211 & ~n477 ) | ( n476 & ~n477 ) ;
  assign n479 = ( ~x211 & n477 ) | ( ~x211 & n478 ) | ( n477 & n478 ) ;
  assign n480 = ( ~n476 & n478 ) | ( ~n476 & n479 ) | ( n478 & n479 ) ;
  assign n481 = n468 & n480 ;
  assign n482 = n460 & n481 ;
  assign n483 = x11 & ~n322 ;
  assign n484 = x11 | x16 ;
  assign n485 = ( x207 & n483 ) | ( x207 & ~n484 ) | ( n483 & ~n484 ) ;
  assign n486 = ( ~x207 & n484 ) | ( ~x207 & n485 ) | ( n484 & n485 ) ;
  assign n487 = ( ~n483 & n485 ) | ( ~n483 & n486 ) | ( n485 & n486 ) ;
  assign n488 = ( x104 & x220 ) | ( x104 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n489 = ( ~x74 & x220 ) | ( ~x74 & x221 ) | ( x220 & x221 ) ;
  assign n490 = n488 & ~n489 ;
  assign n491 = ( x84 & ~x220 ) | ( x84 & x221 ) | ( ~x220 & x221 ) ;
  assign n492 = ( x94 & x220 ) | ( x94 & x221 ) | ( x220 & x221 ) ;
  assign n493 = n491 & n492 ;
  assign n494 = n490 | n493 ;
  assign n495 = x22 & ~n494 ;
  assign n496 = x18 | x22 ;
  assign n497 = ( x210 & n495 ) | ( x210 & ~n496 ) | ( n495 & ~n496 ) ;
  assign n498 = ( ~x210 & n496 ) | ( ~x210 & n497 ) | ( n496 & n497 ) ;
  assign n499 = ( ~n495 & n497 ) | ( ~n495 & n498 ) | ( n497 & n498 ) ;
  assign n500 = x11 & ~n329 ;
  assign n501 = x5 | x11 ;
  assign n502 = ( x208 & n500 ) | ( x208 & ~n501 ) | ( n500 & ~n501 ) ;
  assign n503 = ( ~x208 & n501 ) | ( ~x208 & n502 ) | ( n501 & n502 ) ;
  assign n504 = ( ~n500 & n502 ) | ( ~n500 & n503 ) | ( n502 & n503 ) ;
  assign n505 = x11 & ~n336 ;
  assign n506 = x11 | x17 ;
  assign n507 = ( x209 & n505 ) | ( x209 & ~n506 ) | ( n505 & ~n506 ) ;
  assign n508 = ( ~x209 & n506 ) | ( ~x209 & n507 ) | ( n506 & n507 ) ;
  assign n509 = ( ~n505 & n507 ) | ( ~n505 & n508 ) | ( n507 & n508 ) ;
  assign n510 = n504 & n509 ;
  assign n511 = ( ~n487 & n499 ) | ( ~n487 & n510 ) | ( n499 & n510 ) ;
  assign n512 = n487 & n511 ;
  assign n513 = x11 & ~n280 ;
  assign n514 = x11 | x15 ;
  assign n515 = ( x206 & n513 ) | ( x206 & ~n514 ) | ( n513 & ~n514 ) ;
  assign n516 = ( ~x206 & n514 ) | ( ~x206 & n515 ) | ( n514 & n515 ) ;
  assign n517 = ( ~n513 & n515 ) | ( ~n513 & n516 ) | ( n515 & n516 ) ;
  assign n518 = x11 & ~n344 ;
  assign n519 = x3 | x11 ;
  assign n520 = ( x201 & n518 ) | ( x201 & ~n519 ) | ( n518 & ~n519 ) ;
  assign n521 = ( ~x201 & n519 ) | ( ~x201 & n520 ) | ( n519 & n520 ) ;
  assign n522 = ( ~n518 & n520 ) | ( ~n518 & n521 ) | ( n520 & n521 ) ;
  assign n523 = x11 & ~n287 ;
  assign n524 = x11 | x14 ;
  assign n525 = ( x205 & n523 ) | ( x205 & ~n524 ) | ( n523 & ~n524 ) ;
  assign n526 = ( ~x205 & n524 ) | ( ~x205 & n525 ) | ( n524 & n525 ) ;
  assign n527 = ( ~n523 & n525 ) | ( ~n523 & n526 ) | ( n525 & n526 ) ;
  assign n528 = x11 & ~n316 ;
  assign n529 = x11 | x13 ;
  assign n530 = ( x203 & n528 ) | ( x203 & ~n529 ) | ( n528 & ~n529 ) ;
  assign n531 = ( ~x203 & n529 ) | ( ~x203 & n530 ) | ( n529 & n530 ) ;
  assign n532 = ( ~n528 & n530 ) | ( ~n528 & n531 ) | ( n530 & n531 ) ;
  assign n533 = x11 & ~n294 ;
  assign n534 = x4 | x11 ;
  assign n535 = ( x204 & n533 ) | ( x204 & ~n534 ) | ( n533 & ~n534 ) ;
  assign n536 = ( ~x204 & n534 ) | ( ~x204 & n535 ) | ( n534 & n535 ) ;
  assign n537 = ( ~n533 & n535 ) | ( ~n533 & n536 ) | ( n535 & n536 ) ;
  assign n538 = n532 & n537 ;
  assign n539 = ( ~n522 & n527 ) | ( ~n522 & n538 ) | ( n527 & n538 ) ;
  assign n540 = n522 & n539 ;
  assign n541 = x11 & ~n301 ;
  assign n542 = x11 | x12 ;
  assign n543 = ( x200 & n541 ) | ( x200 & ~n542 ) | ( n541 & ~n542 ) ;
  assign n544 = ( ~x200 & n542 ) | ( ~x200 & n543 ) | ( n542 & n543 ) ;
  assign n545 = ( ~n541 & n543 ) | ( ~n541 & n544 ) | ( n543 & n544 ) ;
  assign n546 = n540 & n545 ;
  assign n547 = ( ~n512 & n517 ) | ( ~n512 & n546 ) | ( n517 & n546 ) ;
  assign n548 = n512 & n547 ;
  assign n549 = n482 & n548 ;
  assign n550 = x8 & n549 ;
  assign n551 = ( n301 & n344 ) | ( n301 & n352 ) | ( n344 & n352 ) ;
  assign n552 = ( n301 & ~n344 ) | ( n301 & n352 ) | ( ~n344 & n352 ) ;
  assign n553 = ( n344 & ~n551 ) | ( n344 & n552 ) | ( ~n551 & n552 ) ;
  assign n554 = ( x72 & x192 ) | ( x72 & ~x195 ) | ( x192 & ~x195 ) ;
  assign n555 = ( ~x40 & x192 ) | ( ~x40 & x195 ) | ( x192 & x195 ) ;
  assign n556 = n554 & ~n555 ;
  assign n557 = ( x61 & ~x192 ) | ( x61 & x195 ) | ( ~x192 & x195 ) ;
  assign n558 = ( x50 & x192 ) | ( x50 & x195 ) | ( x192 & x195 ) ;
  assign n559 = n557 & n558 ;
  assign n560 = n556 | n559 ;
  assign n561 = x197 & ~n553 ;
  assign n562 = ( n553 & n560 ) | ( n553 & ~n561 ) | ( n560 & ~n561 ) ;
  assign n563 = ( n553 & ~n560 ) | ( n553 & n561 ) | ( ~n560 & n561 ) ;
  assign n564 = ( ~n553 & n562 ) | ( ~n553 & n563 ) | ( n562 & n563 ) ;
  assign n565 = n430 & ~n475 ;
  assign n566 = n430 & n475 ;
  assign n567 = ( n475 & n565 ) | ( n475 & ~n566 ) | ( n565 & ~n566 ) ;
  assign n568 = ( x113 & x220 ) | ( x113 & ~x221 ) | ( x220 & ~x221 ) ;
  assign n569 = ( ~x83 & x220 ) | ( ~x83 & x221 ) | ( x220 & x221 ) ;
  assign n570 = n568 & ~n569 ;
  assign n571 = ( x93 & ~x220 ) | ( x93 & x221 ) | ( ~x220 & x221 ) ;
  assign n572 = ( x103 & x220 ) | ( x103 & x221 ) | ( x220 & x221 ) ;
  assign n573 = n571 & n572 ;
  assign n574 = ~n570 & n573 ;
  assign n575 = ( n494 & n570 ) | ( n494 & ~n574 ) | ( n570 & ~n574 ) ;
  assign n576 = ( ~n494 & n570 ) | ( ~n494 & n574 ) | ( n570 & n574 ) ;
  assign n577 = ( ~n570 & n575 ) | ( ~n570 & n576 ) | ( n575 & n576 ) ;
  assign n578 = ( n259 & ~n266 ) | ( n259 & n362 ) | ( ~n266 & n362 ) ;
  assign n579 = ( n259 & n362 ) | ( n259 & ~n578 ) | ( n362 & ~n578 ) ;
  assign n580 = ( n266 & n578 ) | ( n266 & ~n579 ) | ( n578 & ~n579 ) ;
  assign n581 = ~n273 & n447 ;
  assign n582 = n273 & n447 ;
  assign n583 = ( n273 & n581 ) | ( n273 & ~n582 ) | ( n581 & ~n582 ) ;
  assign n584 = ( n577 & ~n580 ) | ( n577 & n583 ) | ( ~n580 & n583 ) ;
  assign n585 = ( n580 & ~n583 ) | ( n580 & n584 ) | ( ~n583 & n584 ) ;
  assign n586 = ( ~n577 & n584 ) | ( ~n577 & n585 ) | ( n584 & n585 ) ;
  assign n587 = n567 & n586 ;
  assign n588 = n567 | n586 ;
  assign n589 = ~n587 & n588 ;
  assign n590 = ~x28 & n589 ;
  assign n591 = ~n301 & n560 ;
  assign n592 = n301 & n560 ;
  assign n593 = ( n301 & n591 ) | ( n301 & ~n592 ) | ( n591 & ~n592 ) ;
  assign n594 = n316 & n344 ;
  assign n595 = ~n316 & n344 ;
  assign n596 = ( n316 & ~n594 ) | ( n316 & n595 ) | ( ~n594 & n595 ) ;
  assign n597 = ( ~n280 & n322 ) | ( ~n280 & n329 ) | ( n322 & n329 ) ;
  assign n598 = ( n280 & ~n322 ) | ( n280 & n597 ) | ( ~n322 & n597 ) ;
  assign n599 = ( ~n329 & n597 ) | ( ~n329 & n598 ) | ( n597 & n598 ) ;
  assign n600 = n336 | n599 ;
  assign n601 = n336 & n599 ;
  assign n602 = n600 & ~n601 ;
  assign n603 = ( n352 & n596 ) | ( n352 & n602 ) | ( n596 & n602 ) ;
  assign n604 = ( n352 & n602 ) | ( n352 & ~n603 ) | ( n602 & ~n603 ) ;
  assign n605 = ( n596 & ~n603 ) | ( n596 & n604 ) | ( ~n603 & n604 ) ;
  assign n606 = n593 & ~n605 ;
  assign n607 = ~n593 & n605 ;
  assign n608 = n606 | n607 ;
  assign n609 = x198 & n608 ;
  assign n610 = x198 | n560 ;
  assign n611 = ( ~x198 & n609 ) | ( ~x198 & n610 ) | ( n609 & n610 ) ;
  assign n612 = ( n287 & n593 ) | ( n287 & n596 ) | ( n593 & n596 ) ;
  assign n613 = ( n593 & n596 ) | ( n593 & ~n612 ) | ( n596 & ~n612 ) ;
  assign n614 = ( n287 & ~n612 ) | ( n287 & n613 ) | ( ~n612 & n613 ) ;
  assign n615 = n294 & ~n614 ;
  assign n616 = ~n294 & n614 ;
  assign n617 = n615 | n616 ;
  assign n618 = ( x28 & n602 ) | ( x28 & ~n617 ) | ( n602 & ~n617 ) ;
  assign n619 = n602 & ~n618 ;
  assign n620 = ( n617 & n618 ) | ( n617 & ~n619 ) | ( n618 & ~n619 ) ;
  assign n621 = x202 | n259 ;
  assign n622 = ( ~x29 & n273 ) | ( ~x29 & n621 ) | ( n273 & n621 ) ;
  assign n623 = n273 & ~n622 ;
  assign n624 = ~x214 & n623 ;
  assign n625 = x203 & ~n623 ;
  assign n626 = ( n623 & ~n624 ) | ( n623 & n625 ) | ( ~n624 & n625 ) ;
  assign n627 = ~x213 & n623 ;
  assign n628 = x201 & ~n623 ;
  assign n629 = ( n623 & ~n627 ) | ( n623 & n628 ) | ( ~n627 & n628 ) ;
  assign n630 = n344 | n629 ;
  assign n631 = ( n316 & n626 ) | ( n316 & ~n630 ) | ( n626 & ~n630 ) ;
  assign n632 = n344 & n629 ;
  assign n633 = ( n316 & n626 ) | ( n316 & ~n632 ) | ( n626 & ~n632 ) ;
  assign n634 = ~n631 & n633 ;
  assign n635 = ( x211 & n301 ) | ( x211 & n623 ) | ( n301 & n623 ) ;
  assign n636 = ( x200 & n301 ) | ( x200 & ~n623 ) | ( n301 & ~n623 ) ;
  assign n637 = n635 | n636 ;
  assign n638 = ( ~x7 & x216 ) | ( ~x7 & n623 ) | ( x216 & n623 ) ;
  assign n639 = ( x7 & ~x205 ) | ( x7 & n623 ) | ( ~x205 & n623 ) ;
  assign n640 = ~n638 & n639 ;
  assign n641 = x7 & n287 ;
  assign n642 = ( ~x7 & x217 ) | ( ~x7 & n623 ) | ( x217 & n623 ) ;
  assign n643 = ( x7 & ~x206 ) | ( x7 & n623 ) | ( ~x206 & n623 ) ;
  assign n644 = ~n642 & n643 ;
  assign n645 = x7 & n280 ;
  assign n646 = n644 & ~n645 ;
  assign n647 = n644 | n645 ;
  assign n648 = ( ~n644 & n646 ) | ( ~n644 & n647 ) | ( n646 & n647 ) ;
  assign n649 = ~x215 & n623 ;
  assign n650 = x204 & ~n623 ;
  assign n651 = ( n623 & ~n649 ) | ( n623 & n650 ) | ( ~n649 & n650 ) ;
  assign n652 = ( n294 & n648 ) | ( n294 & n651 ) | ( n648 & n651 ) ;
  assign n653 = ( x7 & ~x207 ) | ( x7 & n322 ) | ( ~x207 & n322 ) ;
  assign n654 = ( ~x207 & n322 ) | ( ~x207 & n623 ) | ( n322 & n623 ) ;
  assign n655 = n653 & ~n654 ;
  assign n656 = ( n294 & n651 ) | ( n294 & ~n655 ) | ( n651 & ~n655 ) ;
  assign n657 = ~n652 & n656 ;
  assign n658 = ( n640 & ~n641 ) | ( n640 & n657 ) | ( ~n641 & n657 ) ;
  assign n659 = x7 & ~n623 ;
  assign n660 = ~x208 & n659 ;
  assign n661 = n329 & n659 ;
  assign n662 = n660 & ~n661 ;
  assign n663 = n660 | n661 ;
  assign n664 = ( ~n660 & n662 ) | ( ~n660 & n663 ) | ( n662 & n663 ) ;
  assign n665 = ( n640 & ~n641 ) | ( n640 & n664 ) | ( ~n641 & n664 ) ;
  assign n666 = n658 & ~n665 ;
  assign n667 = ( n634 & n637 ) | ( n634 & ~n666 ) | ( n637 & ~n666 ) ;
  assign n668 = ( n316 & n626 ) | ( n316 & n630 ) | ( n626 & n630 ) ;
  assign n669 = n666 & ~n668 ;
  assign n670 = ( n634 & ~n667 ) | ( n634 & n669 ) | ( ~n667 & n669 ) ;
  assign n671 = ( ~n640 & n641 ) | ( ~n640 & n648 ) | ( n641 & n648 ) ;
  assign n672 = n665 | n671 ;
  assign n673 = n294 | n651 ;
  assign n674 = n672 | n673 ;
  assign n675 = n640 & ~n648 ;
  assign n676 = ( ~n641 & n664 ) | ( ~n641 & n675 ) | ( n664 & n675 ) ;
  assign n677 = ~n664 & n676 ;
  assign n678 = ( n646 & ~n655 ) | ( n646 & n664 ) | ( ~n655 & n664 ) ;
  assign n679 = ~n664 & n678 ;
  assign n680 = x7 & ~n322 ;
  assign n681 = ( ~x207 & n623 ) | ( ~x207 & n680 ) | ( n623 & n680 ) ;
  assign n682 = ~n623 & n681 ;
  assign n683 = ( n660 & ~n661 ) | ( n660 & n682 ) | ( ~n661 & n682 ) ;
  assign n684 = n679 | n683 ;
  assign n685 = ( n674 & n677 ) | ( n674 & n684 ) | ( n677 & n684 ) ;
  assign n686 = n655 & ~n684 ;
  assign n687 = ( n674 & ~n685 ) | ( n674 & n686 ) | ( ~n685 & n686 ) ;
  assign n688 = x202 & n273 ;
  assign n689 = x29 & ~n259 ;
  assign n690 = ( ~n273 & n688 ) | ( ~n273 & n689 ) | ( n688 & n689 ) ;
  assign n691 = ~n623 & n690 ;
  assign n692 = ~x213 & n691 ;
  assign n693 = n430 & n691 ;
  assign n694 = n692 & ~n693 ;
  assign n695 = n692 | n693 ;
  assign n696 = ( ~n692 & n694 ) | ( ~n692 & n695 ) | ( n694 & n695 ) ;
  assign n697 = ( ~x211 & n475 ) | ( ~x211 & n690 ) | ( n475 & n690 ) ;
  assign n698 = ( ~x211 & n475 ) | ( ~x211 & n623 ) | ( n475 & n623 ) ;
  assign n699 = n697 & ~n698 ;
  assign n700 = ~x210 & n690 ;
  assign n701 = ( ~n494 & n623 ) | ( ~n494 & n700 ) | ( n623 & n700 ) ;
  assign n702 = ~n623 & n701 ;
  assign n703 = ( n696 & ~n699 ) | ( n696 & n702 ) | ( ~n699 & n702 ) ;
  assign n704 = ( ~x210 & n494 ) | ( ~x210 & n690 ) | ( n494 & n690 ) ;
  assign n705 = ( ~x210 & n494 ) | ( ~x210 & n623 ) | ( n494 & n623 ) ;
  assign n706 = n704 & ~n705 ;
  assign n707 = n336 & ~n623 ;
  assign n708 = n690 & n707 ;
  assign n709 = ~x209 & n691 ;
  assign n710 = ~n708 & n709 ;
  assign n711 = ( n696 & ~n706 ) | ( n696 & n710 ) | ( ~n706 & n710 ) ;
  assign n712 = ~n696 & n711 ;
  assign n713 = ~n699 & n712 ;
  assign n714 = ( ~n696 & n703 ) | ( ~n696 & n713 ) | ( n703 & n713 ) ;
  assign n715 = ~x211 & n690 ;
  assign n716 = ( ~n475 & n623 ) | ( ~n475 & n715 ) | ( n623 & n715 ) ;
  assign n717 = ~n623 & n716 ;
  assign n718 = ( n692 & ~n693 ) | ( n692 & n717 ) | ( ~n693 & n717 ) ;
  assign n719 = n714 | n718 ;
  assign n720 = ( n670 & n687 ) | ( n670 & ~n719 ) | ( n687 & ~n719 ) ;
  assign n721 = n708 & ~n709 ;
  assign n722 = n708 | n709 ;
  assign n723 = ( ~n708 & n721 ) | ( ~n708 & n722 ) | ( n721 & n722 ) ;
  assign n724 = n706 | n723 ;
  assign n725 = ( ~n696 & n699 ) | ( ~n696 & n724 ) | ( n699 & n724 ) ;
  assign n726 = n696 | n725 ;
  assign n727 = ~n719 & n726 ;
  assign n728 = ( ~n670 & n720 ) | ( ~n670 & n727 ) | ( n720 & n727 ) ;
  assign n729 = n402 & ~n590 ;
  assign n730 = n620 & n729 ;
  assign n731 = ~n252 & n423 ;
  assign n732 = ( n387 & n730 ) | ( n387 & n731 ) | ( n730 & n731 ) ;
  assign n733 = ~n387 & n732 ;
  assign y0 = x114 ;
  assign y1 = x115 ;
  assign y2 = x116 ;
  assign y3 = x117 ;
  assign y4 = x118 ;
  assign y5 = x119 ;
  assign y6 = x120 ;
  assign y7 = x121 ;
  assign y8 = x122 ;
  assign y9 = x123 ;
  assign y10 = x124 ;
  assign y11 = x125 ;
  assign y12 = x126 ;
  assign y13 = x127 ;
  assign y14 = x128 ;
  assign y15 = x129 ;
  assign y16 = x130 ;
  assign y17 = x131 ;
  assign y18 = x132 ;
  assign y19 = x133 ;
  assign y20 = x134 ;
  assign y21 = x135 ;
  assign y22 = x136 ;
  assign y23 = x137 ;
  assign y24 = x138 ;
  assign y25 = x139 ;
  assign y26 = x140 ;
  assign y27 = x141 ;
  assign y28 = x142 ;
  assign y29 = x143 ;
  assign y30 = x144 ;
  assign y31 = x145 ;
  assign y32 = x146 ;
  assign y33 = x147 ;
  assign y34 = x148 ;
  assign y35 = x149 ;
  assign y36 = x150 ;
  assign y37 = x151 ;
  assign y38 = x152 ;
  assign y39 = x153 ;
  assign y40 = x154 ;
  assign y41 = x155 ;
  assign y42 = x156 ;
  assign y43 = x157 ;
  assign y44 = x158 ;
  assign y45 = x159 ;
  assign y46 = x160 ;
  assign y47 = x161 ;
  assign y48 = x162 ;
  assign y49 = x163 ;
  assign y50 = x164 ;
  assign y51 = x165 ;
  assign y52 = x166 ;
  assign y53 = x167 ;
  assign y54 = x168 ;
  assign y55 = x169 ;
  assign y56 = x170 ;
  assign y57 = x171 ;
  assign y58 = x172 ;
  assign y59 = x173 ;
  assign y60 = x174 ;
  assign y61 = x175 ;
  assign y62 = x176 ;
  assign y63 = x177 ;
  assign y64 = x178 ;
  assign y65 = x179 ;
  assign y66 = x180 ;
  assign y67 = x181 ;
  assign y68 = x182 ;
  assign y69 = x183 ;
  assign y70 = x184 ;
  assign y71 = x185 ;
  assign y72 = x186 ;
  assign y73 = x187 ;
  assign y74 = x188 ;
  assign y75 = x189 ;
  assign y76 = x190 ;
  assign y77 = x190 ;
  assign y78 = x190 ;
  assign y79 = x199 ;
  assign y80 = x199 ;
  assign y81 = x212 ;
  assign y82 = x212 ;
  assign y83 = x212 ;
  assign y84 = ~x31 ;
  assign y85 = ~x105 ;
  assign y86 = ~x63 ;
  assign y87 = ~x75 ;
  assign y88 = ~x52 ;
  assign y89 = ~x95 ;
  assign y90 = ~x42 ;
  assign y91 = ~x85 ;
  assign y92 = ~n236 ;
  assign y93 = ~n238 ;
  assign y94 = x190 ;
  assign y95 = n239 ;
  assign y96 = ~n240 ;
  assign y97 = ~n241 ;
  assign y98 = ~n242 ;
  assign y99 = n249 ;
  assign y100 = ~n249 ;
  assign y101 = ~n252 ;
  assign y102 = ~n259 ;
  assign y103 = ~n266 ;
  assign y104 = ~n273 ;
  assign y105 = ~n280 ;
  assign y106 = ~n287 ;
  assign y107 = ~n294 ;
  assign y108 = ~n302 ;
  assign y109 = ~n305 ;
  assign y110 = ~n309 ;
  assign y111 = n316 ;
  assign y112 = n294 ;
  assign y113 = n287 ;
  assign y114 = n280 ;
  assign y115 = n322 ;
  assign y116 = n329 ;
  assign y117 = n336 ;
  assign y118 = n346 ;
  assign y119 = n346 ;
  assign y120 = n349 ;
  assign y121 = n349 ;
  assign y122 = n351 ;
  assign y123 = n355 ;
  assign y124 = n355 ;
  assign y125 = ~n365 ;
  assign y126 = n387 ;
  assign y127 = ~n402 ;
  assign y128 = ~n423 ;
  assign y129 = n550 ;
  assign y130 = ~n550 ;
  assign y131 = ~n564 ;
  assign y132 = n590 ;
  assign y133 = n611 ;
  assign y134 = n611 ;
  assign y135 = ~n620 ;
  assign y136 = ~n728 ;
  assign y137 = 1'b0 ;
  assign y138 = n733 ;
  assign y139 = ~n733 ;
endmodule
