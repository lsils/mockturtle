module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 ;
  wire n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 ;
  assign n136 = ( x9 & ~x11 ) | ( x9 & x14 ) | ( ~x11 & x14 ) ;
  assign n137 = ( ~x9 & x11 ) | ( ~x9 & n136 ) | ( x11 & n136 ) ;
  assign n138 = ( ~x14 & n136 ) | ( ~x14 & n137 ) | ( n136 & n137 ) ;
  assign n139 = ( x2 & x5 ) | ( x2 & n138 ) | ( x5 & n138 ) ;
  assign n140 = ( x2 & n138 ) | ( x2 & ~n139 ) | ( n138 & ~n139 ) ;
  assign n141 = ( x5 & ~n139 ) | ( x5 & n140 ) | ( ~n139 & n140 ) ;
  assign n142 = ~x7 & n141 ;
  assign n143 = x7 & ~n141 ;
  assign n144 = n142 | n143 ;
  assign n145 = x18 & ~x32 ;
  assign n146 = x22 & n145 ;
  assign n147 = n144 | n146 ;
  assign n148 = n144 & n146 ;
  assign n149 = n147 & ~n148 ;
  assign n150 = x30 & n149 ;
  assign n151 = ( x27 & n149 ) | ( x27 & n150 ) | ( n149 & n150 ) ;
  assign n152 = ( x27 & ~n149 ) | ( x27 & n150 ) | ( ~n149 & n150 ) ;
  assign n153 = ( n149 & ~n151 ) | ( n149 & n152 ) | ( ~n151 & n152 ) ;
  assign n158 = ( x1 & ~x4 ) | ( x1 & x7 ) | ( ~x4 & x7 ) ;
  assign n159 = ( ~x1 & x4 ) | ( ~x1 & n158 ) | ( x4 & n158 ) ;
  assign n160 = ( ~x7 & n158 ) | ( ~x7 & n159 ) | ( n158 & n159 ) ;
  assign n112 = ( x8 & ~x13 ) | ( x8 & x15 ) | ( ~x13 & x15 ) ;
  assign n113 = ( ~x8 & x13 ) | ( ~x8 & n112 ) | ( x13 & n112 ) ;
  assign n114 = ( ~x15 & n112 ) | ( ~x15 & n113 ) | ( n112 & n113 ) ;
  assign n102 = x23 | x32 ;
  assign n154 = x17 & ~n102 ;
  assign n155 = x14 & ~n154 ;
  assign n156 = ~x14 & n154 ;
  assign n157 = n155 | n156 ;
  assign n161 = ( n114 & n157 ) | ( n114 & n160 ) | ( n157 & n160 ) ;
  assign n162 = ( n114 & n157 ) | ( n114 & ~n161 ) | ( n157 & ~n161 ) ;
  assign n163 = ( n160 & ~n161 ) | ( n160 & n162 ) | ( ~n161 & n162 ) ;
  assign n164 = ~x10 & n163 ;
  assign n165 = x10 & ~n163 ;
  assign n166 = n164 | n165 ;
  assign n167 = x30 & n166 ;
  assign n168 = ( x26 & n166 ) | ( x26 & n167 ) | ( n166 & n167 ) ;
  assign n169 = ( x26 & ~n166 ) | ( x26 & n167 ) | ( ~n166 & n167 ) ;
  assign n170 = ( n166 & ~n168 ) | ( n166 & n169 ) | ( ~n168 & n169 ) ;
  assign n171 = n153 | n170 ;
  assign n36 = x22 & ~x23 ;
  assign n37 = x31 & ~x32 ;
  assign n38 = ( ~x22 & n36 ) | ( ~x22 & n37 ) | ( n36 & n37 ) ;
  assign n34 = ~x23 & x32 ;
  assign n35 = ( ~x22 & x32 ) | ( ~x22 & n34 ) | ( x32 & n34 ) ;
  assign n39 = ( ~x28 & n35 ) | ( ~x28 & n38 ) | ( n35 & n38 ) ;
  assign n40 = x30 & ~n39 ;
  assign n41 = ( x30 & n38 ) | ( x30 & ~n40 ) | ( n38 & ~n40 ) ;
  assign n64 = x16 & x30 ;
  assign n42 = ( x0 & ~x1 ) | ( x0 & x2 ) | ( ~x1 & x2 ) ;
  assign n43 = ( ~x0 & x1 ) | ( ~x0 & n42 ) | ( x1 & n42 ) ;
  assign n44 = ( ~x2 & n42 ) | ( ~x2 & n43 ) | ( n42 & n43 ) ;
  assign n45 = ( x4 & x5 ) | ( x4 & n44 ) | ( x5 & n44 ) ;
  assign n46 = ( x4 & n44 ) | ( x4 & ~n45 ) | ( n44 & ~n45 ) ;
  assign n47 = ( x5 & ~n45 ) | ( x5 & n46 ) | ( ~n45 & n46 ) ;
  assign n48 = ~x6 & n47 ;
  assign n49 = x6 & ~n47 ;
  assign n50 = n48 | n49 ;
  assign n51 = ( ~x3 & x7 ) | ( ~x3 & n50 ) | ( x7 & n50 ) ;
  assign n52 = ( x3 & ~n50 ) | ( x3 & n51 ) | ( ~n50 & n51 ) ;
  assign n53 = ( ~x7 & n51 ) | ( ~x7 & n52 ) | ( n51 & n52 ) ;
  assign n54 = ( x9 & ~x14 ) | ( x9 & x15 ) | ( ~x14 & x15 ) ;
  assign n55 = ( ~x9 & x14 ) | ( ~x9 & n54 ) | ( x14 & n54 ) ;
  assign n56 = ( ~x15 & n54 ) | ( ~x15 & n55 ) | ( n54 & n55 ) ;
  assign n57 = x20 & ~x32 ;
  assign n58 = ( x8 & n56 ) | ( x8 & ~n57 ) | ( n56 & ~n57 ) ;
  assign n59 = ( ~n56 & n57 ) | ( ~n56 & n58 ) | ( n57 & n58 ) ;
  assign n60 = ( ~x8 & n58 ) | ( ~x8 & n59 ) | ( n58 & n59 ) ;
  assign n61 = ~n53 & n60 ;
  assign n62 = n53 & n60 ;
  assign n63 = ( n53 & n61 ) | ( n53 & ~n62 ) | ( n61 & ~n62 ) ;
  assign n65 = ( x16 & x23 ) | ( x16 & x30 ) | ( x23 & x30 ) ;
  assign n66 = n63 & n65 ;
  assign n67 = ( ~x30 & n63 ) | ( ~x30 & n65 ) | ( n63 & n65 ) ;
  assign n68 = ( n64 & ~n66 ) | ( n64 & n67 ) | ( ~n66 & n67 ) ;
  assign n86 = x17 & x30 ;
  assign n87 = ( x17 & x23 ) | ( x17 & n86 ) | ( x23 & n86 ) ;
  assign n72 = x21 & ~x32 ;
  assign n73 = ( x3 & x13 ) | ( x3 & ~n72 ) | ( x13 & ~n72 ) ;
  assign n74 = ( ~x3 & n72 ) | ( ~x3 & n73 ) | ( n72 & n73 ) ;
  assign n75 = ( ~x13 & n73 ) | ( ~x13 & n74 ) | ( n73 & n74 ) ;
  assign n69 = ( x10 & ~x11 ) | ( x10 & x12 ) | ( ~x11 & x12 ) ;
  assign n70 = ( ~x10 & x11 ) | ( ~x10 & n69 ) | ( x11 & n69 ) ;
  assign n71 = ( ~x12 & n69 ) | ( ~x12 & n70 ) | ( n69 & n70 ) ;
  assign n76 = ( n44 & n56 ) | ( n44 & n71 ) | ( n56 & n71 ) ;
  assign n77 = ( n56 & n71 ) | ( n56 & ~n76 ) | ( n71 & ~n76 ) ;
  assign n78 = ( n44 & ~n76 ) | ( n44 & n77 ) | ( ~n76 & n77 ) ;
  assign n79 = n75 & n78 ;
  assign n80 = n75 | n78 ;
  assign n81 = ~n79 & n80 ;
  assign n82 = x30 & n81 ;
  assign n83 = ( x24 & n81 ) | ( x24 & n82 ) | ( n81 & n82 ) ;
  assign n84 = ( x24 & ~n81 ) | ( x24 & n82 ) | ( ~n81 & n82 ) ;
  assign n85 = ( n81 & ~n83 ) | ( n81 & n84 ) | ( ~n83 & n84 ) ;
  assign n88 = x19 & x30 ;
  assign n89 = ( x19 & ~x22 ) | ( x19 & n88 ) | ( ~x22 & n88 ) ;
  assign n90 = n85 & ~n89 ;
  assign n91 = ( n68 & n87 ) | ( n68 & ~n90 ) | ( n87 & ~n90 ) ;
  assign n92 = n68 & ~n91 ;
  assign n93 = n56 & ~n71 ;
  assign n94 = n56 | n71 ;
  assign n95 = ( ~n56 & n93 ) | ( ~n56 & n94 ) | ( n93 & n94 ) ;
  assign n96 = ( x4 & x5 ) | ( x4 & n95 ) | ( x5 & n95 ) ;
  assign n97 = ( x4 & n95 ) | ( x4 & ~n96 ) | ( n95 & ~n96 ) ;
  assign n98 = ( x5 & ~n96 ) | ( x5 & n97 ) | ( ~n96 & n97 ) ;
  assign n99 = ~x6 & n98 ;
  assign n100 = x6 & ~n98 ;
  assign n101 = n99 | n100 ;
  assign n103 = x16 & ~n102 ;
  assign n104 = x0 & ~n103 ;
  assign n105 = ~x0 & n103 ;
  assign n106 = n104 | n105 ;
  assign n107 = ( x25 & n101 ) | ( x25 & n106 ) | ( n101 & n106 ) ;
  assign n108 = ~x30 & n107 ;
  assign n109 = ( n101 & n106 ) | ( n101 & ~n107 ) | ( n106 & ~n107 ) ;
  assign n110 = ~x30 & n109 ;
  assign n111 = ( x25 & ~n108 ) | ( x25 & n110 ) | ( ~n108 & n110 ) ;
  assign n129 = x18 & x30 ;
  assign n115 = ( x3 & x6 ) | ( x3 & n114 ) | ( x6 & n114 ) ;
  assign n116 = ( x3 & n114 ) | ( x3 & ~n115 ) | ( n114 & ~n115 ) ;
  assign n117 = ( x6 & ~n115 ) | ( x6 & n116 ) | ( ~n115 & n116 ) ;
  assign n118 = ~x9 & n117 ;
  assign n119 = x9 & ~n117 ;
  assign n120 = n118 | n119 ;
  assign n121 = x19 & ~x32 ;
  assign n122 = x22 & n121 ;
  assign n123 = x12 & ~n122 ;
  assign n124 = ~x12 & n122 ;
  assign n125 = n123 | n124 ;
  assign n126 = n120 | n125 ;
  assign n127 = n120 & ~n125 ;
  assign n128 = ( ~n120 & n126 ) | ( ~n120 & n127 ) | ( n126 & n127 ) ;
  assign n130 = ( x18 & ~x22 ) | ( x18 & x30 ) | ( ~x22 & x30 ) ;
  assign n131 = n128 & n130 ;
  assign n132 = ( ~x30 & n128 ) | ( ~x30 & n130 ) | ( n128 & n130 ) ;
  assign n133 = ( n129 & ~n131 ) | ( n129 & n132 ) | ( ~n131 & n132 ) ;
  assign n134 = n111 & ~n133 ;
  assign n135 = n92 & n134 ;
  assign n172 = n41 & n135 ;
  assign n173 = ~n171 & n172 ;
  assign n174 = x0 & ~n173 ;
  assign n175 = ~x0 & n173 ;
  assign n176 = n174 | n175 ;
  assign n179 = ~n153 & n170 ;
  assign n177 = n111 | n133 ;
  assign n178 = n92 & ~n177 ;
  assign n180 = n41 & n178 ;
  assign n181 = n179 & n180 ;
  assign n182 = x1 & ~n181 ;
  assign n183 = ~x1 & n181 ;
  assign n184 = n182 | n183 ;
  assign n185 = n153 & ~n170 ;
  assign n186 = n180 & n185 ;
  assign n187 = x2 & ~n186 ;
  assign n188 = ~x2 & n186 ;
  assign n189 = n187 | n188 ;
  assign n190 = ~n111 & n133 ;
  assign n191 = n92 & n190 ;
  assign n192 = n41 & n191 ;
  assign n193 = ~n171 & n192 ;
  assign n194 = x3 & ~n193 ;
  assign n195 = ~x3 & n193 ;
  assign n196 = n194 | n195 ;
  assign n197 = ( ~x29 & n35 ) | ( ~x29 & n38 ) | ( n35 & n38 ) ;
  assign n198 = x30 & ~n197 ;
  assign n199 = ( x30 & n38 ) | ( x30 & ~n198 ) | ( n38 & ~n198 ) ;
  assign n200 = n111 & n133 ;
  assign n201 = n92 & n200 ;
  assign n202 = n199 & n201 ;
  assign n203 = n185 & n202 ;
  assign n204 = x9 & ~n203 ;
  assign n205 = ~x9 & n203 ;
  assign n206 = n204 | n205 ;
  assign n207 = n153 & n170 ;
  assign n208 = n135 & n199 ;
  assign n209 = n207 & n208 ;
  assign n210 = x14 & ~n209 ;
  assign n211 = ~x14 & n209 ;
  assign n212 = n210 | n211 ;
  assign n213 = n179 & n202 ;
  assign n214 = x15 & ~n213 ;
  assign n215 = ~x15 & n213 ;
  assign n216 = n214 | n215 ;
  assign n217 = n85 | n89 ;
  assign n218 = n68 & ~n217 ;
  assign n219 = ~n87 & n218 ;
  assign n220 = n134 & n219 ;
  assign n221 = n41 & n220 ;
  assign n222 = n179 & n221 ;
  assign n223 = x4 & ~n222 ;
  assign n224 = ~x4 & n222 ;
  assign n225 = n223 | n224 ;
  assign n226 = n185 & n221 ;
  assign n227 = x5 & ~n226 ;
  assign n228 = ~x5 & n226 ;
  assign n229 = n227 | n228 ;
  assign n230 = n200 & n219 ;
  assign n231 = n41 & n230 ;
  assign n232 = ~n171 & n231 ;
  assign n233 = x6 & ~n232 ;
  assign n234 = ~x6 & n232 ;
  assign n235 = n233 | n234 ;
  assign n236 = ~n177 & n219 ;
  assign n237 = n41 & n236 ;
  assign n238 = n207 & n237 ;
  assign n239 = x7 & ~n238 ;
  assign n240 = ~x7 & n238 ;
  assign n241 = n239 | n240 ;
  assign n242 = n190 & n219 ;
  assign n243 = n199 & n242 ;
  assign n244 = n179 & n243 ;
  assign n245 = x8 & ~n244 ;
  assign n246 = ~x8 & n244 ;
  assign n247 = n245 | n246 ;
  assign n248 = n68 | n87 ;
  assign n249 = n85 & ~n248 ;
  assign n250 = ~n89 & n249 ;
  assign n251 = n134 & n250 ;
  assign n252 = n199 & n251 ;
  assign n253 = n179 & n252 ;
  assign n254 = x10 & ~n253 ;
  assign n255 = ~x10 & n253 ;
  assign n256 = n254 | n255 ;
  assign n257 = n185 & n252 ;
  assign n258 = x11 & ~n257 ;
  assign n259 = ~x11 & n257 ;
  assign n260 = n258 | n259 ;
  assign n261 = n200 & n250 ;
  assign n262 = n199 & n261 ;
  assign n263 = ~n171 & n262 ;
  assign n264 = x12 & ~n263 ;
  assign n265 = ~x12 & n263 ;
  assign n266 = n264 | n265 ;
  assign n267 = n179 & n250 ;
  assign n268 = ( n190 & ~n199 ) | ( n190 & n267 ) | ( ~n199 & n267 ) ;
  assign n269 = n199 & n268 ;
  assign n270 = ~x13 & n269 ;
  assign n271 = x13 | n269 ;
  assign n272 = ( ~n269 & n270 ) | ( ~n269 & n271 ) | ( n270 & n271 ) ;
  assign n278 = n217 | n248 ;
  assign n279 = n190 & ~n278 ;
  assign n280 = n89 & ~n177 ;
  assign n281 = ( ~n85 & n248 ) | ( ~n85 & n280 ) | ( n248 & n280 ) ;
  assign n282 = ~n248 & n281 ;
  assign n286 = n38 & n179 ;
  assign n287 = ( ~n177 & n278 ) | ( ~n177 & n286 ) | ( n278 & n286 ) ;
  assign n288 = ~n278 & n287 ;
  assign n283 = n38 & ~n177 ;
  assign n284 = ( n185 & n278 ) | ( n185 & n283 ) | ( n278 & n283 ) ;
  assign n285 = ~n278 & n284 ;
  assign n289 = n219 & ~n250 ;
  assign n273 = n38 & ~n171 ;
  assign n290 = ~n177 & n273 ;
  assign n291 = ( n250 & n289 ) | ( n250 & n290 ) | ( n289 & n290 ) ;
  assign n292 = ( n273 & ~n278 ) | ( n273 & n291 ) | ( ~n278 & n291 ) ;
  assign n293 = n134 & ~n292 ;
  assign n294 = ( n134 & n291 ) | ( n134 & ~n293 ) | ( n291 & ~n293 ) ;
  assign n295 = n285 | n294 ;
  assign n296 = n288 | n295 ;
  assign n297 = ( ~n279 & n282 ) | ( ~n279 & n296 ) | ( n282 & n296 ) ;
  assign n298 = n273 | n296 ;
  assign n299 = ( n279 & n297 ) | ( n279 & n298 ) | ( n297 & n298 ) ;
  assign n274 = ~n68 & n87 ;
  assign n275 = ~n217 & n274 ;
  assign n276 = ( n177 & n273 ) | ( n177 & ~n275 ) | ( n273 & ~n275 ) ;
  assign n277 = n273 & ~n276 ;
  assign n300 = n179 & n199 ;
  assign n322 = n201 & ~n300 ;
  assign n301 = ( n41 & ~n171 ) | ( n41 & n181 ) | ( ~n171 & n181 ) ;
  assign n302 = n135 & ~n301 ;
  assign n303 = ( n135 & n181 ) | ( n135 & ~n302 ) | ( n181 & ~n302 ) ;
  assign n304 = n193 | n303 ;
  assign n305 = ( n186 & ~n222 ) | ( n186 & n304 ) | ( ~n222 & n304 ) ;
  assign n306 = n222 | n305 ;
  assign n307 = n232 | n306 ;
  assign n308 = ( n226 & ~n238 ) | ( n226 & n307 ) | ( ~n238 & n307 ) ;
  assign n309 = n238 | n308 ;
  assign n310 = n190 & n250 ;
  assign n311 = n300 & n310 ;
  assign n312 = n185 & n199 ;
  assign n313 = n201 & n312 ;
  assign n314 = n242 | n313 ;
  assign n315 = ( n300 & n313 ) | ( n300 & n314 ) | ( n313 & n314 ) ;
  assign n316 = ( ~n300 & n312 ) | ( ~n300 & n315 ) | ( n312 & n315 ) ;
  assign n317 = n251 | n315 ;
  assign n318 = ( n300 & n316 ) | ( n300 & n317 ) | ( n316 & n317 ) ;
  assign n319 = n209 | n318 ;
  assign n320 = ( ~n263 & n311 ) | ( ~n263 & n319 ) | ( n311 & n319 ) ;
  assign n321 = n263 | n320 ;
  assign n323 = n309 | n321 ;
  assign n324 = ( n201 & ~n322 ) | ( n201 & n323 ) | ( ~n322 & n323 ) ;
  assign n325 = n277 | n324 ;
  assign n326 = n299 | n325 ;
  assign n334 = ~x31 & n326 ;
  assign n330 = n85 | n87 ;
  assign n327 = n133 | n170 ;
  assign n328 = ( n111 & ~n153 ) | ( n111 & n327 ) | ( ~n153 & n327 ) ;
  assign n329 = n153 | n328 ;
  assign n331 = n68 | n329 ;
  assign n332 = ( ~n89 & n330 ) | ( ~n89 & n331 ) | ( n330 & n331 ) ;
  assign n333 = n89 | n332 ;
  assign n335 = ~x32 & n333 ;
  assign n336 = ( ~n326 & n334 ) | ( ~n326 & n335 ) | ( n334 & n335 ) ;
  assign n337 = x30 & n324 ;
  assign n338 = x16 & n337 ;
  assign n339 = ( n53 & ~n60 ) | ( n53 & n338 ) | ( ~n60 & n338 ) ;
  assign n340 = ( n53 & n338 ) | ( n53 & ~n339 ) | ( n338 & ~n339 ) ;
  assign n341 = ( n60 & n339 ) | ( n60 & ~n340 ) | ( n339 & ~n340 ) ;
  assign n342 = ~x32 & n341 ;
  assign n343 = ( x31 & n341 ) | ( x31 & n342 ) | ( n341 & n342 ) ;
  assign n344 = x24 & n324 ;
  assign n345 = x30 & n344 ;
  assign n346 = n81 | n345 ;
  assign n347 = n81 & n345 ;
  assign n348 = n346 & ~n347 ;
  assign n349 = ~x32 & n348 ;
  assign n350 = ( x31 & n348 ) | ( x31 & n349 ) | ( n348 & n349 ) ;
  assign n351 = x26 & n324 ;
  assign n352 = x30 & n351 ;
  assign n353 = n166 | n352 ;
  assign n354 = n166 & n352 ;
  assign n355 = n353 & ~n354 ;
  assign n356 = ~x32 & n355 ;
  assign n357 = ( x31 & n355 ) | ( x31 & n356 ) | ( n355 & n356 ) ;
  assign n358 = x27 & n324 ;
  assign n359 = x30 & n358 ;
  assign n360 = n149 | n359 ;
  assign n361 = n149 & n359 ;
  assign n362 = n360 & ~n361 ;
  assign n363 = ~x32 & n362 ;
  assign n364 = ( x31 & n362 ) | ( x31 & n363 ) | ( n362 & n363 ) ;
  assign n365 = x18 & n337 ;
  assign n366 = ~n128 & n365 ;
  assign n367 = ~x31 & x32 ;
  assign n368 = ( n128 & ~n365 ) | ( n128 & n367 ) | ( ~n365 & n367 ) ;
  assign n369 = ( n366 & ~n367 ) | ( n366 & n368 ) | ( ~n367 & n368 ) ;
  assign n381 = ~x20 & x32 ;
  assign n382 = ( ~x28 & x32 ) | ( ~x28 & n381 ) | ( x32 & n381 ) ;
  assign n370 = n222 | n232 ;
  assign n371 = ( n226 & ~n238 ) | ( n226 & n370 ) | ( ~n238 & n370 ) ;
  assign n372 = n238 | n371 ;
  assign n373 = n186 | n372 ;
  assign n374 = ( ~n193 & n303 ) | ( ~n193 & n373 ) | ( n303 & n373 ) ;
  assign n375 = n193 | n374 ;
  assign n376 = n53 | n375 ;
  assign n377 = ( x32 & n53 ) | ( x32 & ~n375 ) | ( n53 & ~n375 ) ;
  assign n378 = x28 | n53 ;
  assign n379 = ( x32 & n53 ) | ( x32 & n378 ) | ( n53 & n378 ) ;
  assign n380 = ( n376 & n377 ) | ( n376 & ~n379 ) | ( n377 & ~n379 ) ;
  assign n383 = n380 | n382 ;
  assign n384 = ~n380 & n382 ;
  assign n385 = ( ~n382 & n383 ) | ( ~n382 & n384 ) | ( n383 & n384 ) ;
  assign n402 = ~x21 & x32 ;
  assign n403 = ( ~x29 & x32 ) | ( ~x29 & n402 ) | ( x32 & n402 ) ;
  assign n390 = n251 & n300 ;
  assign n391 = ( n251 & n312 ) | ( n251 & n390 ) | ( n312 & n390 ) ;
  assign n386 = n209 | n300 ;
  assign n387 = ( n201 & n209 ) | ( n201 & n386 ) | ( n209 & n386 ) ;
  assign n388 = n263 | n387 ;
  assign n389 = n311 | n388 ;
  assign n392 = n315 | n389 ;
  assign n393 = n391 | n392 ;
  assign n394 = ( ~x8 & x13 ) | ( ~x8 & n95 ) | ( x13 & n95 ) ;
  assign n395 = ( x8 & ~n95 ) | ( x8 & n394 ) | ( ~n95 & n394 ) ;
  assign n396 = ( ~x13 & n394 ) | ( ~x13 & n395 ) | ( n394 & n395 ) ;
  assign n397 = n393 | n396 ;
  assign n398 = ( x32 & ~n393 ) | ( x32 & n396 ) | ( ~n393 & n396 ) ;
  assign n399 = x29 | n396 ;
  assign n400 = ( x32 & n396 ) | ( x32 & n399 ) | ( n396 & n399 ) ;
  assign n401 = ( n397 & n398 ) | ( n397 & ~n400 ) | ( n398 & ~n400 ) ;
  assign n404 = n401 | n403 ;
  assign n405 = ~n401 & n403 ;
  assign n406 = ( ~n403 & n404 ) | ( ~n403 & n405 ) | ( n404 & n405 ) ;
  assign n407 = x25 & n324 ;
  assign n408 = x30 & n407 ;
  assign n409 = n101 & ~n408 ;
  assign n410 = ~n101 & n408 ;
  assign n411 = n409 | n410 ;
  assign n412 = n106 & ~n411 ;
  assign n413 = ( ~n106 & n367 ) | ( ~n106 & n411 ) | ( n367 & n411 ) ;
  assign n414 = ( ~n367 & n412 ) | ( ~n367 & n413 ) | ( n412 & n413 ) ;
  assign y0 = n176 ;
  assign y1 = n184 ;
  assign y2 = n189 ;
  assign y3 = n196 ;
  assign y4 = n206 ;
  assign y5 = n212 ;
  assign y6 = n216 ;
  assign y7 = n225 ;
  assign y8 = n229 ;
  assign y9 = n235 ;
  assign y10 = n241 ;
  assign y11 = n247 ;
  assign y12 = n256 ;
  assign y13 = n260 ;
  assign y14 = n266 ;
  assign y15 = n272 ;
  assign y16 = ~n336 ;
  assign y17 = n343 ;
  assign y18 = n350 ;
  assign y19 = n357 ;
  assign y20 = n364 ;
  assign y21 = n369 ;
  assign y22 = ~n385 ;
  assign y23 = ~n406 ;
  assign y24 = n414 ;
endmodule
